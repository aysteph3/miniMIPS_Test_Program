
module alu_DW01_add_11 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] ,
         \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] ,
         \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419;
  assign SUM[30] = \A[30] ;
  assign \A[30]  = A[30];
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND_GATE U2 ( .I1(n325), .I2(n4), .O(n1) );
  AND_GATE U3 ( .I1(n1), .I2(n2), .O(n283) );
  OR_GATE U4 ( .I1(n3), .I2(n323), .O(n2) );
  INV_GATE U5 ( .I1(n322), .O(n3) );
  AND_GATE U6 ( .I1(n324), .I2(n322), .O(n4) );
  NAND_GATE U7 ( .I1(n248), .I2(n8), .O(n5) );
  AND_GATE U8 ( .I1(n5), .I2(n6), .O(n239) );
  OR_GATE U9 ( .I1(n7), .I2(n247), .O(n6) );
  INV_GATE U10 ( .I1(n242), .O(n7) );
  AND_GATE U11 ( .I1(n249), .I2(n242), .O(n8) );
  NAND_GATE U12 ( .I1(n207), .I2(n12), .O(n9) );
  AND_GATE U13 ( .I1(n9), .I2(n10), .O(n133) );
  OR_GATE U14 ( .I1(n11), .I2(n206), .O(n10) );
  INV_GATE U15 ( .I1(n136), .O(n11) );
  AND_GATE U16 ( .I1(n208), .I2(n136), .O(n12) );
  AND_GATE U17 ( .I1(n351), .I2(n398), .O(n13) );
  AND_GATE U18 ( .I1(n328), .I2(n331), .O(n14) );
  AND_GATE U19 ( .I1(n293), .I2(n297), .O(n15) );
  AND_GATE U20 ( .I1(n262), .I2(n260), .O(n16) );
  AND_GATE U21 ( .I1(n235), .I2(n233), .O(n17) );
  AND_GATE U22 ( .I1(n215), .I2(n213), .O(n18) );
  AND_GATE U23 ( .I1(n208), .I2(n206), .O(n19) );
  AND_GATE U24 ( .I1(n200), .I2(n198), .O(n20) );
  AND_GATE U25 ( .I1(n377), .I2(n369), .O(n21) );
  AND_GATE U26 ( .I1(n364), .I2(n372), .O(n22) );
  AND_GATE U27 ( .I1(n396), .I2(n403), .O(n23) );
  AND_GATE U28 ( .I1(n330), .I2(n322), .O(n24) );
  AND_GATE U29 ( .I1(n329), .I2(n327), .O(n25) );
  AND_GATE U30 ( .I1(n326), .I2(n333), .O(n26) );
  AND_GATE U31 ( .I1(n256), .I2(n254), .O(n27) );
  AND_GATE U32 ( .I1(n249), .I2(n247), .O(n28) );
  AND_GATE U33 ( .I1(n242), .I2(n240), .O(n29) );
  AND_GATE U34 ( .I1(n228), .I2(n226), .O(n30) );
  AND_GATE U35 ( .I1(n221), .I2(n219), .O(n31) );
  AND_GATE U36 ( .I1(n143), .I2(n34), .O(n32) );
  NOR_GATE U37 ( .I1(n32), .I2(n33), .O(n391) );
  AND_GATE U38 ( .I1(n22), .I2(n370), .O(n33) );
  AND_GATE U39 ( .I1(n173), .I2(n22), .O(n34) );
  NAND_GATE U40 ( .I1(n143), .I2(n37), .O(n35) );
  AND_GATE U41 ( .I1(n35), .I2(n36), .O(n409) );
  OR_GATE U42 ( .I1(n411), .I2(n394), .O(n36) );
  AND_GATE U43 ( .I1(n399), .I2(n412), .O(n37) );
  OR_GATE U44 ( .I1(n22), .I2(n370), .O(n38) );
  NAND_GATE U45 ( .I1(n39), .I2(n413), .O(n410) );
  NOR_GATE U46 ( .I1(n127), .I2(n412), .O(n39) );
  OR_GATE U47 ( .I1(n38), .I2(n393), .O(n392) );
  OR_GATE U48 ( .I1(n404), .I2(n23), .O(n406) );
  OR_GATE U49 ( .I1(n356), .I2(n26), .O(n355) );
  OR_GATE U50 ( .I1(n339), .I2(n25), .O(n345) );
  NAND_GATE U51 ( .I1(n404), .I2(n43), .O(n40) );
  AND_GATE U52 ( .I1(n40), .I2(n41), .O(n400) );
  OR_GATE U53 ( .I1(n42), .I2(n403), .O(n41) );
  INV_GATE U54 ( .I1(n13), .O(n42) );
  AND_GATE U55 ( .I1(n396), .I2(n13), .O(n43) );
  NAND_GATE U56 ( .I1(n402), .I2(n44), .O(n401) );
  AND_GATE U57 ( .I1(n403), .I2(n42), .O(n44) );
  AND_GATE U58 ( .I1(n194), .I2(n198), .O(n45) );
  NAND_GATE U59 ( .I1(n197), .I2(n45), .O(n73) );
  NAND_GATE U60 ( .I1(n199), .I2(n48), .O(n46) );
  NAND_GATE U61 ( .I1(n46), .I2(n47), .O(n61) );
  OR_GATE U62 ( .I1(n194), .I2(n198), .O(n47) );
  AND_GATE U63 ( .I1(n200), .I2(n195), .O(n48) );
  AND3_GATE U64 ( .I1(n280), .I2(n188), .I3(n281), .O(n49) );
  NAND_GATE U65 ( .I1(n379), .I2(n52), .O(n50) );
  AND_GATE U66 ( .I1(n50), .I2(n51), .O(n381) );
  OR_GATE U67 ( .I1(n383), .I2(n365), .O(n51) );
  AND_GATE U68 ( .I1(n367), .I2(n53), .O(n52) );
  INV_GATE U69 ( .I1(n383), .O(n53) );
  AND_GATE U70 ( .I1(n383), .I2(n365), .O(n54) );
  NAND_GATE U71 ( .I1(n305), .I2(n57), .O(n55) );
  AND_GATE U72 ( .I1(n55), .I2(n56), .O(n308) );
  OR_GATE U73 ( .I1(n310), .I2(n307), .O(n56) );
  AND_GATE U74 ( .I1(n149), .I2(n58), .O(n57) );
  INV_GATE U75 ( .I1(n310), .O(n58) );
  AND_GATE U76 ( .I1(n307), .I2(n310), .O(n59) );
  AND_GATE U77 ( .I1(n201), .I2(n62), .O(n60) );
  NOR_GATE U78 ( .I1(n60), .I2(n61), .O(n192) );
  AND_GATE U79 ( .I1(n156), .I2(n195), .O(n62) );
  AND_GATE U80 ( .I1(n201), .I2(n65), .O(n63) );
  NOR_GATE U81 ( .I1(n63), .I2(n64), .O(n202) );
  AND_GATE U82 ( .I1(n20), .I2(n199), .O(n64) );
  AND_GATE U83 ( .I1(n151), .I2(n20), .O(n65) );
  AND_GATE U84 ( .I1(n201), .I2(n68), .O(n66) );
  NOR_GATE U85 ( .I1(n66), .I2(n67), .O(n209) );
  AND_GATE U86 ( .I1(n19), .I2(n207), .O(n67) );
  AND_GATE U87 ( .I1(n157), .I2(n19), .O(n68) );
  AND_GATE U88 ( .I1(n201), .I2(n71), .O(n69) );
  NOR_GATE U89 ( .I1(n69), .I2(n70), .O(n236) );
  AND_GATE U90 ( .I1(n17), .I2(n234), .O(n70) );
  AND_GATE U91 ( .I1(n159), .I2(n17), .O(n71) );
  OR_GATE U92 ( .I1(n376), .I2(n72), .O(n373) );
  AND3_GATE U93 ( .I1(n369), .I2(n377), .I3(n378), .O(n72) );
  OR_GATE U94 ( .I1(n204), .I2(n74), .O(n203) );
  OR_GATE U95 ( .I1(n199), .I2(n20), .O(n74) );
  OR_GATE U96 ( .I1(n211), .I2(n75), .O(n210) );
  OR_GATE U97 ( .I1(n207), .I2(n19), .O(n75) );
  OR_GATE U98 ( .I1(n238), .I2(n76), .O(n237) );
  OR_GATE U99 ( .I1(n234), .I2(n17), .O(n76) );
  INV_GATE U100 ( .I1(n337), .O(n77) );
  NAND_GATE U101 ( .I1(n78), .I2(n338), .O(n335) );
  NOR_GATE U102 ( .I1(n77), .I2(n24), .O(n78) );
  NAND_GATE U103 ( .I1(n305), .I2(n82), .O(n79) );
  AND_GATE U104 ( .I1(n79), .I2(n80), .O(n313) );
  OR_GATE U105 ( .I1(n81), .I2(n284), .O(n80) );
  INV_GATE U106 ( .I1(n15), .O(n81) );
  AND_GATE U107 ( .I1(n294), .I2(n15), .O(n82) );
  NAND_GATE U108 ( .I1(n339), .I2(n86), .O(n83) );
  AND_GATE U109 ( .I1(n83), .I2(n84), .O(n341) );
  OR_GATE U110 ( .I1(n85), .I2(n327), .O(n84) );
  INV_GATE U111 ( .I1(n14), .O(n85) );
  AND_GATE U112 ( .I1(n329), .I2(n14), .O(n86) );
  NAND_GATE U113 ( .I1(n315), .I2(n87), .O(n314) );
  AND_GATE U114 ( .I1(n284), .I2(n81), .O(n87) );
  NAND_GATE U115 ( .I1(n343), .I2(n88), .O(n342) );
  AND_GATE U116 ( .I1(n327), .I2(n85), .O(n88) );
  AND_GATE U117 ( .I1(n201), .I2(n91), .O(n89) );
  NOR_GATE U118 ( .I1(n89), .I2(n90), .O(n216) );
  AND_GATE U119 ( .I1(n18), .I2(n214), .O(n90) );
  AND_GATE U120 ( .I1(n152), .I2(n18), .O(n91) );
  AND_GATE U121 ( .I1(n201), .I2(n94), .O(n92) );
  NOR_GATE U122 ( .I1(n92), .I2(n93), .O(n222) );
  AND_GATE U123 ( .I1(n31), .I2(n220), .O(n93) );
  AND_GATE U124 ( .I1(n158), .I2(n31), .O(n94) );
  AND_GATE U125 ( .I1(n201), .I2(n97), .O(n95) );
  NOR_GATE U126 ( .I1(n95), .I2(n96), .O(n229) );
  AND_GATE U127 ( .I1(n30), .I2(n227), .O(n96) );
  AND_GATE U128 ( .I1(n153), .I2(n30), .O(n97) );
  AND_GATE U129 ( .I1(n201), .I2(n100), .O(n98) );
  NOR_GATE U130 ( .I1(n98), .I2(n99), .O(n243) );
  AND_GATE U131 ( .I1(n29), .I2(n241), .O(n99) );
  AND_GATE U132 ( .I1(n154), .I2(n29), .O(n100) );
  AND_GATE U133 ( .I1(n201), .I2(n103), .O(n101) );
  NOR_GATE U134 ( .I1(n101), .I2(n102), .O(n250) );
  AND_GATE U135 ( .I1(n28), .I2(n248), .O(n102) );
  AND_GATE U136 ( .I1(n160), .I2(n28), .O(n103) );
  AND_GATE U137 ( .I1(n201), .I2(n106), .O(n104) );
  NOR_GATE U138 ( .I1(n104), .I2(n105), .O(n257) );
  AND_GATE U139 ( .I1(n27), .I2(n255), .O(n105) );
  AND_GATE U140 ( .I1(n155), .I2(n27), .O(n106) );
  AND_GATE U141 ( .I1(n201), .I2(n109), .O(n107) );
  NOR_GATE U142 ( .I1(n107), .I2(n108), .O(n263) );
  AND_GATE U143 ( .I1(n16), .I2(n261), .O(n108) );
  AND_GATE U144 ( .I1(n146), .I2(n16), .O(n109) );
  NAND_GATE U145 ( .I1(n201), .I2(n112), .O(n110) );
  AND_GATE U146 ( .I1(n110), .I2(n111), .O(n271) );
  OR_GATE U147 ( .I1(n273), .I2(n269), .O(n111) );
  AND_GATE U148 ( .I1(n270), .I2(n274), .O(n112) );
  OR_GATE U149 ( .I1(n302), .I2(n113), .O(n300) );
  AND_GATE U150 ( .I1(n303), .I2(n304), .O(n113) );
  OR_GATE U151 ( .I1(n218), .I2(n114), .O(n217) );
  OR_GATE U152 ( .I1(n214), .I2(n18), .O(n114) );
  OR_GATE U153 ( .I1(n31), .I2(n220), .O(n115) );
  OR_GATE U154 ( .I1(n30), .I2(n227), .O(n116) );
  OR_GATE U155 ( .I1(n29), .I2(n241), .O(n117) );
  OR_GATE U156 ( .I1(n28), .I2(n248), .O(n118) );
  OR_GATE U157 ( .I1(n27), .I2(n255), .O(n119) );
  OR_GATE U158 ( .I1(n16), .I2(n261), .O(n120) );
  INV_GATE U159 ( .I1(n269), .O(n121) );
  NAND_GATE U160 ( .I1(n122), .I2(n275), .O(n272) );
  NOR_GATE U161 ( .I1(n121), .I2(n274), .O(n122) );
  NAND5_GATE U162 ( .I1(n182), .I2(n287), .I3(n156), .I4(n286), .I5(n147), .O(
        n186) );
  NAND3_GATE U163 ( .I1(n366), .I2(n367), .I3(n363), .O(n362) );
  NAND3_GATE U164 ( .I1(B[48]), .I2(A[48]), .I3(n268), .O(n266) );
  NAND4_GATE U165 ( .I1(n352), .I2(n351), .I3(n396), .I4(n290), .O(n371) );
  NAND3_GATE U166 ( .I1(n219), .I2(n138), .I3(n137), .O(n214) );
  NAND_GATE U167 ( .I1(B[31]), .I2(A[31]), .O(n123) );
  AND_GATE U168 ( .I1(n150), .I2(A[31]), .O(n124) );
  INV_GATE U169 ( .I1(n303), .O(n125) );
  NAND_GATE U170 ( .I1(n126), .I2(n304), .O(n301) );
  NOR_GATE U171 ( .I1(n125), .I2(n166), .O(n126) );
  AND_GATE U172 ( .I1(B[32]), .I2(A[32]), .O(n127) );
  AND3_GATE U173 ( .I1(n320), .I2(n283), .I3(n321), .O(n128) );
  NAND_GATE U174 ( .I1(n266), .I2(n132), .O(n129) );
  AND_GATE U175 ( .I1(n129), .I2(n130), .O(n255) );
  OR_GATE U176 ( .I1(n131), .I2(n262), .O(n130) );
  INV_GATE U177 ( .I1(n260), .O(n131) );
  AND_GATE U178 ( .I1(n267), .I2(n260), .O(n132) );
  AND_GATE U179 ( .I1(n133), .I2(n134), .O(n181) );
  OR_GATE U180 ( .I1(n135), .I2(n198), .O(n134) );
  INV_GATE U181 ( .I1(n182), .O(n135) );
  AND_GATE U182 ( .I1(n200), .I2(n182), .O(n136) );
  NAND_GATE U183 ( .I1(n227), .I2(n140), .O(n137) );
  OR_GATE U184 ( .I1(n139), .I2(n226), .O(n138) );
  INV_GATE U185 ( .I1(n221), .O(n139) );
  AND_GATE U186 ( .I1(n228), .I2(n221), .O(n140) );
  AND_GATE U187 ( .I1(n378), .I2(n21), .O(n375) );
  AND3_GATE U188 ( .I1(n389), .I2(n364), .I3(n390), .O(n141) );
  OR_GATE U189 ( .I1(n73), .I2(n196), .O(n193) );
  AND4_GATE U190 ( .I1(n360), .I2(n366), .I3(n367), .I4(n372), .O(n142) );
  INV_GATE U191 ( .I1(n142), .O(n285) );
  AND_GATE U192 ( .I1(B[31]), .I2(A[31]), .O(n143) );
  AND_GATE U193 ( .I1(n142), .I2(n173), .O(n144) );
  AND_GATE U194 ( .I1(n173), .I2(n147), .O(n145) );
  AND_GATE U195 ( .I1(n270), .I2(n268), .O(n146) );
  AND4_GATE U196 ( .I1(n292), .I2(n190), .I3(n293), .I4(n294), .O(n147) );
  NAND_GATE U197 ( .I1(n190), .I2(n189), .O(n171) );
  OR_GATE U198 ( .I1(n297), .I2(n148), .O(n296) );
  INV_GATE U199 ( .I1(n292), .O(n148) );
  AND_GATE U200 ( .I1(n294), .I2(n293), .O(n149) );
  AND4_GATE U201 ( .I1(n322), .I2(n328), .I3(n329), .I4(n333), .O(n150) );
  AND_GATE U202 ( .I1(n157), .I2(n208), .O(n151) );
  AND_GATE U203 ( .I1(n158), .I2(n221), .O(n152) );
  AND_GATE U204 ( .I1(n159), .I2(n235), .O(n153) );
  AND_GATE U205 ( .I1(n160), .I2(n249), .O(n154) );
  AND_GATE U206 ( .I1(n146), .I2(n262), .O(n155) );
  AND_GATE U207 ( .I1(n151), .I2(n200), .O(n156) );
  AND_GATE U208 ( .I1(n152), .I2(n215), .O(n157) );
  AND_GATE U209 ( .I1(n153), .I2(n228), .O(n158) );
  AND_GATE U210 ( .I1(n154), .I2(n242), .O(n159) );
  AND_GATE U211 ( .I1(n155), .I2(n256), .O(n160) );
  NOR_GATE U212 ( .I1(1'b0), .I2(n419), .O(SUM[31]) );
  NAND_GATE U213 ( .I1(n283), .I2(n165), .O(n162) );
  NAND_GATE U214 ( .I1(n162), .I2(n163), .O(n280) );
  OR_GATE U215 ( .I1(n164), .I2(n172), .O(n163) );
  INV_GATE U216 ( .I1(n171), .O(n164) );
  AND_GATE U217 ( .I1(n284), .I2(n171), .O(n165) );
  INV_GATE U218 ( .I1(n302), .O(n166) );
  NAND_GATE U219 ( .I1(n359), .I2(n170), .O(n167) );
  NAND_GATE U220 ( .I1(n167), .I2(n168), .O(n287) );
  OR_GATE U221 ( .I1(n169), .I2(n285), .O(n168) );
  INV_GATE U222 ( .I1(n150), .O(n169) );
  AND_GATE U223 ( .I1(n360), .I2(n150), .O(n170) );
  AND_GATE U224 ( .I1(n147), .I2(n190), .O(n172) );
  OR_GATE U225 ( .I1(n115), .I2(n224), .O(n223) );
  OR_GATE U226 ( .I1(n116), .I2(n231), .O(n230) );
  OR_GATE U227 ( .I1(n117), .I2(n245), .O(n244) );
  OR_GATE U228 ( .I1(n118), .I2(n252), .O(n251) );
  OR_GATE U229 ( .I1(n119), .I2(n259), .O(n258) );
  OR_GATE U230 ( .I1(n120), .I2(n265), .O(n264) );
  AND4_GATE U231 ( .I1(n399), .I2(n352), .I3(n396), .I4(n351), .O(n173) );
  AND_GATE U233 ( .I1(n174), .I2(n175), .O(SUM[61]) );
  NAND_GATE U234 ( .I1(B[61]), .I2(n176), .O(n175) );
  OR_GATE U235 ( .I1(B[61]), .I2(n176), .O(n174) );
  NAND5_GATE U236 ( .I1(n177), .I2(n178), .I3(n179), .I4(n180), .I5(n181), .O(
        n176) );
  NAND5_GATE U237 ( .I1(n150), .I2(n143), .I3(n183), .I4(n184), .I5(n145), .O(
        n180) );
  AND_GATE U238 ( .I1(n185), .I2(n186), .O(n179) );
  NAND3_GATE U239 ( .I1(n189), .I2(n190), .I3(n184), .O(n178) );
  INV_GATE U240 ( .I1(n187), .O(n184) );
  OR_GATE U241 ( .I1(n187), .I2(n191), .O(n177) );
  NAND_GATE U242 ( .I1(n156), .I2(n182), .O(n187) );
  AND_GATE U243 ( .I1(n192), .I2(n193), .O(SUM[60]) );
  NAND_GATE U244 ( .I1(n199), .I2(n200), .O(n197) );
  AND_GATE U245 ( .I1(n156), .I2(n201), .O(n196) );
  INV_GATE U246 ( .I1(n194), .O(n195) );
  NAND_GATE U247 ( .I1(n185), .I2(n182), .O(n194) );
  OR_GATE U248 ( .I1(A[60]), .I2(B[60]), .O(n182) );
  NAND_GATE U249 ( .I1(B[60]), .I2(A[60]), .O(n185) );
  AND_GATE U250 ( .I1(n202), .I2(n203), .O(SUM[59]) );
  NAND_GATE U251 ( .I1(n205), .I2(n206), .O(n199) );
  NAND_GATE U252 ( .I1(n207), .I2(n208), .O(n205) );
  AND_GATE U253 ( .I1(n151), .I2(n201), .O(n204) );
  NAND_GATE U254 ( .I1(B[59]), .I2(A[59]), .O(n198) );
  OR_GATE U255 ( .I1(A[59]), .I2(B[59]), .O(n200) );
  AND_GATE U256 ( .I1(n209), .I2(n210), .O(SUM[58]) );
  NAND_GATE U257 ( .I1(n212), .I2(n213), .O(n207) );
  NAND_GATE U258 ( .I1(n214), .I2(n215), .O(n212) );
  AND_GATE U259 ( .I1(n157), .I2(n201), .O(n211) );
  NAND_GATE U260 ( .I1(B[58]), .I2(A[58]), .O(n206) );
  OR_GATE U261 ( .I1(A[58]), .I2(B[58]), .O(n208) );
  AND_GATE U262 ( .I1(n216), .I2(n217), .O(SUM[57]) );
  AND_GATE U263 ( .I1(n152), .I2(n201), .O(n218) );
  NAND_GATE U264 ( .I1(B[57]), .I2(A[57]), .O(n213) );
  OR_GATE U265 ( .I1(A[57]), .I2(B[57]), .O(n215) );
  AND_GATE U266 ( .I1(n222), .I2(n223), .O(SUM[56]) );
  NAND_GATE U267 ( .I1(n225), .I2(n226), .O(n220) );
  NAND_GATE U268 ( .I1(n227), .I2(n228), .O(n225) );
  AND_GATE U269 ( .I1(n158), .I2(n201), .O(n224) );
  NAND_GATE U270 ( .I1(B[56]), .I2(A[56]), .O(n219) );
  OR_GATE U271 ( .I1(A[56]), .I2(B[56]), .O(n221) );
  AND_GATE U272 ( .I1(n229), .I2(n230), .O(SUM[55]) );
  NAND_GATE U273 ( .I1(n232), .I2(n233), .O(n227) );
  NAND_GATE U274 ( .I1(n234), .I2(n235), .O(n232) );
  AND_GATE U275 ( .I1(n153), .I2(n201), .O(n231) );
  NAND_GATE U276 ( .I1(B[55]), .I2(A[55]), .O(n226) );
  OR_GATE U277 ( .I1(A[55]), .I2(B[55]), .O(n228) );
  AND_GATE U278 ( .I1(n236), .I2(n237), .O(SUM[54]) );
  NAND_GATE U279 ( .I1(n239), .I2(n240), .O(n234) );
  AND_GATE U280 ( .I1(n159), .I2(n201), .O(n238) );
  NAND_GATE U281 ( .I1(B[54]), .I2(A[54]), .O(n233) );
  OR_GATE U282 ( .I1(A[54]), .I2(B[54]), .O(n235) );
  AND_GATE U283 ( .I1(n243), .I2(n244), .O(SUM[53]) );
  NAND_GATE U284 ( .I1(n246), .I2(n247), .O(n241) );
  NAND_GATE U285 ( .I1(n248), .I2(n249), .O(n246) );
  AND_GATE U286 ( .I1(n154), .I2(n201), .O(n245) );
  NAND_GATE U287 ( .I1(B[53]), .I2(A[53]), .O(n240) );
  OR_GATE U288 ( .I1(A[53]), .I2(B[53]), .O(n242) );
  AND_GATE U289 ( .I1(n250), .I2(n251), .O(SUM[52]) );
  NAND_GATE U290 ( .I1(n253), .I2(n254), .O(n248) );
  NAND_GATE U291 ( .I1(n255), .I2(n256), .O(n253) );
  AND_GATE U292 ( .I1(n160), .I2(n201), .O(n252) );
  NAND_GATE U293 ( .I1(B[52]), .I2(A[52]), .O(n247) );
  OR_GATE U294 ( .I1(A[52]), .I2(B[52]), .O(n249) );
  AND_GATE U295 ( .I1(n257), .I2(n258), .O(SUM[51]) );
  AND_GATE U296 ( .I1(n155), .I2(n201), .O(n259) );
  NAND_GATE U297 ( .I1(B[51]), .I2(A[51]), .O(n254) );
  OR_GATE U298 ( .I1(A[51]), .I2(B[51]), .O(n256) );
  AND_GATE U299 ( .I1(n263), .I2(n264), .O(SUM[50]) );
  NAND_GATE U300 ( .I1(n266), .I2(n267), .O(n261) );
  AND_GATE U301 ( .I1(n146), .I2(n201), .O(n265) );
  NAND_GATE U302 ( .I1(B[50]), .I2(A[50]), .O(n260) );
  OR_GATE U303 ( .I1(A[50]), .I2(B[50]), .O(n262) );
  AND_GATE U304 ( .I1(n271), .I2(n272), .O(SUM[49]) );
  NAND_GATE U305 ( .I1(n201), .I2(n270), .O(n275) );
  INV_GATE U306 ( .I1(n273), .O(n274) );
  NAND_GATE U307 ( .I1(n268), .I2(n267), .O(n273) );
  NAND_GATE U308 ( .I1(B[49]), .I2(A[49]), .O(n267) );
  OR_GATE U309 ( .I1(A[49]), .I2(B[49]), .O(n268) );
  AND_GATE U310 ( .I1(n276), .I2(n277), .O(SUM[48]) );
  NAND_GATE U311 ( .I1(n49), .I2(n278), .O(n277) );
  NAND_GATE U312 ( .I1(n279), .I2(n201), .O(n276) );
  NAND3_GATE U313 ( .I1(n280), .I2(n188), .I3(n281), .O(n201) );
  NAND3_GATE U314 ( .I1(n145), .I2(n183), .I3(n282), .O(n281) );
  AND_GATE U315 ( .I1(n124), .I2(B[31]), .O(n282) );
  NAND3_GATE U316 ( .I1(n283), .I2(n284), .I3(n285), .O(n183) );
  NAND3_GATE U317 ( .I1(n147), .I2(n286), .I3(n287), .O(n188) );
  NAND3_GATE U318 ( .I1(n288), .I2(n371), .I3(n289), .O(n286) );
  NAND_GATE U319 ( .I1(n147), .I2(n291), .O(n191) );
  NAND_GATE U320 ( .I1(n284), .I2(n283), .O(n291) );
  NAND_GATE U321 ( .I1(n295), .I2(n296), .O(n189) );
  AND_GATE U322 ( .I1(n298), .I2(n299), .O(n295) );
  INV_GATE U323 ( .I1(n278), .O(n279) );
  NAND_GATE U324 ( .I1(n270), .I2(n269), .O(n278) );
  NAND_GATE U325 ( .I1(B[48]), .I2(A[48]), .O(n269) );
  OR_GATE U326 ( .I1(A[48]), .I2(B[48]), .O(n270) );
  AND_GATE U327 ( .I1(n300), .I2(n301), .O(SUM[47]) );
  NAND3_GATE U328 ( .I1(n149), .I2(n292), .I3(n305), .O(n304) );
  NAND_GATE U329 ( .I1(n306), .I2(n292), .O(n303) );
  NAND_GATE U330 ( .I1(n307), .I2(n299), .O(n306) );
  NAND_GATE U331 ( .I1(n298), .I2(n190), .O(n302) );
  OR_GATE U332 ( .I1(A[47]), .I2(B[47]), .O(n190) );
  NAND_GATE U333 ( .I1(B[47]), .I2(A[47]), .O(n298) );
  AND_GATE U334 ( .I1(n308), .I2(n309), .O(SUM[46]) );
  NAND_GATE U335 ( .I1(n59), .I2(n311), .O(n309) );
  NAND_GATE U336 ( .I1(n149), .I2(n305), .O(n311) );
  NAND_GATE U337 ( .I1(n312), .I2(n293), .O(n307) );
  NAND_GATE U338 ( .I1(n284), .I2(n297), .O(n312) );
  NAND_GATE U339 ( .I1(n292), .I2(n299), .O(n310) );
  NAND_GATE U340 ( .I1(B[46]), .I2(A[46]), .O(n299) );
  OR_GATE U341 ( .I1(A[46]), .I2(B[46]), .O(n292) );
  AND_GATE U342 ( .I1(n313), .I2(n314), .O(SUM[45]) );
  NAND_GATE U343 ( .I1(n305), .I2(n294), .O(n315) );
  NAND_GATE U344 ( .I1(B[45]), .I2(A[45]), .O(n297) );
  OR_GATE U345 ( .I1(A[45]), .I2(B[45]), .O(n293) );
  AND_GATE U346 ( .I1(n316), .I2(n317), .O(SUM[44]) );
  NAND_GATE U347 ( .I1(n128), .I2(n318), .O(n317) );
  NAND_GATE U348 ( .I1(n319), .I2(n305), .O(n316) );
  NAND3_GATE U349 ( .I1(n320), .I2(n283), .I3(n321), .O(n305) );
  NAND3_GATE U350 ( .I1(n150), .I2(n143), .I3(n144), .O(n321) );
  NAND_GATE U351 ( .I1(n326), .I2(n327), .O(n325) );
  AND_GATE U352 ( .I1(n328), .I2(n329), .O(n324) );
  AND_GATE U353 ( .I1(n330), .I2(n331), .O(n323) );
  NAND_GATE U354 ( .I1(n332), .I2(n150), .O(n320) );
  INV_GATE U355 ( .I1(n318), .O(n319) );
  NAND_GATE U356 ( .I1(n294), .I2(n284), .O(n318) );
  NAND_GATE U357 ( .I1(B[44]), .I2(A[44]), .O(n284) );
  OR_GATE U358 ( .I1(A[44]), .I2(B[44]), .O(n294) );
  AND_GATE U359 ( .I1(n334), .I2(n335), .O(SUM[43]) );
  NAND_GATE U360 ( .I1(n24), .I2(n336), .O(n334) );
  NAND_GATE U361 ( .I1(n337), .I2(n338), .O(n336) );
  NAND3_GATE U362 ( .I1(n328), .I2(n329), .I3(n339), .O(n338) );
  NAND_GATE U363 ( .I1(n340), .I2(n328), .O(n337) );
  NAND_GATE U364 ( .I1(n327), .I2(n331), .O(n340) );
  OR_GATE U365 ( .I1(A[43]), .I2(B[43]), .O(n322) );
  NAND_GATE U366 ( .I1(B[43]), .I2(A[43]), .O(n330) );
  AND_GATE U367 ( .I1(n341), .I2(n342), .O(SUM[42]) );
  NAND_GATE U368 ( .I1(n339), .I2(n329), .O(n343) );
  NAND_GATE U369 ( .I1(B[42]), .I2(A[42]), .O(n331) );
  OR_GATE U370 ( .I1(A[42]), .I2(B[42]), .O(n328) );
  AND_GATE U371 ( .I1(n344), .I2(n345), .O(SUM[41]) );
  NAND_GATE U372 ( .I1(n25), .I2(n339), .O(n344) );
  NAND3_GATE U373 ( .I1(n346), .I2(n326), .I3(n347), .O(n339) );
  NAND3_GATE U374 ( .I1(n143), .I2(n333), .I3(n144), .O(n347) );
  NAND_GATE U375 ( .I1(n332), .I2(n333), .O(n346) );
  NAND3_GATE U376 ( .I1(n348), .I2(n288), .I3(n349), .O(n332) );
  NAND4_GATE U377 ( .I1(n142), .I2(n396), .I3(n350), .I4(n290), .O(n349) );
  AND_GATE U378 ( .I1(n351), .I2(n352), .O(n350) );
  NAND_GATE U379 ( .I1(n142), .I2(n353), .O(n348) );
  NAND_GATE U380 ( .I1(B[41]), .I2(A[41]), .O(n327) );
  OR_GATE U381 ( .I1(A[41]), .I2(B[41]), .O(n329) );
  AND_GATE U382 ( .I1(n354), .I2(n355), .O(SUM[40]) );
  NAND_GATE U383 ( .I1(n26), .I2(n356), .O(n354) );
  NAND3_GATE U384 ( .I1(n357), .I2(n288), .I3(n358), .O(n356) );
  NAND_GATE U385 ( .I1(n144), .I2(n143), .O(n358) );
  NAND_GATE U386 ( .I1(n359), .I2(n360), .O(n288) );
  NAND_GATE U387 ( .I1(n361), .I2(n362), .O(n359) );
  NAND_GATE U388 ( .I1(n364), .I2(n365), .O(n363) );
  AND_GATE U389 ( .I1(n368), .I2(n369), .O(n361) );
  NAND_GATE U390 ( .I1(n142), .I2(n370), .O(n357) );
  NAND_GATE U391 ( .I1(n289), .I2(n371), .O(n370) );
  OR_GATE U392 ( .I1(A[40]), .I2(B[40]), .O(n333) );
  NAND_GATE U393 ( .I1(B[40]), .I2(A[40]), .O(n326) );
  AND_GATE U394 ( .I1(n373), .I2(n374), .O(SUM[39]) );
  NAND_GATE U395 ( .I1(n375), .I2(n376), .O(n374) );
  NAND3_GATE U396 ( .I1(n366), .I2(n367), .I3(n379), .O(n378) );
  NAND_GATE U397 ( .I1(n380), .I2(n366), .O(n377) );
  INV_GATE U398 ( .I1(n365), .O(n380) );
  NAND_GATE U399 ( .I1(n368), .I2(n360), .O(n376) );
  OR_GATE U400 ( .I1(A[39]), .I2(B[39]), .O(n360) );
  NAND_GATE U401 ( .I1(B[39]), .I2(A[39]), .O(n368) );
  AND_GATE U402 ( .I1(n381), .I2(n382), .O(SUM[38]) );
  NAND_GATE U403 ( .I1(n54), .I2(n384), .O(n382) );
  NAND_GATE U404 ( .I1(n367), .I2(n379), .O(n384) );
  NAND_GATE U405 ( .I1(n366), .I2(n369), .O(n383) );
  NAND_GATE U406 ( .I1(B[38]), .I2(A[38]), .O(n369) );
  OR_GATE U407 ( .I1(A[38]), .I2(B[38]), .O(n366) );
  AND_GATE U408 ( .I1(n385), .I2(n386), .O(SUM[37]) );
  NAND_GATE U409 ( .I1(n141), .I2(n387), .O(n386) );
  NAND_GATE U410 ( .I1(n388), .I2(n379), .O(n385) );
  NAND3_GATE U411 ( .I1(n389), .I2(n364), .I3(n390), .O(n379) );
  NAND3_GATE U412 ( .I1(n173), .I2(n372), .I3(n143), .O(n390) );
  NAND_GATE U413 ( .I1(n370), .I2(n372), .O(n389) );
  INV_GATE U414 ( .I1(n387), .O(n388) );
  NAND_GATE U415 ( .I1(n367), .I2(n365), .O(n387) );
  NAND_GATE U416 ( .I1(B[37]), .I2(A[37]), .O(n365) );
  OR_GATE U417 ( .I1(A[37]), .I2(B[37]), .O(n367) );
  AND_GATE U418 ( .I1(n391), .I2(n392), .O(SUM[36]) );
  NAND_GATE U419 ( .I1(n394), .I2(n395), .O(n290) );
  OR_GATE U420 ( .I1(A[34]), .I2(B[34]), .O(n396) );
  INV_GATE U421 ( .I1(n353), .O(n289) );
  NAND_GATE U422 ( .I1(n397), .I2(n398), .O(n353) );
  NAND3_GATE U423 ( .I1(B[34]), .I2(n351), .I3(A[34]), .O(n397) );
  AND_GATE U424 ( .I1(n173), .I2(n143), .O(n393) );
  OR_GATE U425 ( .I1(A[36]), .I2(B[36]), .O(n372) );
  NAND_GATE U426 ( .I1(B[36]), .I2(A[36]), .O(n364) );
  AND_GATE U427 ( .I1(n400), .I2(n401), .O(SUM[35]) );
  NAND_GATE U428 ( .I1(n396), .I2(n404), .O(n402) );
  NAND_GATE U429 ( .I1(B[35]), .I2(A[35]), .O(n398) );
  OR_GATE U430 ( .I1(A[35]), .I2(B[35]), .O(n351) );
  AND_GATE U431 ( .I1(n405), .I2(n406), .O(SUM[34]) );
  NAND_GATE U432 ( .I1(n23), .I2(n404), .O(n405) );
  NAND3_GATE U433 ( .I1(n395), .I2(n407), .I3(n408), .O(n404) );
  NAND3_GATE U434 ( .I1(n399), .I2(n352), .I3(n143), .O(n408) );
  NAND_GATE U435 ( .I1(n127), .I2(n352), .O(n407) );
  NAND_GATE U436 ( .I1(B[34]), .I2(A[34]), .O(n403) );
  AND_GATE U437 ( .I1(n409), .I2(n410), .O(SUM[33]) );
  NAND_GATE U438 ( .I1(n143), .I2(n399), .O(n413) );
  INV_GATE U439 ( .I1(n411), .O(n412) );
  NAND_GATE U440 ( .I1(n352), .I2(n395), .O(n411) );
  NAND_GATE U441 ( .I1(B[33]), .I2(A[33]), .O(n395) );
  OR_GATE U442 ( .I1(A[33]), .I2(B[33]), .O(n352) );
  AND_GATE U443 ( .I1(n414), .I2(n415), .O(SUM[32]) );
  NAND_GATE U444 ( .I1(n123), .I2(n416), .O(n415) );
  NAND_GATE U445 ( .I1(n417), .I2(n143), .O(n414) );
  INV_GATE U446 ( .I1(n416), .O(n417) );
  NAND_GATE U447 ( .I1(n399), .I2(n394), .O(n416) );
  NAND_GATE U448 ( .I1(B[32]), .I2(A[32]), .O(n394) );
  OR_GATE U449 ( .I1(A[32]), .I2(B[32]), .O(n399) );
  NAND_GATE U450 ( .I1(n418), .I2(n123), .O(n419) );
  OR_GATE U451 ( .I1(A[31]), .I2(B[31]), .O(n418) );
endmodule


module alu_DW01_add_10 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455;
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND_GATE U2 ( .I1(n209), .I2(n4), .O(n1) );
  NAND_GATE U3 ( .I1(n1), .I2(n2), .O(n443) );
  OR_GATE U4 ( .I1(n3), .I2(n43), .O(n2) );
  INV_GATE U5 ( .I1(n42), .O(n3) );
  AND_GATE U6 ( .I1(n210), .I2(n42), .O(n4) );
  OR_GATE U7 ( .I1(n215), .I2(n5), .O(n202) );
  INV_GATE U8 ( .I1(n187), .O(n5) );
  NAND3_GATE U9 ( .I1(n322), .I2(n321), .I3(n320), .O(n6) );
  NAND_GATE U10 ( .I1(n238), .I2(n10), .O(n7) );
  AND_GATE U11 ( .I1(n7), .I2(n8), .O(n226) );
  OR_GATE U12 ( .I1(n9), .I2(n234), .O(n8) );
  INV_GATE U13 ( .I1(n232), .O(n9) );
  AND_GATE U14 ( .I1(n239), .I2(n232), .O(n10) );
  NAND_GATE U15 ( .I1(n240), .I2(n14), .O(n11) );
  NAND_GATE U16 ( .I1(n11), .I2(n12), .O(n121) );
  OR_GATE U17 ( .I1(n13), .I2(n239), .O(n12) );
  INV_GATE U18 ( .I1(n35), .O(n13) );
  AND_GATE U19 ( .I1(n241), .I2(n35), .O(n14) );
  NAND_GATE U20 ( .I1(n281), .I2(n18), .O(n15) );
  AND_GATE U21 ( .I1(n15), .I2(n16), .O(n111) );
  OR_GATE U22 ( .I1(n17), .I2(n280), .O(n16) );
  INV_GATE U23 ( .I1(n114), .O(n17) );
  AND_GATE U24 ( .I1(n282), .I2(n114), .O(n18) );
  AND_GATE U25 ( .I1(n354), .I2(n351), .O(n19) );
  AND_GATE U26 ( .I1(n320), .I2(n328), .O(n20) );
  AND_GATE U27 ( .I1(n327), .I2(n212), .O(n21) );
  AND_GATE U28 ( .I1(n289), .I2(n287), .O(n22) );
  AND_GATE U29 ( .I1(n282), .I2(n280), .O(n23) );
  AND_GATE U30 ( .I1(n275), .I2(n273), .O(n24) );
  AND_GATE U31 ( .I1(n268), .I2(n266), .O(n25) );
  AND_GATE U32 ( .I1(n262), .I2(n260), .O(n26) );
  AND_GATE U33 ( .I1(n255), .I2(n253), .O(n27) );
  AND_GATE U34 ( .I1(n248), .I2(n246), .O(n28) );
  AND_GATE U35 ( .I1(n241), .I2(n239), .O(n29) );
  AND_GATE U36 ( .I1(n227), .I2(n225), .O(n30) );
  AND_GATE U37 ( .I1(n429), .I2(n428), .O(n31) );
  AND_GATE U38 ( .I1(n361), .I2(n355), .O(n32) );
  AND_GATE U39 ( .I1(n322), .I2(n332), .O(n33) );
  AND_GATE U40 ( .I1(n386), .I2(n390), .O(n34) );
  AND_GATE U41 ( .I1(n234), .I2(n232), .O(n35) );
  AND_GATE U42 ( .I1(B[30]), .I2(A[30]), .O(n36) );
  AND_GATE U43 ( .I1(n210), .I2(n312), .O(n37) );
  OR_GATE U44 ( .I1(n36), .I2(n37), .O(n453) );
  AND_GATE U45 ( .I1(n389), .I2(n396), .O(n38) );
  AND_GATE U46 ( .I1(n208), .I2(n41), .O(n39) );
  NOR_GATE U47 ( .I1(n39), .I2(n40), .O(n415) );
  AND_GATE U48 ( .I1(n38), .I2(n385), .O(n40) );
  AND_GATE U49 ( .I1(n207), .I2(n38), .O(n41) );
  OR_GATE U50 ( .I1(n445), .I2(n442), .O(n42) );
  AND_GATE U51 ( .I1(n429), .I2(n446), .O(n43) );
  OR_GATE U52 ( .I1(n38), .I2(n385), .O(n44) );
  NAND_GATE U53 ( .I1(n45), .I2(n447), .O(n444) );
  NOR_GATE U54 ( .I1(n441), .I2(n446), .O(n45) );
  OR_GATE U55 ( .I1(n44), .I2(n417), .O(n416) );
  NAND_GATE U56 ( .I1(n226), .I2(n48), .O(n46) );
  NAND_GATE U57 ( .I1(n46), .I2(n47), .O(n126) );
  OR_GATE U58 ( .I1(n222), .I2(n225), .O(n47) );
  AND_GATE U59 ( .I1(n227), .I2(n127), .O(n48) );
  NAND_GATE U60 ( .I1(n224), .I2(n49), .O(n118) );
  AND_GATE U61 ( .I1(n225), .I2(n222), .O(n49) );
  AND_GATE U62 ( .I1(n345), .I2(n332), .O(n50) );
  NAND_GATE U63 ( .I1(n50), .I2(n347), .O(n76) );
  NAND_GATE U64 ( .I1(n326), .I2(n53), .O(n51) );
  NAND_GATE U65 ( .I1(n51), .I2(n52), .O(n64) );
  OR_GATE U66 ( .I1(n345), .I2(n332), .O(n52) );
  AND_GATE U67 ( .I1(n322), .I2(n65), .O(n53) );
  AND_GATE U68 ( .I1(n339), .I2(n56), .O(n54) );
  NOR_GATE U69 ( .I1(n54), .I2(n55), .O(n340) );
  AND_GATE U70 ( .I1(n20), .I2(n338), .O(n55) );
  AND_GATE U71 ( .I1(n172), .I2(n20), .O(n56) );
  OR_GATE U72 ( .I1(n342), .I2(n57), .O(n341) );
  OR_GATE U73 ( .I1(n338), .I2(n20), .O(n57) );
  NAND_GATE U74 ( .I1(n434), .I2(n60), .O(n58) );
  AND_GATE U75 ( .I1(n58), .I2(n59), .O(n430) );
  OR_GATE U76 ( .I1(n432), .I2(n426), .O(n59) );
  AND_GATE U77 ( .I1(n419), .I2(n61), .O(n60) );
  INV_GATE U78 ( .I1(n432), .O(n61) );
  AND_GATE U79 ( .I1(n432), .I2(n426), .O(n62) );
  AND_GATE U80 ( .I1(n339), .I2(n66), .O(n63) );
  NOR_GATE U81 ( .I1(n63), .I2(n64), .O(n343) );
  INV_GATE U82 ( .I1(n345), .O(n65) );
  AND_GATE U83 ( .I1(n171), .I2(n65), .O(n66) );
  AND_GATE U84 ( .I1(n339), .I2(n69), .O(n67) );
  NOR_GATE U85 ( .I1(n67), .I2(n68), .O(n348) );
  AND_GATE U86 ( .I1(n33), .I2(n326), .O(n68) );
  AND_GATE U87 ( .I1(n170), .I2(n33), .O(n69) );
  AND_GATE U88 ( .I1(n339), .I2(n72), .O(n70) );
  NOR_GATE U89 ( .I1(n70), .I2(n71), .O(n370) );
  AND_GATE U90 ( .I1(n32), .I2(n369), .O(n71) );
  AND_GATE U91 ( .I1(n174), .I2(n32), .O(n72) );
  NAND_GATE U92 ( .I1(n339), .I2(n75), .O(n73) );
  AND_GATE U93 ( .I1(n73), .I2(n74), .O(n374) );
  OR_GATE U94 ( .I1(n376), .I2(n360), .O(n74) );
  AND_GATE U95 ( .I1(n363), .I2(n377), .O(n75) );
  OR_GATE U96 ( .I1(n346), .I2(n76), .O(n344) );
  OR_GATE U97 ( .I1(n33), .I2(n326), .O(n77) );
  OR_GATE U98 ( .I1(n32), .I2(n369), .O(n78) );
  INV_GATE U99 ( .I1(n360), .O(n79) );
  NAND_GATE U100 ( .I1(n80), .I2(n378), .O(n375) );
  NOR_GATE U101 ( .I1(n79), .I2(n377), .O(n80) );
  NAND_GATE U102 ( .I1(n403), .I2(n83), .O(n81) );
  AND_GATE U103 ( .I1(n81), .I2(n82), .O(n405) );
  OR_GATE U104 ( .I1(n407), .I2(n394), .O(n82) );
  AND_GATE U105 ( .I1(n388), .I2(n84), .O(n83) );
  INV_GATE U106 ( .I1(n407), .O(n84) );
  AND_GATE U107 ( .I1(n394), .I2(n407), .O(n85) );
  NAND_GATE U108 ( .I1(n226), .I2(n89), .O(n86) );
  AND_GATE U109 ( .I1(n86), .I2(n87), .O(n200) );
  OR_GATE U110 ( .I1(n88), .I2(n225), .O(n87) );
  INV_GATE U111 ( .I1(n214), .O(n88) );
  AND_GATE U112 ( .I1(n227), .I2(n214), .O(n89) );
  AND_GATE U113 ( .I1(n195), .I2(n310), .O(n90) );
  NAND_GATE U114 ( .I1(n358), .I2(n94), .O(n91) );
  NAND_GATE U115 ( .I1(n91), .I2(n92), .O(n96) );
  OR_GATE U116 ( .I1(n93), .I2(n355), .O(n92) );
  INV_GATE U117 ( .I1(n137), .O(n93) );
  AND_GATE U118 ( .I1(n357), .I2(n137), .O(n94) );
  OR3_GATE U119 ( .I1(n136), .I2(n95), .I3(n96), .O(n213) );
  NOR_GATE U120 ( .I1(n6), .I2(n351), .O(n95) );
  NOR3_GATE U121 ( .I1(n311), .I2(n383), .I3(n384), .O(n97) );
  NAND3_GATE U122 ( .I1(n311), .I2(n187), .I3(n310), .O(n205) );
  NAND5_GATE U123 ( .I1(n98), .I2(n201), .I3(n200), .I4(n202), .I5(n203), .O(
        n196) );
  INV_GATE U124 ( .I1(n198), .O(n98) );
  NAND3_GATE U125 ( .I1(n330), .I2(n100), .I3(n99), .O(n338) );
  AND3_GATE U126 ( .I1(n115), .I2(n104), .I3(n103), .O(n337) );
  NAND4_GATE U127 ( .I1(n307), .I2(n211), .I3(n309), .I4(n215), .O(n228) );
  NAND3_GATE U128 ( .I1(n266), .I2(n112), .I3(n111), .O(n261) );
  AND4_GATE U129 ( .I1(n419), .I2(n420), .I3(n428), .I4(n429), .O(n207) );
  NAND_GATE U130 ( .I1(n326), .I2(n102), .O(n99) );
  OR_GATE U131 ( .I1(n101), .I2(n332), .O(n100) );
  INV_GATE U132 ( .I1(n321), .O(n101) );
  AND_GATE U133 ( .I1(n322), .I2(n321), .O(n102) );
  NAND_GATE U134 ( .I1(n326), .I2(n106), .O(n103) );
  OR_GATE U135 ( .I1(n105), .I2(n332), .O(n104) );
  INV_GATE U136 ( .I1(n117), .O(n105) );
  AND_GATE U137 ( .I1(n322), .I2(n117), .O(n106) );
  OR_GATE U138 ( .I1(n265), .I2(n107), .O(n264) );
  OR_GATE U139 ( .I1(n261), .I2(n26), .O(n107) );
  AND_GATE U140 ( .I1(n228), .I2(n110), .O(n108) );
  NOR_GATE U141 ( .I1(n108), .I2(n109), .O(n263) );
  AND_GATE U142 ( .I1(n26), .I2(n261), .O(n109) );
  AND_GATE U143 ( .I1(n184), .I2(n26), .O(n110) );
  OR_GATE U144 ( .I1(n113), .I2(n273), .O(n112) );
  INV_GATE U145 ( .I1(n268), .O(n113) );
  AND_GATE U146 ( .I1(n275), .I2(n268), .O(n114) );
  OR_GATE U147 ( .I1(n116), .I2(n330), .O(n115) );
  INV_GATE U148 ( .I1(n320), .O(n116) );
  AND_GATE U149 ( .I1(n321), .I2(n320), .O(n117) );
  OR_GATE U150 ( .I1(n223), .I2(n118), .O(n221) );
  OR_GATE U151 ( .I1(n231), .I2(n119), .O(n230) );
  OR_GATE U152 ( .I1(n226), .I2(n30), .O(n119) );
  AND_GATE U153 ( .I1(n228), .I2(n122), .O(n120) );
  NOR_GATE U154 ( .I1(n120), .I2(n121), .O(n235) );
  AND_GATE U155 ( .I1(n180), .I2(n35), .O(n122) );
  NAND_GATE U156 ( .I1(n208), .I2(n31), .O(n440) );
  AND3_GATE U157 ( .I1(n421), .I2(n439), .I3(n440), .O(n123) );
  AND_GATE U158 ( .I1(n209), .I2(n210), .O(n124) );
  AND_GATE U159 ( .I1(n228), .I2(n128), .O(n125) );
  NOR_GATE U160 ( .I1(n125), .I2(n126), .O(n220) );
  INV_GATE U161 ( .I1(n222), .O(n127) );
  AND_GATE U162 ( .I1(n178), .I2(n127), .O(n128) );
  AND_GATE U163 ( .I1(n228), .I2(n131), .O(n129) );
  NOR_GATE U164 ( .I1(n129), .I2(n130), .O(n229) );
  AND_GATE U165 ( .I1(n30), .I2(n226), .O(n130) );
  AND_GATE U166 ( .I1(n179), .I2(n30), .O(n131) );
  OR_GATE U167 ( .I1(n35), .I2(n233), .O(n132) );
  NAND_GATE U168 ( .I1(n228), .I2(n135), .O(n133) );
  AND_GATE U169 ( .I1(n133), .I2(n134), .O(n298) );
  OR_GATE U170 ( .I1(n300), .I2(n296), .O(n134) );
  AND_GATE U171 ( .I1(n297), .I2(n301), .O(n135) );
  NAND3_GATE U172 ( .I1(n323), .I2(n324), .I3(n325), .O(n136) );
  AND_GATE U173 ( .I1(n354), .I2(n169), .O(n137) );
  INV_GATE U174 ( .I1(n296), .O(n138) );
  NAND_GATE U175 ( .I1(n139), .I2(n302), .O(n299) );
  NOR_GATE U176 ( .I1(n138), .I2(n301), .O(n139) );
  AND3_GATE U177 ( .I1(n307), .I2(n215), .I3(n308), .O(n140) );
  AND_GATE U178 ( .I1(n228), .I2(n143), .O(n141) );
  NOR_GATE U179 ( .I1(n141), .I2(n142), .O(n242) );
  AND_GATE U180 ( .I1(n29), .I2(n240), .O(n142) );
  AND_GATE U181 ( .I1(n181), .I2(n29), .O(n143) );
  AND_GATE U182 ( .I1(n228), .I2(n146), .O(n144) );
  NOR_GATE U183 ( .I1(n144), .I2(n145), .O(n249) );
  AND_GATE U184 ( .I1(n28), .I2(n247), .O(n145) );
  AND_GATE U185 ( .I1(n182), .I2(n28), .O(n146) );
  AND_GATE U186 ( .I1(n228), .I2(n149), .O(n147) );
  NOR_GATE U187 ( .I1(n147), .I2(n148), .O(n256) );
  AND_GATE U188 ( .I1(n27), .I2(n254), .O(n148) );
  AND_GATE U189 ( .I1(n183), .I2(n27), .O(n149) );
  AND_GATE U190 ( .I1(n228), .I2(n152), .O(n150) );
  NOR_GATE U191 ( .I1(n150), .I2(n151), .O(n269) );
  AND_GATE U192 ( .I1(n25), .I2(n267), .O(n151) );
  AND_GATE U193 ( .I1(n185), .I2(n25), .O(n152) );
  AND_GATE U194 ( .I1(n228), .I2(n155), .O(n153) );
  NOR_GATE U195 ( .I1(n153), .I2(n154), .O(n276) );
  AND_GATE U196 ( .I1(n24), .I2(n274), .O(n154) );
  AND_GATE U197 ( .I1(n186), .I2(n24), .O(n155) );
  OR_GATE U198 ( .I1(n285), .I2(n156), .O(n284) );
  OR_GATE U199 ( .I1(n281), .I2(n23), .O(n156) );
  AND_GATE U200 ( .I1(n228), .I2(n159), .O(n157) );
  NOR_GATE U201 ( .I1(n157), .I2(n158), .O(n290) );
  AND_GATE U202 ( .I1(n22), .I2(n288), .O(n158) );
  AND_GATE U203 ( .I1(n175), .I2(n22), .O(n159) );
  OR_GATE U204 ( .I1(n29), .I2(n240), .O(n160) );
  OR_GATE U205 ( .I1(n28), .I2(n247), .O(n161) );
  OR_GATE U206 ( .I1(n27), .I2(n254), .O(n162) );
  OR_GATE U207 ( .I1(n25), .I2(n267), .O(n163) );
  OR_GATE U208 ( .I1(n24), .I2(n274), .O(n164) );
  OR_GATE U209 ( .I1(n22), .I2(n288), .O(n165) );
  NAND3_GATE U210 ( .I1(n166), .I2(n312), .I3(n167), .O(n309) );
  NAND_GATE U211 ( .I1(n210), .I2(n209), .O(n166) );
  NOR_GATE U212 ( .I1(n314), .I2(n427), .O(n167) );
  OR_GATE U213 ( .I1(n77), .I2(n350), .O(n349) );
  OR_GATE U214 ( .I1(n78), .I2(n372), .O(n371) );
  AND3_GATE U215 ( .I1(n396), .I2(n413), .I3(n414), .O(n168) );
  OR_GATE U216 ( .I1(n366), .I2(n19), .O(n365) );
  AND3_GATE U217 ( .I1(n322), .I2(n321), .I3(n320), .O(n169) );
  AND4_GATE U218 ( .I1(n354), .I2(n361), .I3(n362), .I4(n363), .O(n170) );
  AND_GATE U219 ( .I1(n170), .I2(n322), .O(n171) );
  AND_GATE U220 ( .I1(n171), .I2(n321), .O(n172) );
  OR_GATE U221 ( .I1(n360), .I2(n173), .O(n373) );
  INV_GATE U222 ( .I1(n362), .O(n173) );
  AND_GATE U223 ( .I1(n362), .I2(n363), .O(n174) );
  AND_GATE U224 ( .I1(n297), .I2(n295), .O(n175) );
  OR_GATE U225 ( .I1(n296), .I2(n176), .O(n293) );
  INV_GATE U226 ( .I1(n295), .O(n176) );
  AND_GATE U227 ( .I1(n175), .I2(n289), .O(n177) );
  AND_GATE U228 ( .I1(n179), .I2(n227), .O(n178) );
  AND_GATE U229 ( .I1(n180), .I2(n234), .O(n179) );
  AND_GATE U230 ( .I1(n181), .I2(n241), .O(n180) );
  AND_GATE U231 ( .I1(n182), .I2(n248), .O(n181) );
  AND_GATE U232 ( .I1(n183), .I2(n255), .O(n182) );
  AND_GATE U233 ( .I1(n184), .I2(n262), .O(n183) );
  AND_GATE U234 ( .I1(n185), .I2(n268), .O(n184) );
  AND_GATE U235 ( .I1(n186), .I2(n275), .O(n185) );
  AND_GATE U236 ( .I1(n177), .I2(n282), .O(n186) );
  AND_GATE U237 ( .I1(n178), .I2(n214), .O(n187) );
  NOR_GATE U238 ( .I1(1'b0), .I2(n455), .O(SUM[30]) );
  NAND_GATE U239 ( .I1(n209), .I2(n210), .O(n208) );
  AND_GATE U240 ( .I1(n228), .I2(n191), .O(n189) );
  NOR_GATE U241 ( .I1(n189), .I2(n190), .O(n283) );
  AND_GATE U242 ( .I1(n23), .I2(n281), .O(n190) );
  AND_GATE U243 ( .I1(n177), .I2(n23), .O(n191) );
  AND_GATE U244 ( .I1(n207), .I2(n195), .O(n192) );
  AND_GATE U245 ( .I1(n208), .I2(n192), .O(n383) );
  OR_GATE U246 ( .I1(n400), .I2(n34), .O(n399) );
  OR_GATE U247 ( .I1(n335), .I2(n21), .O(n334) );
  OR_GATE U248 ( .I1(n132), .I2(n237), .O(n236) );
  OR_GATE U249 ( .I1(n160), .I2(n244), .O(n243) );
  OR_GATE U250 ( .I1(n161), .I2(n251), .O(n250) );
  AND_GATE U251 ( .I1(n421), .I2(n422), .O(n193) );
  OR_GATE U252 ( .I1(n162), .I2(n258), .O(n257) );
  AND_GATE U253 ( .I1(n423), .I2(n421), .O(n194) );
  OR3_GATE U254 ( .I1(n194), .I2(n193), .I3(n319), .O(n418) );
  OR_GATE U255 ( .I1(n163), .I2(n271), .O(n270) );
  OR_GATE U256 ( .I1(n164), .I2(n278), .O(n277) );
  OR_GATE U257 ( .I1(n165), .I2(n292), .O(n291) );
  AND4_GATE U258 ( .I1(n386), .I2(n387), .I3(n388), .I4(n389), .O(n195) );
  AND_GATE U260 ( .I1(n196), .I2(n197), .O(SUM[61]) );
  NAND_GATE U261 ( .I1(n198), .I2(n199), .O(n197) );
  NAND4_GATE U262 ( .I1(n200), .I2(n201), .I3(n202), .I4(n203), .O(n199) );
  AND3_GATE U263 ( .I1(n204), .I2(n205), .I3(n206), .O(n203) );
  NAND4_GATE U264 ( .I1(n187), .I2(n90), .I3(n207), .I4(n208), .O(n206) );
  NAND3_GATE U265 ( .I1(n187), .I2(n212), .I3(n213), .O(n204) );
  NAND_GATE U266 ( .I1(n216), .I2(n217), .O(n198) );
  NAND_GATE U267 ( .I1(B[61]), .I2(n218), .O(n217) );
  INV_GATE U268 ( .I1(A[61]), .O(n218) );
  NAND_GATE U269 ( .I1(A[61]), .I2(n219), .O(n216) );
  INV_GATE U270 ( .I1(B[61]), .O(n219) );
  AND_GATE U271 ( .I1(n220), .I2(n221), .O(SUM[60]) );
  NAND_GATE U272 ( .I1(n226), .I2(n227), .O(n224) );
  AND_GATE U273 ( .I1(n178), .I2(n228), .O(n223) );
  NAND_GATE U274 ( .I1(n201), .I2(n214), .O(n222) );
  OR_GATE U275 ( .I1(A[60]), .I2(B[60]), .O(n214) );
  NAND_GATE U276 ( .I1(B[60]), .I2(A[60]), .O(n201) );
  AND_GATE U277 ( .I1(n229), .I2(n230), .O(SUM[59]) );
  AND_GATE U278 ( .I1(n179), .I2(n228), .O(n231) );
  NAND_GATE U279 ( .I1(B[59]), .I2(A[59]), .O(n225) );
  OR_GATE U280 ( .I1(A[59]), .I2(B[59]), .O(n227) );
  AND_GATE U281 ( .I1(n235), .I2(n236), .O(SUM[58]) );
  NAND_GATE U282 ( .I1(n238), .I2(n239), .O(n233) );
  NAND_GATE U283 ( .I1(n240), .I2(n241), .O(n238) );
  AND_GATE U284 ( .I1(n180), .I2(n228), .O(n237) );
  NAND_GATE U285 ( .I1(B[58]), .I2(A[58]), .O(n232) );
  OR_GATE U286 ( .I1(A[58]), .I2(B[58]), .O(n234) );
  AND_GATE U287 ( .I1(n242), .I2(n243), .O(SUM[57]) );
  NAND_GATE U288 ( .I1(n245), .I2(n246), .O(n240) );
  NAND_GATE U289 ( .I1(n247), .I2(n248), .O(n245) );
  AND_GATE U290 ( .I1(n181), .I2(n228), .O(n244) );
  NAND_GATE U291 ( .I1(B[57]), .I2(A[57]), .O(n239) );
  OR_GATE U292 ( .I1(A[57]), .I2(B[57]), .O(n241) );
  AND_GATE U293 ( .I1(n249), .I2(n250), .O(SUM[56]) );
  NAND_GATE U294 ( .I1(n252), .I2(n253), .O(n247) );
  NAND_GATE U295 ( .I1(n254), .I2(n255), .O(n252) );
  AND_GATE U296 ( .I1(n182), .I2(n228), .O(n251) );
  NAND_GATE U297 ( .I1(B[56]), .I2(A[56]), .O(n246) );
  OR_GATE U298 ( .I1(A[56]), .I2(B[56]), .O(n248) );
  AND_GATE U299 ( .I1(n256), .I2(n257), .O(SUM[55]) );
  NAND_GATE U300 ( .I1(n259), .I2(n260), .O(n254) );
  NAND_GATE U301 ( .I1(n261), .I2(n262), .O(n259) );
  AND_GATE U302 ( .I1(n183), .I2(n228), .O(n258) );
  NAND_GATE U303 ( .I1(B[55]), .I2(A[55]), .O(n253) );
  OR_GATE U304 ( .I1(A[55]), .I2(B[55]), .O(n255) );
  AND_GATE U305 ( .I1(n263), .I2(n264), .O(SUM[54]) );
  AND_GATE U306 ( .I1(n184), .I2(n228), .O(n265) );
  NAND_GATE U307 ( .I1(B[54]), .I2(A[54]), .O(n260) );
  OR_GATE U308 ( .I1(A[54]), .I2(B[54]), .O(n262) );
  AND_GATE U309 ( .I1(n269), .I2(n270), .O(SUM[53]) );
  NAND_GATE U310 ( .I1(n272), .I2(n273), .O(n267) );
  NAND_GATE U311 ( .I1(n274), .I2(n275), .O(n272) );
  AND_GATE U312 ( .I1(n185), .I2(n228), .O(n271) );
  NAND_GATE U313 ( .I1(B[53]), .I2(A[53]), .O(n266) );
  OR_GATE U314 ( .I1(A[53]), .I2(B[53]), .O(n268) );
  AND_GATE U315 ( .I1(n276), .I2(n277), .O(SUM[52]) );
  NAND_GATE U316 ( .I1(n279), .I2(n280), .O(n274) );
  NAND_GATE U317 ( .I1(n281), .I2(n282), .O(n279) );
  AND_GATE U318 ( .I1(n186), .I2(n228), .O(n278) );
  NAND_GATE U319 ( .I1(B[52]), .I2(A[52]), .O(n273) );
  OR_GATE U320 ( .I1(A[52]), .I2(B[52]), .O(n275) );
  AND_GATE U321 ( .I1(n283), .I2(n284), .O(SUM[51]) );
  NAND_GATE U322 ( .I1(n286), .I2(n287), .O(n281) );
  NAND_GATE U323 ( .I1(n288), .I2(n289), .O(n286) );
  AND_GATE U324 ( .I1(n177), .I2(n228), .O(n285) );
  NAND_GATE U325 ( .I1(B[51]), .I2(A[51]), .O(n280) );
  OR_GATE U326 ( .I1(A[51]), .I2(B[51]), .O(n282) );
  AND_GATE U327 ( .I1(n290), .I2(n291), .O(SUM[50]) );
  NAND_GATE U328 ( .I1(n293), .I2(n294), .O(n288) );
  AND_GATE U329 ( .I1(n175), .I2(n228), .O(n292) );
  NAND_GATE U330 ( .I1(B[50]), .I2(A[50]), .O(n287) );
  OR_GATE U331 ( .I1(A[50]), .I2(B[50]), .O(n289) );
  AND_GATE U332 ( .I1(n298), .I2(n299), .O(SUM[49]) );
  NAND_GATE U333 ( .I1(n228), .I2(n297), .O(n302) );
  INV_GATE U334 ( .I1(n300), .O(n301) );
  NAND_GATE U335 ( .I1(n295), .I2(n294), .O(n300) );
  NAND_GATE U336 ( .I1(B[49]), .I2(A[49]), .O(n294) );
  OR_GATE U337 ( .I1(A[49]), .I2(B[49]), .O(n295) );
  AND_GATE U338 ( .I1(n303), .I2(n304), .O(SUM[48]) );
  NAND_GATE U339 ( .I1(n140), .I2(n305), .O(n304) );
  NAND_GATE U340 ( .I1(n306), .I2(n228), .O(n303) );
  AND_GATE U341 ( .I1(n309), .I2(n211), .O(n308) );
  NAND_GATE U342 ( .I1(n310), .I2(n311), .O(n211) );
  OR_GATE U343 ( .I1(A[30]), .I2(B[30]), .O(n313) );
  NAND_GATE U344 ( .I1(n195), .I2(n310), .O(n314) );
  NAND5_GATE U345 ( .I1(n195), .I2(n310), .I3(n315), .I4(n316), .I5(n317), .O(
        n215) );
  NAND_GATE U346 ( .I1(n318), .I2(n319), .O(n317) );
  NAND_GATE U347 ( .I1(n193), .I2(n318), .O(n316) );
  NAND_GATE U348 ( .I1(n194), .I2(n318), .O(n315) );
  AND5_GATE U349 ( .I1(n320), .I2(n212), .I3(n321), .I4(n322), .I5(n170), .O(
        n310) );
  NAND_GATE U350 ( .I1(n213), .I2(n212), .O(n307) );
  AND_GATE U351 ( .I1(n327), .I2(n328), .O(n325) );
  NAND_GATE U352 ( .I1(n329), .I2(n320), .O(n324) );
  INV_GATE U353 ( .I1(n330), .O(n329) );
  NAND3_GATE U354 ( .I1(n320), .I2(n331), .I3(n321), .O(n323) );
  INV_GATE U355 ( .I1(n332), .O(n331) );
  INV_GATE U356 ( .I1(n305), .O(n306) );
  NAND_GATE U357 ( .I1(n297), .I2(n296), .O(n305) );
  NAND_GATE U358 ( .I1(B[48]), .I2(A[48]), .O(n296) );
  OR_GATE U359 ( .I1(A[48]), .I2(B[48]), .O(n297) );
  AND_GATE U360 ( .I1(n333), .I2(n334), .O(SUM[47]) );
  NAND_GATE U361 ( .I1(n21), .I2(n335), .O(n333) );
  NAND3_GATE U362 ( .I1(n328), .I2(n336), .I3(n337), .O(n335) );
  NAND3_GATE U363 ( .I1(n172), .I2(n320), .I3(n339), .O(n336) );
  OR_GATE U364 ( .I1(A[47]), .I2(B[47]), .O(n212) );
  NAND_GATE U365 ( .I1(B[47]), .I2(A[47]), .O(n327) );
  AND_GATE U366 ( .I1(n340), .I2(n341), .O(SUM[46]) );
  AND_GATE U367 ( .I1(n172), .I2(n339), .O(n342) );
  NAND_GATE U368 ( .I1(B[46]), .I2(A[46]), .O(n328) );
  OR_GATE U369 ( .I1(A[46]), .I2(B[46]), .O(n320) );
  AND_GATE U370 ( .I1(n343), .I2(n344), .O(SUM[45]) );
  NAND_GATE U371 ( .I1(n326), .I2(n322), .O(n347) );
  AND_GATE U372 ( .I1(n171), .I2(n339), .O(n346) );
  NAND_GATE U373 ( .I1(n321), .I2(n330), .O(n345) );
  NAND_GATE U374 ( .I1(B[45]), .I2(A[45]), .O(n330) );
  OR_GATE U375 ( .I1(A[45]), .I2(B[45]), .O(n321) );
  AND_GATE U376 ( .I1(n348), .I2(n349), .O(SUM[44]) );
  NAND_GATE U377 ( .I1(n351), .I2(n352), .O(n326) );
  NAND_GATE U378 ( .I1(n353), .I2(n354), .O(n352) );
  NAND_GATE U379 ( .I1(n355), .I2(n356), .O(n353) );
  NAND_GATE U380 ( .I1(n357), .I2(n358), .O(n356) );
  NAND_GATE U381 ( .I1(n359), .I2(n360), .O(n358) );
  AND_GATE U382 ( .I1(n361), .I2(n362), .O(n357) );
  AND_GATE U383 ( .I1(n170), .I2(n339), .O(n350) );
  NAND_GATE U384 ( .I1(B[44]), .I2(A[44]), .O(n332) );
  OR_GATE U385 ( .I1(A[44]), .I2(B[44]), .O(n322) );
  AND_GATE U386 ( .I1(n364), .I2(n365), .O(SUM[43]) );
  NAND_GATE U387 ( .I1(n19), .I2(n366), .O(n364) );
  NAND3_GATE U388 ( .I1(n355), .I2(n367), .I3(n368), .O(n366) );
  NAND3_GATE U389 ( .I1(n174), .I2(n361), .I3(n339), .O(n368) );
  NAND_GATE U390 ( .I1(n369), .I2(n361), .O(n367) );
  NAND_GATE U391 ( .I1(B[43]), .I2(A[43]), .O(n351) );
  OR_GATE U392 ( .I1(A[43]), .I2(B[43]), .O(n354) );
  AND_GATE U393 ( .I1(n370), .I2(n371), .O(SUM[42]) );
  NAND_GATE U394 ( .I1(n373), .I2(n359), .O(n369) );
  AND_GATE U395 ( .I1(n174), .I2(n339), .O(n372) );
  NAND_GATE U396 ( .I1(B[42]), .I2(A[42]), .O(n355) );
  OR_GATE U397 ( .I1(A[42]), .I2(B[42]), .O(n361) );
  AND_GATE U398 ( .I1(n374), .I2(n375), .O(SUM[41]) );
  NAND_GATE U399 ( .I1(n339), .I2(n363), .O(n378) );
  INV_GATE U400 ( .I1(n376), .O(n377) );
  NAND_GATE U401 ( .I1(n362), .I2(n359), .O(n376) );
  NAND_GATE U402 ( .I1(B[41]), .I2(A[41]), .O(n359) );
  OR_GATE U403 ( .I1(A[41]), .I2(B[41]), .O(n362) );
  AND_GATE U404 ( .I1(n379), .I2(n380), .O(SUM[40]) );
  NAND_GATE U405 ( .I1(n97), .I2(n381), .O(n380) );
  NAND_GATE U406 ( .I1(n382), .I2(n339), .O(n379) );
  OR3_GATE U407 ( .I1(n311), .I2(n383), .I3(n384), .O(n339) );
  AND_GATE U408 ( .I1(n195), .I2(n385), .O(n384) );
  NAND_GATE U409 ( .I1(n390), .I2(n391), .O(n311) );
  NAND3_GATE U410 ( .I1(n386), .I2(n392), .I3(n393), .O(n391) );
  NAND3_GATE U411 ( .I1(n394), .I2(n395), .I3(n396), .O(n393) );
  NAND_GATE U412 ( .I1(n397), .I2(n395), .O(n392) );
  NAND_GATE U413 ( .I1(n387), .I2(n388), .O(n397) );
  INV_GATE U414 ( .I1(n381), .O(n382) );
  NAND_GATE U415 ( .I1(n363), .I2(n360), .O(n381) );
  NAND_GATE U416 ( .I1(B[40]), .I2(A[40]), .O(n360) );
  OR_GATE U417 ( .I1(A[40]), .I2(B[40]), .O(n363) );
  AND_GATE U418 ( .I1(n398), .I2(n399), .O(SUM[39]) );
  NAND_GATE U419 ( .I1(n34), .I2(n400), .O(n398) );
  NAND3_GATE U420 ( .I1(n395), .I2(n401), .I3(n402), .O(n400) );
  NAND3_GATE U421 ( .I1(n387), .I2(n388), .I3(n403), .O(n402) );
  NAND_GATE U422 ( .I1(n404), .I2(n387), .O(n401) );
  INV_GATE U423 ( .I1(n394), .O(n404) );
  NAND_GATE U424 ( .I1(B[39]), .I2(A[39]), .O(n390) );
  OR_GATE U425 ( .I1(A[39]), .I2(B[39]), .O(n386) );
  AND_GATE U426 ( .I1(n405), .I2(n406), .O(SUM[38]) );
  NAND_GATE U427 ( .I1(n85), .I2(n408), .O(n406) );
  NAND_GATE U428 ( .I1(n403), .I2(n388), .O(n408) );
  NAND_GATE U429 ( .I1(n387), .I2(n395), .O(n407) );
  NAND_GATE U430 ( .I1(B[38]), .I2(A[38]), .O(n395) );
  OR_GATE U431 ( .I1(A[38]), .I2(B[38]), .O(n387) );
  AND_GATE U432 ( .I1(n409), .I2(n410), .O(SUM[37]) );
  NAND_GATE U433 ( .I1(n168), .I2(n411), .O(n410) );
  NAND_GATE U434 ( .I1(n412), .I2(n403), .O(n409) );
  NAND3_GATE U435 ( .I1(n396), .I2(n413), .I3(n414), .O(n403) );
  NAND_GATE U436 ( .I1(n385), .I2(n389), .O(n414) );
  NAND3_GATE U437 ( .I1(n207), .I2(n389), .I3(n208), .O(n413) );
  INV_GATE U438 ( .I1(n411), .O(n412) );
  NAND_GATE U439 ( .I1(n388), .I2(n394), .O(n411) );
  NAND_GATE U440 ( .I1(B[37]), .I2(A[37]), .O(n394) );
  OR_GATE U441 ( .I1(A[37]), .I2(B[37]), .O(n388) );
  AND_GATE U442 ( .I1(n415), .I2(n416), .O(SUM[36]) );
  NAND_GATE U443 ( .I1(n318), .I2(n418), .O(n385) );
  NAND3_GATE U444 ( .I1(n419), .I2(n420), .I3(n428), .O(n319) );
  INV_GATE U445 ( .I1(A[32]), .O(n422) );
  INV_GATE U446 ( .I1(B[32]), .O(n423) );
  NAND_GATE U447 ( .I1(n424), .I2(n420), .O(n318) );
  NAND_GATE U448 ( .I1(n425), .I2(n426), .O(n424) );
  AND_GATE U449 ( .I1(n207), .I2(n208), .O(n417) );
  NAND4_GATE U450 ( .I1(n419), .I2(n420), .I3(n428), .I4(n429), .O(n427) );
  NAND_GATE U451 ( .I1(B[36]), .I2(A[36]), .O(n396) );
  OR_GATE U452 ( .I1(A[36]), .I2(B[36]), .O(n389) );
  AND_GATE U453 ( .I1(n430), .I2(n431), .O(SUM[35]) );
  NAND_GATE U454 ( .I1(n62), .I2(n433), .O(n431) );
  NAND_GATE U455 ( .I1(n434), .I2(n419), .O(n433) );
  NAND_GATE U456 ( .I1(n425), .I2(n420), .O(n432) );
  OR_GATE U457 ( .I1(A[35]), .I2(B[35]), .O(n420) );
  NAND_GATE U458 ( .I1(B[35]), .I2(A[35]), .O(n425) );
  AND_GATE U459 ( .I1(n435), .I2(n436), .O(SUM[34]) );
  NAND_GATE U460 ( .I1(n123), .I2(n437), .O(n436) );
  NAND_GATE U461 ( .I1(n438), .I2(n434), .O(n435) );
  NAND3_GATE U462 ( .I1(n421), .I2(n439), .I3(n440), .O(n434) );
  NAND_GATE U463 ( .I1(n441), .I2(n428), .O(n439) );
  INV_GATE U464 ( .I1(n442), .O(n441) );
  INV_GATE U465 ( .I1(n437), .O(n438) );
  NAND_GATE U466 ( .I1(n419), .I2(n426), .O(n437) );
  NAND_GATE U467 ( .I1(B[34]), .I2(A[34]), .O(n426) );
  OR_GATE U468 ( .I1(A[34]), .I2(B[34]), .O(n419) );
  AND_GATE U469 ( .I1(n443), .I2(n444), .O(SUM[33]) );
  NAND_GATE U470 ( .I1(n208), .I2(n429), .O(n447) );
  INV_GATE U471 ( .I1(n445), .O(n446) );
  NAND_GATE U472 ( .I1(n428), .I2(n421), .O(n445) );
  NAND_GATE U473 ( .I1(B[33]), .I2(A[33]), .O(n421) );
  OR_GATE U474 ( .I1(A[33]), .I2(B[33]), .O(n428) );
  AND_GATE U475 ( .I1(n448), .I2(n449), .O(SUM[32]) );
  NAND_GATE U476 ( .I1(n124), .I2(n450), .O(n449) );
  NAND_GATE U477 ( .I1(n451), .I2(n208), .O(n448) );
  NAND3_GATE U478 ( .I1(A[30]), .I2(B[30]), .I3(n312), .O(n209) );
  INV_GATE U479 ( .I1(n450), .O(n451) );
  NAND_GATE U480 ( .I1(n429), .I2(n442), .O(n450) );
  NAND_GATE U481 ( .I1(B[32]), .I2(A[32]), .O(n442) );
  OR_GATE U482 ( .I1(A[32]), .I2(B[32]), .O(n429) );
  AND_GATE U483 ( .I1(n452), .I2(n453), .O(SUM[31]) );
  NAND_GATE U484 ( .I1(n37), .I2(n36), .O(n452) );
  OR_GATE U485 ( .I1(A[31]), .I2(B[31]), .O(n312) );
  NAND_GATE U486 ( .I1(B[31]), .I2(A[31]), .O(n210) );
  NAND_GATE U487 ( .I1(n313), .I2(n454), .O(n455) );
  NAND_GATE U488 ( .I1(B[30]), .I2(A[30]), .O(n454) );
endmodule


module alu_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] ,
         \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] ,
         \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] ,
         \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] ,
         \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] ,
         \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] ,
         \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[61] , \A2[60] ,
         \A2[59] , \A2[57] , \A2[55] , \A2[53] , \A2[51] , \A2[49] , \A2[47] ,
         \A2[45] , \A2[43] , \A2[41] , \A2[39] , \A2[38] , \A2[37] , \A2[36] ,
         \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15379;

  alu_DW01_add_11 FS_1 ( .A({1'b0, \A1[60] , \A1[59] , \A1[58] , \A1[57] , 
        \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , 
        \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , 
        \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , 
        \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , 
        \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , 
        \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , 
        \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[61] , \A2[60] , \A2[59] , n15376, \A2[57] , n15373, \A2[55] , 
        n15374, \A2[53] , n15372, \A2[51] , n15370, \A2[49] , n15371, \A2[47] , 
        n15375, \A2[45] , n15369, \A2[43] , n15368, \A2[41] , n15367, \A2[39] , 
        \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , 
        \A2[31] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM(PRODUCT[63:2]) );
  AND3_GATE U2 ( .I1(n4855), .I2(n4854), .I3(n4853), .O(n3) );
  AND3_GATE U3 ( .I1(n8904), .I2(n8903), .I3(n8902), .O(n4) );
  AND3_GATE U4 ( .I1(n9724), .I2(n9732), .I3(n9543), .O(n5) );
  AND_GATE U5 ( .I1(n2046), .I2(n1884), .O(n6) );
  AND_GATE U6 ( .I1(n2035), .I2(n1859), .O(n7) );
  AND_GATE U7 ( .I1(n2899), .I2(n2898), .O(n8) );
  AND3_GATE U8 ( .I1(n8839), .I2(n8838), .I3(n8683), .O(n9) );
  NAND_GATE U9 ( .I1(n9772), .I2(n13), .O(n10) );
  AND_GATE U10 ( .I1(n10), .I2(n11), .O(n9756) );
  OR_GATE U11 ( .I1(n12), .I2(n9517), .O(n11) );
  INV_GATE U12 ( .I1(n9758), .O(n12) );
  AND_GATE U13 ( .I1(n9774), .I2(n9758), .O(n13) );
  NOR_GATE U14 ( .I1(n1212), .I2(n1045), .O(n14) );
  AND_GATE U15 ( .I1(n10088), .I2(n10087), .O(n15) );
  AND3_GATE U16 ( .I1(n12261), .I2(n12254), .I3(n12253), .O(n16) );
  AND3_GATE U17 ( .I1(n4434), .I2(n4433), .I3(n4432), .O(n17) );
  AND3_GATE U18 ( .I1(n7986), .I2(n7985), .I3(n7729), .O(n18) );
  AND_GATE U19 ( .I1(n9517), .I2(n9516), .O(n19) );
  AND_GATE U20 ( .I1(n6451), .I2(n6450), .O(n20) );
  INV_GATE U21 ( .I1(n20), .O(n6544) );
  AND3_GATE U22 ( .I1(n14873), .I2(n14872), .I3(n14871), .O(n21) );
  AND_GATE U23 ( .I1(n15042), .I2(n15024), .O(n22) );
  OR_GATE U24 ( .I1(n633), .I2(n26), .O(n23) );
  AND_GATE U25 ( .I1(n23), .I2(n24), .O(n9979) );
  OR_GATE U26 ( .I1(n25), .I2(n9976), .O(n24) );
  INV_GATE U27 ( .I1(n9978), .O(n25) );
  OR_GATE U28 ( .I1(n9975), .I2(n25), .O(n26) );
  AND_GATE U29 ( .I1(n10220), .I2(n10218), .O(n27) );
  NAND_GATE U30 ( .I1(n552), .I2(n27), .O(n29) );
  NAND_GATE U31 ( .I1(n10216), .I2(n30), .O(n28) );
  AND_GATE U32 ( .I1(n28), .I2(n29), .O(n10221) );
  AND_GATE U33 ( .I1(n10215), .I2(n10220), .O(n30) );
  NAND_GATE U34 ( .I1(n10221), .I2(n34), .O(n31) );
  AND_GATE U35 ( .I1(n31), .I2(n32), .O(n10695) );
  OR_GATE U36 ( .I1(n33), .I2(n10224), .O(n32) );
  INV_GATE U37 ( .I1(n10349), .O(n33) );
  AND_GATE U38 ( .I1(n10222), .I2(n10349), .O(n34) );
  NAND_GATE U39 ( .I1(n11105), .I2(n38), .O(n35) );
  AND_GATE U40 ( .I1(n35), .I2(n36), .O(n11108) );
  OR_GATE U41 ( .I1(n37), .I2(n11106), .O(n36) );
  INV_GATE U42 ( .I1(n11107), .O(n37) );
  AND_GATE U43 ( .I1(n11104), .I2(n11107), .O(n38) );
  AND_GATE U44 ( .I1(n11291), .I2(n11288), .O(n39) );
  NAND_GATE U45 ( .I1(n11289), .I2(n39), .O(n70) );
  AND_GATE U46 ( .I1(n11734), .I2(n11733), .O(n40) );
  NAND_GATE U47 ( .I1(n11978), .I2(n41), .O(n43) );
  AND_GATE U48 ( .I1(n11976), .I2(n40), .O(n41) );
  NAND_GATE U49 ( .I1(n11974), .I2(n44), .O(n42) );
  AND_GATE U50 ( .I1(n42), .I2(n43), .O(n11979) );
  AND_GATE U51 ( .I1(n11973), .I2(n11978), .O(n44) );
  NAND_GATE U52 ( .I1(n13517), .I2(n48), .O(n45) );
  AND_GATE U53 ( .I1(n45), .I2(n46), .O(n13924) );
  OR_GATE U54 ( .I1(n47), .I2(n13669), .O(n46) );
  INV_GATE U55 ( .I1(n13519), .O(n47) );
  AND_GATE U56 ( .I1(n13672), .I2(n13519), .O(n48) );
  AND_GATE U57 ( .I1(n13518), .I2(n13669), .O(n49) );
  AND_GATE U58 ( .I1(n13516), .I2(n13515), .O(n50) );
  NAND_GATE U59 ( .I1(n13670), .I2(n13675), .O(n62) );
  NAND_GATE U60 ( .I1(n12837), .I2(n54), .O(n51) );
  AND_GATE U61 ( .I1(n51), .I2(n52), .O(n13510) );
  OR_GATE U62 ( .I1(n53), .I2(n12840), .O(n52) );
  INV_GATE U63 ( .I1(n12842), .O(n53) );
  AND_GATE U64 ( .I1(n12838), .I2(n12842), .O(n54) );
  AND_GATE U65 ( .I1(n13284), .I2(n13286), .O(n55) );
  NAND_GATE U66 ( .I1(n13283), .I2(n55), .O(n57) );
  NAND_GATE U67 ( .I1(n13281), .I2(n58), .O(n56) );
  AND_GATE U68 ( .I1(n56), .I2(n57), .O(n13287) );
  AND_GATE U69 ( .I1(n13280), .I2(n13286), .O(n58) );
  OR_GATE U70 ( .I1(n13672), .I2(n62), .O(n59) );
  AND_GATE U71 ( .I1(n59), .I2(n60), .O(n13676) );
  OR_GATE U72 ( .I1(n61), .I2(n13673), .O(n60) );
  INV_GATE U73 ( .I1(n13675), .O(n61) );
  AND3_GATE U74 ( .I1(n13922), .I2(n14361), .I3(n14360), .O(n63) );
  NAND_GATE U75 ( .I1(n11799), .I2(n64), .O(n66) );
  NOR_GATE U76 ( .I1(n11804), .I2(n67), .O(n64) );
  NAND_GATE U77 ( .I1(n11797), .I2(n68), .O(n65) );
  AND_GATE U78 ( .I1(n65), .I2(n66), .O(n11801) );
  INV_GATE U79 ( .I1(n11800), .O(n67) );
  AND_GATE U80 ( .I1(n11804), .I2(n11800), .O(n68) );
  NAND_GATE U81 ( .I1(n11286), .I2(n71), .O(n69) );
  AND_GATE U82 ( .I1(n69), .I2(n70), .O(n11292) );
  AND_GATE U83 ( .I1(n11287), .I2(n11291), .O(n71) );
  OR_GATE U84 ( .I1(n6857), .I2(n87), .O(n6853) );
  OR_GATE U85 ( .I1(n6873), .I2(n83), .O(n6869) );
  NAND_GATE U86 ( .I1(n8706), .I2(n75), .O(n72) );
  AND_GATE U87 ( .I1(n72), .I2(n73), .O(n8710) );
  OR_GATE U88 ( .I1(n74), .I2(n8708), .O(n73) );
  INV_GATE U89 ( .I1(n8709), .O(n74) );
  AND_GATE U90 ( .I1(n8707), .I2(n8709), .O(n75) );
  NAND_GATE U91 ( .I1(n8710), .I2(n79), .O(n76) );
  AND_GATE U92 ( .I1(n76), .I2(n77), .O(n8816) );
  OR_GATE U93 ( .I1(n78), .I2(n8713), .O(n77) );
  INV_GATE U94 ( .I1(n8714), .O(n78) );
  AND_GATE U95 ( .I1(n8711), .I2(n8714), .O(n79) );
  AND3_GATE U96 ( .I1(n8817), .I2(n8816), .I3(n8715), .O(n80) );
  OR_GATE U97 ( .I1(n6861), .I2(n6872), .O(n6866) );
  NAND_GATE U98 ( .I1(n6871), .I2(n84), .O(n81) );
  AND_GATE U99 ( .I1(n81), .I2(n82), .O(n7070) );
  OR_GATE U100 ( .I1(n83), .I2(n6873), .O(n82) );
  INV_GATE U101 ( .I1(n6874), .O(n83) );
  AND_GATE U102 ( .I1(n6872), .I2(n6874), .O(n84) );
  OR_GATE U103 ( .I1(n6856), .I2(n6848), .O(n6850) );
  NAND_GATE U104 ( .I1(n6855), .I2(n88), .O(n85) );
  AND_GATE U105 ( .I1(n85), .I2(n86), .O(n7081) );
  OR_GATE U106 ( .I1(n87), .I2(n6857), .O(n86) );
  INV_GATE U107 ( .I1(n6858), .O(n87) );
  AND_GATE U108 ( .I1(n6856), .I2(n6858), .O(n88) );
  AND3_GATE U109 ( .I1(n7078), .I2(n7077), .I3(n6859), .O(n89) );
  AND_GATE U110 ( .I1(n7757), .I2(n7457), .O(n90) );
  NAND_GATE U111 ( .I1(n7782), .I2(n94), .O(n91) );
  AND_GATE U112 ( .I1(n91), .I2(n92), .O(n7939) );
  OR_GATE U113 ( .I1(n93), .I2(n7785), .O(n92) );
  INV_GATE U114 ( .I1(n7786), .O(n93) );
  AND_GATE U115 ( .I1(n7783), .I2(n7786), .O(n94) );
  AND3_GATE U116 ( .I1(n8806), .I2(n8805), .I3(n8731), .O(n95) );
  NAND_GATE U117 ( .I1(n15335), .I2(n99), .O(n96) );
  AND_GATE U118 ( .I1(n96), .I2(n97), .O(n15339) );
  OR_GATE U119 ( .I1(n98), .I2(n15337), .O(n97) );
  INV_GATE U120 ( .I1(n15338), .O(n98) );
  AND_GATE U121 ( .I1(n15336), .I2(n15338), .O(n99) );
  OR_GATE U122 ( .I1(n11574), .I2(n11572), .O(n11583) );
  AND3_GATE U123 ( .I1(n10205), .I2(n10206), .I3(n10212), .O(n100) );
  AND3_GATE U124 ( .I1(n11093), .I2(n11094), .I3(n11100), .O(n101) );
  NAND_GATE U125 ( .I1(n11567), .I2(n102), .O(n119) );
  AND_GATE U126 ( .I1(n101), .I2(n11565), .O(n102) );
  OR_GATE U127 ( .I1(n11573), .I2(n103), .O(n864) );
  NAND_GATE U128 ( .I1(n11577), .I2(n11579), .O(n103) );
  NAND_GATE U129 ( .I1(n11272), .I2(n107), .O(n104) );
  AND_GATE U130 ( .I1(n104), .I2(n105), .O(n11275) );
  OR_GATE U131 ( .I1(n106), .I2(n11273), .O(n105) );
  INV_GATE U132 ( .I1(n11274), .O(n106) );
  AND_GATE U133 ( .I1(n11271), .I2(n11274), .O(n107) );
  NAND_GATE U134 ( .I1(n11950), .I2(n108), .O(n122) );
  AND_GATE U135 ( .I1(n11955), .I2(n686), .O(n108) );
  OR_GATE U136 ( .I1(n11541), .I2(n11547), .O(n11539) );
  NAND_GATE U137 ( .I1(n11546), .I2(n112), .O(n109) );
  AND_GATE U138 ( .I1(n109), .I2(n110), .O(n11938) );
  OR_GATE U139 ( .I1(n111), .I2(n11548), .O(n110) );
  INV_GATE U140 ( .I1(n11549), .O(n111) );
  AND_GATE U141 ( .I1(n11547), .I2(n11549), .O(n112) );
  AND_GATE U142 ( .I1(n11948), .I2(n11756), .O(n113) );
  NOR_GATE U143 ( .I1(n12398), .I2(n12399), .O(n115) );
  NAND_GATE U144 ( .I1(n12180), .I2(n12181), .O(n114) );
  NAND_GATE U145 ( .I1(n114), .I2(n115), .O(n12396) );
  AND_GATE U146 ( .I1(n12807), .I2(n12660), .O(n116) );
  NAND_GATE U147 ( .I1(n11573), .I2(n117), .O(n865) );
  NOR_GATE U148 ( .I1(n11577), .I2(n11575), .O(n117) );
  NAND_GATE U149 ( .I1(n11562), .I2(n120), .O(n118) );
  AND_GATE U150 ( .I1(n118), .I2(n119), .O(n11568) );
  AND_GATE U151 ( .I1(n11563), .I2(n11567), .O(n120) );
  NAND_GATE U152 ( .I1(n11955), .I2(n121), .O(n123) );
  NOR_GATE U153 ( .I1(n11950), .I2(n686), .O(n121) );
  AND_GATE U154 ( .I1(n122), .I2(n123), .O(n11956) );
  AND3_GATE U155 ( .I1(n12658), .I2(n13073), .I3(n13072), .O(n124) );
  OR_GATE U156 ( .I1(n13248), .I2(n125), .O(n373) );
  NAND_GATE U157 ( .I1(n13249), .I2(n13250), .O(n125) );
  NAND_GATE U158 ( .I1(n11963), .I2(n129), .O(n126) );
  AND_GATE U159 ( .I1(n126), .I2(n127), .O(n11967) );
  OR_GATE U160 ( .I1(n128), .I2(n11965), .O(n127) );
  INV_GATE U161 ( .I1(n11966), .O(n128) );
  AND_GATE U162 ( .I1(n11964), .I2(n11966), .O(n129) );
  OR_GATE U163 ( .I1(n10450), .I2(n10455), .O(n10460) );
  AND_GATE U164 ( .I1(n8652), .I2(n8651), .O(n130) );
  NAND_GATE U165 ( .I1(n11568), .I2(n134), .O(n131) );
  AND_GATE U166 ( .I1(n131), .I2(n132), .O(n12152) );
  OR_GATE U167 ( .I1(n133), .I2(n11571), .O(n132) );
  INV_GATE U168 ( .I1(n11753), .O(n133) );
  AND_GATE U169 ( .I1(n11569), .I2(n11753), .O(n134) );
  NAND_GATE U170 ( .I1(n12419), .I2(n135), .O(n688) );
  AND_GATE U171 ( .I1(n12418), .I2(n136), .O(n135) );
  INV_GATE U172 ( .I1(n12420), .O(n136) );
  OR_GATE U173 ( .I1(n137), .I2(n10416), .O(n10414) );
  INV_GATE U174 ( .I1(n10413), .O(n137) );
  NAND_GATE U175 ( .I1(n12692), .I2(n141), .O(n138) );
  AND_GATE U176 ( .I1(n138), .I2(n139), .O(n12779) );
  OR_GATE U177 ( .I1(n140), .I2(n13123), .O(n139) );
  INV_GATE U178 ( .I1(n12778), .O(n140) );
  AND_GATE U179 ( .I1(n13124), .I2(n12778), .O(n141) );
  AND_GATE U180 ( .I1(n12210), .I2(n12211), .O(n142) );
  NAND_GATE U181 ( .I1(n12209), .I2(n142), .O(n144) );
  NAND_GATE U182 ( .I1(n12207), .I2(n145), .O(n143) );
  AND_GATE U183 ( .I1(n143), .I2(n144), .O(n12212) );
  AND_GATE U184 ( .I1(n12208), .I2(n12211), .O(n145) );
  NAND_GATE U185 ( .I1(n11398), .I2(n149), .O(n146) );
  AND_GATE U186 ( .I1(n146), .I2(n147), .O(n11365) );
  OR_GATE U187 ( .I1(n148), .I2(n11393), .O(n147) );
  INV_GATE U188 ( .I1(n11401), .O(n148) );
  AND_GATE U189 ( .I1(n11385), .I2(n11401), .O(n149) );
  NAND_GATE U190 ( .I1(n11398), .I2(n153), .O(n150) );
  AND_GATE U191 ( .I1(n150), .I2(n151), .O(n11366) );
  OR_GATE U192 ( .I1(n152), .I2(n11393), .O(n151) );
  INV_GATE U193 ( .I1(n11386), .O(n152) );
  AND_GATE U194 ( .I1(n11385), .I2(n11386), .O(n153) );
  AND_GATE U195 ( .I1(n11342), .I2(n10920), .O(n154) );
  INV_GATE U196 ( .I1(n154), .O(n11001) );
  AND_GATE U197 ( .I1(n5870), .I2(n5871), .O(n155) );
  AND_GATE U198 ( .I1(n6087), .I2(n6086), .O(n156) );
  AND_GATE U199 ( .I1(n12741), .I2(n12712), .O(n157) );
  INV_GATE U200 ( .I1(n157), .O(n12726) );
  NAND3_GATE U201 ( .I1(n8114), .I2(n8113), .I3(n8112), .O(n158) );
  INV_GATE U202 ( .I1(n158), .O(n874) );
  OR_GATE U203 ( .I1(n746), .I2(n159), .O(n8560) );
  INV_GATE U204 ( .I1(n8979), .O(n159) );
  NAND_GATE U205 ( .I1(n8564), .I2(n163), .O(n160) );
  AND_GATE U206 ( .I1(n160), .I2(n161), .O(n8568) );
  OR_GATE U207 ( .I1(n162), .I2(n8562), .O(n161) );
  INV_GATE U208 ( .I1(n8567), .O(n162) );
  AND_GATE U209 ( .I1(n8571), .I2(n8567), .O(n163) );
  OR_GATE U210 ( .I1(n10661), .I2(n170), .O(n10665) );
  AND_GATE U211 ( .I1(n10033), .I2(n10166), .O(n164) );
  INV_GATE U212 ( .I1(n164), .O(n10168) );
  AND3_GATE U213 ( .I1(n8092), .I2(n7628), .I3(n8091), .O(n165) );
  AND_GATE U214 ( .I1(n8223), .I2(n8222), .O(n166) );
  AND_GATE U215 ( .I1(n12785), .I2(n12363), .O(n167) );
  AND3_GATE U216 ( .I1(n8962), .I2(n8576), .I3(n8961), .O(n168) );
  AND_GATE U217 ( .I1(n5670), .I2(n5669), .O(n169) );
  OR_GATE U218 ( .I1(n9834), .I2(n632), .O(n9467) );
  OR_GATE U219 ( .I1(n4505), .I2(n820), .O(n4725) );
  AND_GATE U220 ( .I1(n10671), .I2(n10368), .O(n170) );
  INV_GATE U221 ( .I1(n170), .O(n10667) );
  OR3_GATE U222 ( .I1(n171), .I2(n9836), .I3(n172), .O(n9839) );
  INV_GATE U223 ( .I1(n9473), .O(n171) );
  INV_GATE U224 ( .I1(n9837), .O(n172) );
  AND_GATE U225 ( .I1(n7618), .I2(n7617), .O(n173) );
  AND_GATE U226 ( .I1(n4749), .I2(n4748), .O(n174) );
  AND_GATE U227 ( .I1(n8318), .I2(n8317), .O(n175) );
  INV_GATE U228 ( .I1(n175), .O(n8644) );
  AND_GATE U229 ( .I1(n9528), .I2(n9206), .O(n176) );
  INV_GATE U230 ( .I1(n176), .O(n9536) );
  OR_GATE U231 ( .I1(n177), .I2(n5809), .O(n5807) );
  AND3_GATE U232 ( .I1(n5550), .I2(n5549), .I3(n5370), .O(n177) );
  NAND_GATE U233 ( .I1(n178), .I2(n8876), .O(n8878) );
  NOR_GATE U234 ( .I1(n8887), .I2(n8886), .O(n178) );
  NAND_GATE U235 ( .I1(n4841), .I2(n182), .O(n179) );
  AND_GATE U236 ( .I1(n179), .I2(n180), .O(n5371) );
  OR_GATE U237 ( .I1(n181), .I2(n4843), .O(n180) );
  INV_GATE U238 ( .I1(n5375), .O(n181) );
  AND_GATE U239 ( .I1(n258), .I2(n5375), .O(n182) );
  AND_GATE U240 ( .I1(n9714), .I2(n9715), .O(n183) );
  AND_GATE U241 ( .I1(n9716), .I2(n183), .O(n10443) );
  AND3_GATE U242 ( .I1(n7398), .I2(n6747), .I3(n6746), .O(n184) );
  INV_GATE U243 ( .I1(n184), .O(n7174) );
  NOR_GATE U244 ( .I1(n2003), .I2(n1307), .O(n185) );
  INV_GATE U245 ( .I1(n185), .O(n2797) );
  AND_GATE U246 ( .I1(n8602), .I2(n8599), .O(n186) );
  INV_GATE U247 ( .I1(n186), .O(n9180) );
  AND3_GATE U248 ( .I1(n11879), .I2(n11813), .I3(n11880), .O(n187) );
  INV_GATE U249 ( .I1(n187), .O(n11875) );
  AND_GATE U250 ( .I1(n11803), .I2(n11314), .O(n188) );
  INV_GATE U251 ( .I1(n188), .O(n11495) );
  AND3_GATE U252 ( .I1(n7344), .I2(n7534), .I3(n7535), .O(n189) );
  INV_GATE U253 ( .I1(n189), .O(n7624) );
  NOR_GATE U254 ( .I1(n11894), .I2(n11895), .O(n190) );
  INV_GATE U255 ( .I1(n190), .O(n11899) );
  NAND_GATE U256 ( .I1(n6678), .I2(n194), .O(n191) );
  AND_GATE U257 ( .I1(n191), .I2(n192), .O(n6683) );
  OR_GATE U258 ( .I1(n193), .I2(n6682), .O(n192) );
  INV_GATE U259 ( .I1(n7248), .O(n193) );
  AND_GATE U260 ( .I1(n6679), .I2(n7248), .O(n194) );
  NAND_GATE U261 ( .I1(n11313), .I2(n198), .O(n195) );
  AND_GATE U262 ( .I1(n195), .I2(n196), .O(n11490) );
  OR_GATE U263 ( .I1(n197), .I2(n11803), .O(n196) );
  INV_GATE U264 ( .I1(n11489), .O(n197) );
  AND_GATE U265 ( .I1(n11804), .I2(n11489), .O(n198) );
  AND_GATE U266 ( .I1(n4738), .I2(n4739), .O(n199) );
  OR3_GATE U267 ( .I1(n201), .I2(n200), .I3(n3874), .O(n3878) );
  INV_GATE U268 ( .I1(n3875), .O(n200) );
  AND_GATE U269 ( .I1(n3873), .I2(n3872), .O(n201) );
  NAND_GATE U270 ( .I1(n808), .I2(n809), .O(n202) );
  INV_GATE U271 ( .I1(n202), .O(n8284) );
  NAND_GATE U272 ( .I1(n813), .I2(n206), .O(n203) );
  AND_GATE U273 ( .I1(n203), .I2(n204), .O(n5523) );
  OR_GATE U274 ( .I1(n205), .I2(n4821), .O(n204) );
  INV_GATE U275 ( .I1(n5513), .O(n205) );
  AND_GATE U276 ( .I1(n4823), .I2(n5513), .O(n206) );
  AND_GATE U277 ( .I1(n7371), .I2(n7370), .O(n207) );
  AND3_GATE U278 ( .I1(n6448), .I2(n6447), .I3(n6446), .O(n208) );
  AND_GATE U279 ( .I1(n7425), .I2(n827), .O(n209) );
  AND3_GATE U280 ( .I1(n9202), .I2(n9201), .I3(n9200), .O(n210) );
  NAND_GATE U281 ( .I1(n4842), .I2(n214), .O(n211) );
  AND_GATE U282 ( .I1(n211), .I2(n212), .O(n4846) );
  OR_GATE U283 ( .I1(n213), .I2(n4844), .O(n212) );
  INV_GATE U284 ( .I1(n5375), .O(n213) );
  AND_GATE U285 ( .I1(n706), .I2(n5375), .O(n214) );
  AND_GATE U286 ( .I1(n2792), .I2(n2791), .O(n215) );
  AND_GATE U287 ( .I1(n4591), .I2(n4588), .O(n216) );
  AND4_GATE U288 ( .I1(n1875), .I2(n1874), .I3(n1873), .I4(n1872), .O(n217) );
  AND3_GATE U289 ( .I1(n9737), .I2(n9534), .I3(n9533), .O(n218) );
  NAND_GATE U290 ( .I1(n5812), .I2(n6288), .O(n219) );
  INV_GATE U291 ( .I1(n219), .O(n259) );
  OR_GATE U292 ( .I1(n6390), .I2(n6398), .O(n5764) );
  OR_GATE U293 ( .I1(n220), .I2(n794), .O(n5760) );
  INV_GATE U294 ( .I1(n6390), .O(n220) );
  AND3_GATE U295 ( .I1(n7032), .I2(n7031), .I3(n6926), .O(n221) );
  AND_GATE U296 ( .I1(n3048), .I2(n2821), .O(n222) );
  AND_GATE U297 ( .I1(n3073), .I2(n3072), .O(n223) );
  AND3_GATE U298 ( .I1(n2698), .I2(n2697), .I3(n2696), .O(n224) );
  AND_GATE U299 ( .I1(n2034), .I2(n2029), .O(n225) );
  INV_GATE U300 ( .I1(n225), .O(n2024) );
  OR4_GATE U301 ( .I1(n226), .I2(n227), .I3(n805), .I4(n228), .O(n3537) );
  NOR_GATE U302 ( .I1(n3059), .I2(n3546), .O(n226) );
  AND_GATE U303 ( .I1(n3548), .I2(n3058), .O(n227) );
  AND_GATE U304 ( .I1(n3543), .I2(n818), .O(n228) );
  AND_GATE U305 ( .I1(n7611), .I2(n917), .O(n229) );
  AND3_GATE U306 ( .I1(n467), .I2(n523), .I3(n477), .O(n230) );
  AND_GATE U307 ( .I1(n12379), .I2(n12378), .O(n231) );
  AND_GATE U308 ( .I1(n12186), .I2(n11777), .O(n232) );
  AND_GATE U309 ( .I1(n11076), .I2(n11075), .O(n233) );
  AND_GATE U310 ( .I1(n11761), .I2(n11299), .O(n234) );
  OR_GATE U311 ( .I1(n6423), .I2(n784), .O(n6421) );
  AND_GATE U312 ( .I1(n3018), .I2(n3015), .O(n235) );
  INV_GATE U313 ( .I1(n235), .O(n3579) );
  NAND_GATE U314 ( .I1(n10169), .I2(n239), .O(n236) );
  AND_GATE U315 ( .I1(n236), .I2(n237), .O(n10371) );
  OR_GATE U316 ( .I1(n238), .I2(n10176), .O(n237) );
  INV_GATE U317 ( .I1(n11060), .O(n238) );
  AND_GATE U318 ( .I1(n164), .I2(n11060), .O(n239) );
  AND3_GATE U319 ( .I1(n12795), .I2(n12780), .I3(n12781), .O(n240) );
  NAND_GATE U320 ( .I1(n11000), .I2(n11004), .O(n241) );
  AND_GATE U321 ( .I1(n10912), .I2(n10402), .O(n242) );
  AND3_GATE U322 ( .I1(n10609), .I2(n10608), .I3(n10607), .O(n243) );
  AND_GATE U323 ( .I1(n10138), .I2(n10137), .O(n244) );
  AND_GATE U324 ( .I1(n7680), .I2(n7679), .O(n245) );
  AND_GATE U325 ( .I1(n9482), .I2(n9168), .O(n246) );
  AND_GATE U326 ( .I1(n12694), .I2(n12779), .O(n247) );
  AND_GATE U327 ( .I1(n12693), .I2(n247), .O(n528) );
  NAND_GATE U328 ( .I1(n8925), .I2(n251), .O(n248) );
  AND_GATE U329 ( .I1(n248), .I2(n249), .O(n8930) );
  OR_GATE U330 ( .I1(n250), .I2(n8922), .O(n249) );
  INV_GATE U331 ( .I1(n8613), .O(n250) );
  AND_GATE U332 ( .I1(n8920), .I2(n8613), .O(n251) );
  NAND_GATE U333 ( .I1(n8302), .I2(n8301), .O(n252) );
  OR_GATE U334 ( .I1(n3888), .I2(n253), .O(n4484) );
  OR_GATE U335 ( .I1(n254), .I2(n3889), .O(n253) );
  INV_GATE U336 ( .I1(n4482), .O(n254) );
  AND_GATE U337 ( .I1(n6717), .I2(n6716), .O(n255) );
  OR_GATE U338 ( .I1(n876), .I2(n256), .O(n9514) );
  AND_GATE U339 ( .I1(n9764), .I2(n9763), .O(n256) );
  AND3_GATE U340 ( .I1(n8348), .I2(n8281), .I3(n8280), .O(n257) );
  INV_GATE U341 ( .I1(n257), .O(n8603) );
  OR_GATE U342 ( .I1(n4829), .I2(n277), .O(n4832) );
  OR_GATE U343 ( .I1(n277), .I2(n216), .O(n4596) );
  AND3_GATE U344 ( .I1(n4596), .I2(n4595), .I3(n4832), .O(n258) );
  INV_GATE U345 ( .I1(n258), .O(n4842) );
  AND3_GATE U346 ( .I1(n7502), .I2(n7500), .I3(n7395), .O(n260) );
  INV_GATE U347 ( .I1(n260), .O(n7495) );
  AND_GATE U348 ( .I1(n8302), .I2(n8301), .O(n261) );
  NAND_GATE U349 ( .I1(n4845), .I2(n5380), .O(n262) );
  AND_GATE U350 ( .I1(n11392), .I2(n10950), .O(n263) );
  NAND_GATE U351 ( .I1(n4837), .I2(n266), .O(n264) );
  NAND_GATE U352 ( .I1(n264), .I2(n265), .O(n1270) );
  OR_GATE U353 ( .I1(n5387), .I2(n4838), .O(n265) );
  AND_GATE U354 ( .I1(n5532), .I2(n4845), .O(n266) );
  NAND_GATE U355 ( .I1(n267), .I2(n10960), .O(n10963) );
  NOR_GATE U356 ( .I1(n10503), .I2(n10961), .O(n267) );
  NAND_GATE U357 ( .I1(n3947), .I2(n271), .O(n268) );
  AND_GATE U358 ( .I1(n268), .I2(n269), .O(n3955) );
  OR_GATE U359 ( .I1(n270), .I2(n3946), .O(n269) );
  INV_GATE U360 ( .I1(n3954), .O(n270) );
  AND_GATE U361 ( .I1(n3948), .I2(n3954), .O(n271) );
  AND_GATE U362 ( .I1(n7740), .I2(n7455), .O(n272) );
  AND3_GATE U363 ( .I1(n2719), .I2(n2718), .I3(n2717), .O(n273) );
  AND_GATE U364 ( .I1(n2060), .I2(n2059), .O(n274) );
  AND_GATE U365 ( .I1(n10484), .I2(n10483), .O(n275) );
  NAND3_GATE U366 ( .I1(n5869), .I2(n6502), .I3(n155), .O(n6215) );
  AND_GATE U367 ( .I1(n7703), .I2(n7706), .O(n276) );
  INV_GATE U368 ( .I1(n276), .O(n7704) );
  OR_GATE U369 ( .I1(n2794), .I2(n185), .O(n2798) );
  AND_GATE U370 ( .I1(n4580), .I2(n4579), .O(n277) );
  NOR_GATE U371 ( .I1(n7009), .I2(n7017), .O(n278) );
  AND3_GATE U372 ( .I1(n10165), .I2(n1328), .I3(n10164), .O(n279) );
  AND_GATE U373 ( .I1(n2685), .I2(n800), .O(n280) );
  NOR_GATE U374 ( .I1(n881), .I2(n14061), .O(n281) );
  AND_GATE U375 ( .I1(n221), .I2(n7029), .O(n282) );
  AND_GATE U376 ( .I1(n6127), .I2(n6126), .O(n283) );
  AND_GATE U377 ( .I1(n9633), .I2(n9223), .O(n284) );
  AND_GATE U378 ( .I1(n8765), .I2(n8336), .O(n285) );
  AND_GATE U379 ( .I1(n4247), .I2(n4246), .O(n286) );
  AND_GATE U380 ( .I1(n3366), .I2(n3365), .O(n287) );
  AND_GATE U381 ( .I1(n2467), .I2(n2466), .O(n288) );
  AND_GATE U382 ( .I1(n12290), .I2(n12289), .O(n289) );
  AND3_GATE U383 ( .I1(n14465), .I2(n14464), .I3(n14463), .O(n290) );
  AND_GATE U384 ( .I1(A[1]), .I2(B[0]), .O(n291) );
  AND_GATE U385 ( .I1(n14851), .I2(n14964), .O(n292) );
  NAND_GATE U386 ( .I1(n14940), .I2(n293), .O(n298) );
  AND_GATE U387 ( .I1(n1260), .I2(n14935), .O(n293) );
  AND_GATE U388 ( .I1(n378), .I2(n296), .O(n294) );
  OR_GATE U389 ( .I1(n294), .I2(n295), .O(n299) );
  AND_GATE U390 ( .I1(n14937), .I2(n14939), .O(n295) );
  AND_GATE U391 ( .I1(n379), .I2(n14937), .O(n296) );
  NAND_GATE U392 ( .I1(n14936), .I2(n299), .O(n297) );
  AND_GATE U393 ( .I1(n297), .I2(n298), .O(\A1[26] ) );
  AND_GATE U394 ( .I1(n14972), .I2(n307), .O(n300) );
  NAND_GATE U395 ( .I1(n308), .I2(n303), .O(n301) );
  AND_GATE U396 ( .I1(n301), .I2(n302), .O(n869) );
  OR_GATE U397 ( .I1(n14972), .I2(n307), .O(n302) );
  AND_GATE U398 ( .I1(n14830), .I2(n14968), .O(n303) );
  OR_GATE U399 ( .I1(n14985), .I2(n14998), .O(n304) );
  OR_GATE U400 ( .I1(n828), .I2(n14998), .O(n15001) );
  NAND_GATE U401 ( .I1(n14890), .I2(n14889), .O(n305) );
  NAND_GATE U402 ( .I1(n14830), .I2(n308), .O(n306) );
  AND_GATE U403 ( .I1(n306), .I2(n307), .O(n14989) );
  OR_GATE U404 ( .I1(n828), .I2(n304), .O(n307) );
  AND_GATE U405 ( .I1(n15003), .I2(n14979), .O(n308) );
  NAND_GATE U406 ( .I1(n14831), .I2(n309), .O(n14832) );
  AND_GATE U407 ( .I1(n15001), .I2(n14985), .O(n309) );
  NAND_GATE U408 ( .I1(n14913), .I2(n313), .O(n310) );
  AND_GATE U409 ( .I1(n310), .I2(n311), .O(\A1[28] ) );
  OR_GATE U410 ( .I1(n312), .I2(n14915), .O(n311) );
  INV_GATE U411 ( .I1(n14917), .O(n312) );
  AND_GATE U412 ( .I1(n14914), .I2(n14917), .O(n313) );
  NAND_GATE U413 ( .I1(n907), .I2(n11961), .O(n11965) );
  AND5_GATE U414 ( .I1(n14376), .I2(n555), .I3(n554), .I4(n536), .I5(n535), 
        .O(n314) );
  OR_GATE U415 ( .I1(n14081), .I2(n315), .O(n14082) );
  INV_GATE U416 ( .I1(n14080), .O(n315) );
  NAND_GATE U417 ( .I1(n14081), .I2(n316), .O(n682) );
  NOR_GATE U418 ( .I1(n14080), .I2(n684), .O(n316) );
  NAND_GATE U419 ( .I1(n13091), .I2(n319), .O(n317) );
  NAND_GATE U420 ( .I1(n317), .I2(n318), .O(n1336) );
  OR_GATE U421 ( .I1(n13240), .I2(n13089), .O(n318) );
  AND_GATE U422 ( .I1(n13090), .I2(n13100), .O(n319) );
  NAND_GATE U423 ( .I1(n1325), .I2(n320), .O(n322) );
  AND_GATE U424 ( .I1(n13092), .I2(n13096), .O(n320) );
  NAND_GATE U425 ( .I1(n13091), .I2(n323), .O(n321) );
  AND_GATE U426 ( .I1(n321), .I2(n322), .O(n13097) );
  AND_GATE U427 ( .I1(n13090), .I2(n13096), .O(n323) );
  NAND_GATE U428 ( .I1(n12670), .I2(n326), .O(n324) );
  AND_GATE U429 ( .I1(n324), .I2(n325), .O(n12796) );
  OR_GATE U430 ( .I1(n12802), .I2(n12673), .O(n325) );
  AND_GATE U431 ( .I1(n12671), .I2(n12674), .O(n326) );
  NAND_GATE U432 ( .I1(n374), .I2(n327), .O(n13252) );
  AND_GATE U433 ( .I1(n13251), .I2(n373), .O(n327) );
  AND_GATE U434 ( .I1(n12392), .I2(n13089), .O(n328) );
  NAND_GATE U435 ( .I1(n13095), .I2(n332), .O(n329) );
  AND_GATE U436 ( .I1(n329), .I2(n330), .O(n13238) );
  OR_GATE U437 ( .I1(n331), .I2(n13098), .O(n330) );
  INV_GATE U438 ( .I1(n13099), .O(n331) );
  AND_GATE U439 ( .I1(n13096), .I2(n13099), .O(n332) );
  NAND_GATE U440 ( .I1(n12676), .I2(n335), .O(n333) );
  AND_GATE U441 ( .I1(n333), .I2(n334), .O(n13102) );
  OR_GATE U442 ( .I1(n13109), .I2(n13088), .O(n334) );
  AND_GATE U443 ( .I1(n13092), .I2(n13103), .O(n335) );
  AND_GATE U444 ( .I1(n13088), .I2(n12689), .O(n336) );
  OR_GATE U445 ( .I1(n13123), .I2(n337), .O(n13125) );
  INV_GATE U446 ( .I1(n13124), .O(n337) );
  NAND_GATE U447 ( .I1(n12680), .I2(n338), .O(n346) );
  NOR_GATE U448 ( .I1(n12685), .I2(n339), .O(n338) );
  INV_GATE U449 ( .I1(n12681), .O(n339) );
  NAND_GATE U450 ( .I1(n14849), .I2(n342), .O(n340) );
  NAND_GATE U451 ( .I1(n340), .I2(n341), .O(n383) );
  OR_GATE U452 ( .I1(n1260), .I2(n1298), .O(n341) );
  AND_GATE U453 ( .I1(n14975), .I2(n14937), .O(n342) );
  NAND_GATE U454 ( .I1(n14848), .I2(n14976), .O(n343) );
  NAND_GATE U455 ( .I1(n343), .I2(n344), .O(n14850) );
  AND_GATE U456 ( .I1(n14960), .I2(n14975), .O(n344) );
  NAND_GATE U457 ( .I1(n12678), .I2(n347), .O(n345) );
  AND_GATE U458 ( .I1(n345), .I2(n346), .O(n12682) );
  AND_GATE U459 ( .I1(n12685), .I2(n12681), .O(n347) );
  AND_GATE U460 ( .I1(n14890), .I2(n14889), .O(n348) );
  NAND_GATE U461 ( .I1(n12812), .I2(n351), .O(n349) );
  AND_GATE U462 ( .I1(n349), .I2(n350), .O(n12815) );
  OR_GATE U463 ( .I1(n12809), .I2(n12813), .O(n350) );
  AND_GATE U464 ( .I1(n12811), .I2(n12814), .O(n351) );
  NAND_GATE U465 ( .I1(n14929), .I2(n354), .O(n352) );
  AND_GATE U466 ( .I1(n352), .I2(n353), .O(n14916) );
  OR_GATE U467 ( .I1(n14914), .I2(n14927), .O(n353) );
  AND_GATE U468 ( .I1(n14875), .I2(n1342), .O(n354) );
  AND_GATE U469 ( .I1(n12411), .I2(n12410), .O(n355) );
  NAND_GATE U470 ( .I1(n629), .I2(n355), .O(n363) );
  OR_GATE U471 ( .I1(n12821), .I2(n12819), .O(n12829) );
  NAND_GATE U472 ( .I1(n12826), .I2(n359), .O(n356) );
  AND_GATE U473 ( .I1(n356), .I2(n357), .O(n13525) );
  OR_GATE U474 ( .I1(n358), .I2(n12828), .O(n357) );
  INV_GATE U475 ( .I1(n12829), .O(n358) );
  AND_GATE U476 ( .I1(n12827), .I2(n12829), .O(n359) );
  AND_GATE U477 ( .I1(n12656), .I2(n12819), .O(n360) );
  AND_GATE U478 ( .I1(n13532), .I2(n13654), .O(n361) );
  NAND_GATE U479 ( .I1(n12408), .I2(n364), .O(n362) );
  AND_GATE U480 ( .I1(n362), .I2(n363), .O(n12412) );
  AND_GATE U481 ( .I1(n12409), .I2(n12411), .O(n364) );
  AND_GATE U482 ( .I1(n13546), .I2(n13641), .O(n365) );
  OR_GATE U483 ( .I1(n13240), .I2(n13250), .O(n366) );
  NOR_GATE U484 ( .I1(n13248), .I2(n13250), .O(n367) );
  INV_GATE U485 ( .I1(n367), .O(n13245) );
  NAND_GATE U486 ( .I1(n314), .I2(n368), .O(n683) );
  AND_GATE U487 ( .I1(n14080), .I2(n14083), .O(n368) );
  NAND_GATE U488 ( .I1(n13086), .I2(n371), .O(n369) );
  AND_GATE U489 ( .I1(n369), .I2(n370), .O(n13235) );
  OR_GATE U490 ( .I1(n13248), .I2(n366), .O(n370) );
  AND_GATE U491 ( .I1(n13249), .I2(n13100), .O(n371) );
  AND_GATE U492 ( .I1(n13245), .I2(n13087), .O(n372) );
  OR_GATE U493 ( .I1(n13247), .I2(n13246), .O(n374) );
  NAND_GATE U494 ( .I1(n13630), .I2(n375), .O(n13970) );
  INV_GATE U495 ( .I1(n13629), .O(n375) );
  NAND_GATE U496 ( .I1(n13630), .I2(n376), .O(n464) );
  NOR_GATE U497 ( .I1(n13629), .I2(n466), .O(n376) );
  NAND_GATE U498 ( .I1(n14943), .I2(n377), .O(n379) );
  NOR_GATE U499 ( .I1(n14946), .I2(n14937), .O(n377) );
  OR_GATE U500 ( .I1(n1264), .I2(n13628), .O(n13968) );
  NAND_GATE U501 ( .I1(n14862), .I2(n380), .O(n378) );
  AND_GATE U502 ( .I1(n378), .I2(n379), .O(n14938) );
  AND_GATE U503 ( .I1(n14950), .I2(n1260), .O(n380) );
  NAND_GATE U504 ( .I1(n14851), .I2(n383), .O(n381) );
  NAND_GATE U505 ( .I1(n381), .I2(n382), .O(n646) );
  OR_GATE U506 ( .I1(n1260), .I2(n14942), .O(n382) );
  OR_GATE U507 ( .I1(n372), .I2(n13238), .O(n13241) );
  OR_GATE U508 ( .I1(n13992), .I2(n506), .O(n13994) );
  AND_GATE U509 ( .I1(n14477), .I2(n14476), .O(n384) );
  NAND_GATE U510 ( .I1(n4940), .I2(n388), .O(n385) );
  AND_GATE U511 ( .I1(n385), .I2(n386), .O(n5272) );
  OR_GATE U512 ( .I1(n387), .I2(n4943), .O(n386) );
  INV_GATE U513 ( .I1(n4944), .O(n387) );
  AND_GATE U514 ( .I1(n4941), .I2(n4944), .O(n388) );
  NAND_GATE U515 ( .I1(n4942), .I2(n391), .O(n389) );
  AND_GATE U516 ( .I1(n389), .I2(n390), .O(n5268) );
  OR_GATE U517 ( .I1(n5274), .I2(n4944), .O(n390) );
  AND_GATE U518 ( .I1(n4943), .I2(n4945), .O(n391) );
  AND3_GATE U519 ( .I1(n5269), .I2(n5268), .I3(n4946), .O(n392) );
  NAND_GATE U520 ( .I1(n4017), .I2(n395), .O(n393) );
  AND_GATE U521 ( .I1(n393), .I2(n394), .O(n4375) );
  OR_GATE U522 ( .I1(n4382), .I2(n4020), .O(n394) );
  AND_GATE U523 ( .I1(n4018), .I2(n4021), .O(n395) );
  AND_GATE U524 ( .I1(n4020), .I2(n4019), .O(n396) );
  AND3_GATE U525 ( .I1(n4398), .I2(n4397), .I3(n3991), .O(n397) );
  AND3_GATE U526 ( .I1(n4389), .I2(n4390), .I3(n4396), .O(n398) );
  AND_GATE U527 ( .I1(n3531), .I2(n3530), .O(n399) );
  OR_GATE U528 ( .I1(n6982), .I2(n15323), .O(n6983) );
  OR_GATE U529 ( .I1(n221), .I2(n7025), .O(n7022) );
  OR_GATE U530 ( .I1(n6877), .I2(n6882), .O(n6879) );
  AND3_GATE U531 ( .I1(n12698), .I2(n12697), .I3(n12759), .O(n400) );
  AND_GATE U532 ( .I1(n13974), .I2(n13555), .O(n401) );
  NAND_GATE U533 ( .I1(n13989), .I2(n404), .O(n402) );
  AND_GATE U534 ( .I1(n402), .I2(n403), .O(n14035) );
  OR_GATE U535 ( .I1(n14042), .I2(n14424), .O(n403) );
  AND_GATE U536 ( .I1(n14427), .I2(n14001), .O(n404) );
  OR_GATE U537 ( .I1(n13558), .I2(n407), .O(n405) );
  AND_GATE U538 ( .I1(n405), .I2(n406), .O(n13995) );
  OR_GATE U539 ( .I1(n13991), .I2(n506), .O(n406) );
  OR_GATE U540 ( .I1(n13200), .I2(n13991), .O(n407) );
  AND3_GATE U541 ( .I1(n12230), .I2(n12229), .I3(n12228), .O(n408) );
  OR_GATE U542 ( .I1(n12741), .I2(n12737), .O(n12743) );
  OR_GATE U543 ( .I1(n14083), .I2(n14396), .O(n409) );
  OR_GATE U544 ( .I1(n14083), .I2(n14080), .O(n14078) );
  AND_GATE U545 ( .I1(n13262), .I2(n13260), .O(n410) );
  NAND_GATE U546 ( .I1(n13261), .I2(n410), .O(n412) );
  NAND_GATE U547 ( .I1(n13259), .I2(n413), .O(n411) );
  AND_GATE U548 ( .I1(n411), .I2(n412), .O(n13263) );
  AND_GATE U549 ( .I1(n13258), .I2(n13262), .O(n413) );
  NAND_GATE U550 ( .I1(n13947), .I2(n416), .O(n414) );
  AND_GATE U551 ( .I1(n414), .I2(n415), .O(n14391) );
  OR_GATE U552 ( .I1(n14080), .I2(n409), .O(n415) );
  AND_GATE U553 ( .I1(n14081), .I2(n13949), .O(n416) );
  AND_GATE U554 ( .I1(n13948), .I2(n417), .O(n723) );
  AND_GATE U555 ( .I1(n14078), .I2(n13949), .O(n417) );
  AND_GATE U556 ( .I1(n13948), .I2(n14078), .O(n418) );
  AND_GATE U557 ( .I1(n13648), .I2(n13649), .O(n419) );
  NAND_GATE U558 ( .I1(n13647), .I2(n419), .O(n421) );
  NAND_GATE U559 ( .I1(n13645), .I2(n422), .O(n420) );
  AND_GATE U560 ( .I1(n420), .I2(n421), .O(n13650) );
  AND_GATE U561 ( .I1(n13646), .I2(n13649), .O(n422) );
  NAND_GATE U562 ( .I1(n14876), .I2(n426), .O(n423) );
  NAND_GATE U563 ( .I1(n423), .I2(n424), .O(n1318) );
  OR_GATE U564 ( .I1(n425), .I2(n14919), .O(n424) );
  INV_GATE U565 ( .I1(n14902), .O(n425) );
  AND_GATE U566 ( .I1(n14938), .I2(n14902), .O(n426) );
  NAND_GATE U567 ( .I1(n14876), .I2(n429), .O(n427) );
  NAND_GATE U568 ( .I1(n427), .I2(n428), .O(n598) );
  OR_GATE U569 ( .I1(n1342), .I2(n14919), .O(n428) );
  AND_GATE U570 ( .I1(n14938), .I2(n14914), .O(n429) );
  NAND_GATE U571 ( .I1(n14074), .I2(n432), .O(n430) );
  AND_GATE U572 ( .I1(n430), .I2(n431), .O(n14496) );
  OR_GATE U573 ( .I1(n14492), .I2(n14077), .O(n431) );
  AND_GATE U574 ( .I1(n14075), .I2(n14403), .O(n432) );
  NAND_GATE U575 ( .I1(n14074), .I2(n436), .O(n433) );
  AND_GATE U576 ( .I1(n433), .I2(n434), .O(n14404) );
  OR_GATE U577 ( .I1(n435), .I2(n14077), .O(n434) );
  INV_GATE U578 ( .I1(n14495), .O(n435) );
  AND_GATE U579 ( .I1(n14075), .I2(n14495), .O(n436) );
  NAND_GATE U580 ( .I1(n13637), .I2(n440), .O(n437) );
  NAND_GATE U581 ( .I1(n437), .I2(n438), .O(n1333) );
  OR_GATE U582 ( .I1(n439), .I2(n13639), .O(n438) );
  INV_GATE U583 ( .I1(n13640), .O(n439) );
  AND_GATE U584 ( .I1(n13638), .I2(n13640), .O(n440) );
  AND_GATE U585 ( .I1(n14408), .I2(n14852), .O(n441) );
  NAND_GATE U586 ( .I1(n14483), .I2(n442), .O(n520) );
  AND_GATE U587 ( .I1(n14438), .I2(n14422), .O(n442) );
  OR_GATE U588 ( .I1(n653), .I2(n443), .O(n6478) );
  AND3_GATE U589 ( .I1(n5804), .I2(n6475), .I3(n6474), .O(n443) );
  OR_GATE U590 ( .I1(n13209), .I2(n444), .O(n13211) );
  INV_GATE U591 ( .I1(n13210), .O(n444) );
  NAND_GATE U592 ( .I1(n13628), .I2(n445), .O(n465) );
  NOR_GATE U593 ( .I1(n13627), .I2(n466), .O(n445) );
  NAND_GATE U594 ( .I1(n13589), .I2(n448), .O(n446) );
  AND_GATE U595 ( .I1(n446), .I2(n447), .O(n13594) );
  OR_GATE U596 ( .I1(n13591), .I2(n514), .O(n447) );
  AND_GATE U597 ( .I1(n1201), .I2(n13593), .O(n448) );
  OR_GATE U598 ( .I1(n6751), .I2(n6752), .O(n7166) );
  OR_GATE U599 ( .I1(n6734), .I2(n6743), .O(n6732) );
  OR_GATE U600 ( .I1(n4921), .I2(n4920), .O(n4918) );
  OR_GATE U601 ( .I1(n399), .I2(n3996), .O(n3994) );
  NAND_GATE U602 ( .I1(n4001), .I2(n451), .O(n449) );
  AND_GATE U603 ( .I1(n449), .I2(n450), .O(n4387) );
  OR_GATE U604 ( .I1(n4393), .I2(n4004), .O(n450) );
  AND_GATE U605 ( .I1(n4002), .I2(n4005), .O(n451) );
  AND_GATE U606 ( .I1(n13209), .I2(n13130), .O(n452) );
  OR_GATE U607 ( .I1(n13195), .I2(n456), .O(n453) );
  AND_GATE U608 ( .I1(n453), .I2(n454), .O(n13563) );
  OR_GATE U609 ( .I1(n455), .I2(n13198), .O(n454) );
  INV_GATE U610 ( .I1(n13991), .O(n455) );
  OR_GATE U611 ( .I1(n13197), .I2(n455), .O(n456) );
  OR3_GATE U612 ( .I1(n12742), .I2(n1213), .I3(n12733), .O(n12738) );
  AND_GATE U613 ( .I1(n13578), .I2(n12743), .O(n457) );
  NAND_GATE U614 ( .I1(n12745), .I2(n12746), .O(n458) );
  NAND_GATE U615 ( .I1(n458), .I2(n459), .O(n461) );
  AND_GATE U616 ( .I1(n13163), .I2(n624), .O(n459) );
  NAND_GATE U617 ( .I1(n13159), .I2(n463), .O(n460) );
  AND_GATE U618 ( .I1(n460), .I2(n461), .O(n13165) );
  INV_GATE U619 ( .I1(n13163), .O(n462) );
  AND_GATE U620 ( .I1(n13160), .I2(n13163), .O(n463) );
  AND_GATE U621 ( .I1(n464), .I2(n465), .O(n13965) );
  INV_GATE U622 ( .I1(n14412), .O(n466) );
  NAND3_GATE U623 ( .I1(n13132), .I2(n13131), .I3(n13195), .O(n467) );
  OR_GATE U624 ( .I1(n4952), .I2(n4951), .O(n4949) );
  NAND_GATE U625 ( .I1(n13606), .I2(n470), .O(n468) );
  AND_GATE U626 ( .I1(n468), .I2(n469), .O(n13611) );
  OR_GATE U627 ( .I1(n230), .I2(n13608), .O(n469) );
  AND_GATE U628 ( .I1(n13607), .I2(n13609), .O(n470) );
  AND_GATE U629 ( .I1(n7002), .I2(n7001), .O(n471) );
  NOR_GATE U630 ( .I1(n7019), .I2(n278), .O(n472) );
  NOR_GATE U631 ( .I1(n12758), .I2(n13135), .O(n473) );
  NAND_GATE U632 ( .I1(n473), .I2(n474), .O(n476) );
  AND_GATE U633 ( .I1(n13607), .I2(n13133), .O(n474) );
  OR_GATE U634 ( .I1(n12759), .I2(n478), .O(n475) );
  AND_GATE U635 ( .I1(n475), .I2(n476), .O(n12762) );
  INV_GATE U636 ( .I1(n13607), .O(n477) );
  OR_GATE U637 ( .I1(n13133), .I2(n477), .O(n478) );
  AND_GATE U638 ( .I1(n11848), .I2(n11847), .O(n479) );
  NAND_GATE U639 ( .I1(n11853), .I2(n482), .O(n480) );
  AND_GATE U640 ( .I1(n480), .I2(n481), .O(n15352) );
  OR_GATE U641 ( .I1(n1220), .I2(n15350), .O(n481) );
  AND_GATE U642 ( .I1(n11854), .I2(n15351), .O(n482) );
  AND_GATE U643 ( .I1(n11845), .I2(n15351), .O(n483) );
  NAND_GATE U644 ( .I1(n11843), .I2(n486), .O(n484) );
  AND_GATE U645 ( .I1(n484), .I2(n485), .O(n487) );
  OR_GATE U646 ( .I1(n1220), .I2(n11845), .O(n485) );
  AND_GATE U647 ( .I1(n12267), .I2(n15351), .O(n486) );
  OR_GATE U648 ( .I1(n11852), .I2(n487), .O(n1218) );
  OR_GATE U649 ( .I1(n488), .I2(n15356), .O(n12715) );
  AND_GATE U650 ( .I1(n12281), .I2(n12280), .O(n488) );
  NAND_GATE U651 ( .I1(n11852), .I2(n489), .O(n1219) );
  AND_GATE U652 ( .I1(n483), .I2(n11844), .O(n489) );
  NAND_GATE U653 ( .I1(n11414), .I2(n492), .O(n490) );
  AND_GATE U654 ( .I1(n490), .I2(n491), .O(n11419) );
  OR_GATE U655 ( .I1(n11355), .I2(n11416), .O(n491) );
  AND_GATE U656 ( .I1(n621), .I2(n11417), .O(n492) );
  NAND3_GATE U657 ( .I1(n12255), .I2(n12256), .I3(n16), .O(n12259) );
  OR_GATE U658 ( .I1(n15358), .I2(n13149), .O(n13151) );
  AND3_GATE U659 ( .I1(n11388), .I2(n11366), .I3(n11365), .O(n493) );
  NAND_GATE U660 ( .I1(n11841), .I2(n496), .O(n494) );
  AND_GATE U661 ( .I1(n494), .I2(n495), .O(n498) );
  OR_GATE U662 ( .I1(n12271), .I2(n12242), .O(n495) );
  AND_GATE U663 ( .I1(n12243), .I2(n12250), .O(n496) );
  NAND_GATE U664 ( .I1(n11427), .I2(n499), .O(n497) );
  AND_GATE U665 ( .I1(n497), .I2(n498), .O(n12265) );
  AND_GATE U666 ( .I1(n11426), .I2(n12250), .O(n499) );
  OR_GATE U667 ( .I1(n7722), .I2(n858), .O(n7450) );
  OR_GATE U668 ( .I1(n7732), .I2(n500), .O(n7737) );
  AND_GATE U669 ( .I1(n7734), .I2(n7733), .O(n500) );
  OR_GATE U670 ( .I1(n791), .I2(n501), .O(n8322) );
  AND_GATE U671 ( .I1(n8659), .I2(n8662), .O(n501) );
  NAND3_GATE U672 ( .I1(n2782), .I2(n2019), .I3(n2020), .O(n2015) );
  AND3_GATE U673 ( .I1(n10665), .I2(n10370), .I3(n10666), .O(n10866) );
  NAND3_GATE U674 ( .I1(n1879), .I2(n2024), .I3(n1981), .O(n795) );
  NAND4_GATE U675 ( .I1(n2710), .I2(n2724), .I3(n2044), .I4(n2045), .O(n2713)
         );
  NAND3_GATE U676 ( .I1(n13478), .I2(n13479), .I3(n13485), .O(n13697) );
  NAND3_GATE U677 ( .I1(n614), .I2(n5445), .I3(n5721), .O(n5711) );
  NAND3_GATE U678 ( .I1(n10031), .I2(n10032), .I3(n10166), .O(n10173) );
  NAND4_GATE U679 ( .I1(n466), .I2(n13972), .I3(n13970), .I4(n13971), .O(
        n14409) );
  NAND4_GATE U680 ( .I1(n11864), .I2(n11832), .I3(n11831), .I4(n11833), .O(
        n11868) );
  NAND3_GATE U681 ( .I1(n13626), .I2(n13232), .I3(n13233), .O(n13552) );
  AND3_GATE U682 ( .I1(n11528), .I2(n11297), .I3(n11529), .O(n11766) );
  AND3_GATE U683 ( .I1(n13937), .I2(n13938), .I3(n13534), .O(n13646) );
  NAND3_GATE U684 ( .I1(n6090), .I2(n6091), .I3(n6097), .O(n6970) );
  AND3_GATE U685 ( .I1(n12326), .I2(n12335), .I3(n12223), .O(n12336) );
  NAND_GATE U686 ( .I1(n10421), .I2(n10095), .O(n10119) );
  AND_GATE U687 ( .I1(n7065), .I2(n7064), .O(n7809) );
  NAND3_GATE U688 ( .I1(n7461), .I2(n7788), .I3(n7806), .O(n7811) );
  NAND3_GATE U689 ( .I1(n7101), .I2(n7102), .I3(n7108), .O(n7747) );
  AND_GATE U690 ( .I1(n7076), .I2(n7075), .O(n7793) );
  NAND3_GATE U691 ( .I1(n7459), .I2(n7772), .I3(n7790), .O(n7795) );
  AND_GATE U692 ( .I1(n7087), .I2(n7086), .O(n7776) );
  NAND3_GATE U693 ( .I1(n11550), .I2(n11280), .I3(n11551), .O(n11542) );
  AND_GATE U694 ( .I1(n11815), .I2(n11816), .O(n11862) );
  NAND3_GATE U695 ( .I1(n11832), .I2(n11831), .I3(n11833), .O(n666) );
  AND_GATE U696 ( .I1(n6205), .I2(n6204), .O(n6828) );
  NAND4_GATE U697 ( .I1(n14838), .I2(n14502), .I3(n14503), .I4(n14389), .O(
        n14836) );
  NAND3_GATE U698 ( .I1(n13178), .I2(n12751), .I3(n12752), .O(n12706) );
  NAND3_GATE U699 ( .I1(n13155), .I2(n13172), .I3(n13156), .O(n14012) );
  AND_GATE U700 ( .I1(n7474), .I2(n471), .O(n15371) );
  AND3_GATE U701 ( .I1(n3549), .I2(n3550), .I3(n502), .O(n1296) );
  INV_GATE U702 ( .I1(n803), .O(n502) );
  AND_GATE U703 ( .I1(n3563), .I2(n3562), .O(n3944) );
  AND3_GATE U704 ( .I1(n7418), .I2(n7419), .I3(n7440), .O(n7705) );
  NAND3_GATE U705 ( .I1(n10928), .I2(n10929), .I3(n11415), .O(n11416) );
  NAND3_GATE U706 ( .I1(n5808), .I2(n5807), .I3(n6293), .O(n6283) );
  NAND3_GATE U707 ( .I1(n6430), .I2(n5520), .I3(n5519), .O(n5792) );
  AND_GATE U708 ( .I1(n2759), .I2(n2758), .O(n2763) );
  NAND3_GATE U709 ( .I1(n12125), .I2(n12126), .I3(n12132), .O(n12445) );
  AND_GATE U710 ( .I1(n13575), .I2(n13587), .O(n14011) );
  NAND3_GATE U711 ( .I1(n12762), .I2(n467), .I3(n12763), .O(n13139) );
  AND3_GATE U712 ( .I1(n10438), .I2(n10439), .I3(n10539), .O(n10946) );
  AND3_GATE U713 ( .I1(n11428), .I2(n11353), .I3(n11354), .O(n11418) );
  NAND3_GATE U714 ( .I1(n13882), .I2(n13883), .I3(n13889), .O(n14133) );
  OR_GATE U715 ( .I1(n2750), .I2(n2751), .O(n2753) );
  AND3_GATE U716 ( .I1(n13537), .I2(n13538), .I3(n13544), .O(n13647) );
  NAND3_GATE U717 ( .I1(n12300), .I2(n12299), .I3(n12308), .O(n12314) );
  NAND3_GATE U718 ( .I1(n10432), .I2(n10431), .I3(n10528), .O(n10534) );
  NAND3_GATE U719 ( .I1(n14333), .I2(n14334), .I3(n14340), .O(n14590) );
  AND3_GATE U720 ( .I1(n13074), .I2(n13075), .I3(n13081), .O(n13260) );
  NAND4_GATE U721 ( .I1(n13269), .I2(n13067), .I3(n13066), .I4(n13271), .O(
        n13277) );
  NAND3_GATE U722 ( .I1(n13045), .I2(n13046), .I3(n13052), .O(n13280) );
  NAND3_GATE U723 ( .I1(n13523), .I2(n13524), .I3(n13530), .O(n13656) );
  NAND5_GATE U724 ( .I1(n5317), .I2(n5318), .I3(n5337), .I4(n4872), .I5(n5338), 
        .O(n5323) );
  NAND3_GATE U725 ( .I1(n3819), .I2(n3815), .I3(n3816), .O(n3898) );
  AND3_GATE U726 ( .I1(n13521), .I2(n13522), .I3(n13071), .O(n13259) );
  AND_GATE U727 ( .I1(n2814), .I2(n3011), .O(n1150) );
  NAND4_GATE U728 ( .I1(n13268), .I2(n13505), .I3(n13506), .I4(n13056), .O(
        n13272) );
  AND3_GATE U729 ( .I1(n11923), .I2(n11775), .I3(n11924), .O(n12188) );
  NAND3_GATE U730 ( .I1(n13551), .I2(n13232), .I3(n13233), .O(n13627) );
  NAND4_GATE U731 ( .I1(n13535), .I2(n13536), .I3(n13085), .I4(n13248), .O(
        n13246) );
  AND_GATE U732 ( .I1(n14063), .I2(n13962), .O(n14062) );
  NAND4_GATE U733 ( .I1(n12721), .I2(n12289), .I3(n12290), .I4(n12291), .O(
        n12725) );
  NAND3_GATE U734 ( .I1(n3038), .I2(n3039), .I3(n3567), .O(n3565) );
  NAND4_GATE U735 ( .I1(n3570), .I2(n3574), .I3(n3023), .I4(n3024), .O(n3566)
         );
  NAND3_GATE U736 ( .I1(n9581), .I2(n846), .I3(n845), .O(n9582) );
  NAND3_GATE U737 ( .I1(n6824), .I2(n657), .I3(n656), .O(n6825) );
  AND_GATE U738 ( .I1(n7109), .I2(n7108), .O(n7745) );
  NAND4_GATE U739 ( .I1(n15363), .I2(n14007), .I3(n14008), .I4(n14009), .O(
        n14020) );
  NAND3_GATE U740 ( .I1(n13215), .I2(n13113), .I3(n13114), .O(n13218) );
  NAND3_GATE U741 ( .I1(n13125), .I2(n13214), .I3(n13126), .O(n13219) );
  AND3_GATE U742 ( .I1(n14390), .I2(n14391), .I3(n13950), .O(n14067) );
  AND3_GATE U743 ( .I1(n12796), .I2(n12675), .I3(n12797), .O(n13090) );
  NAND3_GATE U744 ( .I1(n9829), .I2(n9830), .I3(n9841), .O(n10163) );
  AND_GATE U745 ( .I1(n11314), .I2(n11803), .O(n11493) );
  NAND3_GATE U746 ( .I1(n7661), .I2(n7358), .I3(n7659), .O(n8232) );
  NAND3_GATE U747 ( .I1(n8403), .I2(n8248), .I3(n8404), .O(n8396) );
  NAND3_GATE U748 ( .I1(n7350), .I2(n7356), .I3(n7648), .O(n7654) );
  AND3_GATE U749 ( .I1(n12352), .I2(n12220), .I3(n12221), .O(n12341) );
  NAND3_GATE U750 ( .I1(n12337), .I2(n1231), .I3(n1230), .O(n12334) );
  AND3_GATE U751 ( .I1(n10145), .I2(n10061), .I3(n10062), .O(n10393) );
  AND_GATE U752 ( .I1(n12784), .I2(n13123), .O(n12791) );
  NAND4_GATE U753 ( .I1(n13127), .I2(n13215), .I3(n13113), .I4(n13114), .O(
        n13222) );
  AND3_GATE U754 ( .I1(n7660), .I2(n7359), .I3(n7658), .O(n7509) );
  NAND3_GATE U755 ( .I1(n3000), .I2(n3002), .I3(n3003), .O(n3001) );
  AND_GATE U756 ( .I1(n9213), .I2(n9560), .O(n9577) );
  NAND4_GATE U757 ( .I1(n11522), .I2(n11301), .I3(n11523), .I4(n11780), .O(
        n11778) );
  NAND4_GATE U758 ( .I1(n13127), .I2(n13125), .I3(n13214), .I4(n13126), .O(
        n13221) );
  AND3_GATE U759 ( .I1(n13221), .I2(n13222), .I3(n13217), .O(n13977) );
  AND_GATE U760 ( .I1(n1139), .I2(n3904), .O(n3908) );
  NAND4_GATE U761 ( .I1(n9547), .I2(n8871), .I3(n8873), .I4(n8872), .O(n9544)
         );
  AND3_GATE U762 ( .I1(n11515), .I2(n11516), .I3(n11517), .O(n12210) );
  NAND3_GATE U763 ( .I1(n10171), .I2(n10033), .I3(n10167), .O(n10176) );
  AND_GATE U764 ( .I1(n12691), .I2(n13102), .O(n13118) );
  NAND3_GATE U765 ( .I1(n4790), .I2(n4794), .I3(n5397), .O(n5402) );
  AND_GATE U766 ( .I1(n3001), .I2(n3004), .O(n1034) );
  AND_GATE U767 ( .I1(n4643), .I2(n4642), .O(n4859) );
  AND3_GATE U768 ( .I1(n8018), .I2(n8019), .I3(n8020), .O(n8635) );
  AND3_GATE U769 ( .I1(n7921), .I2(n7922), .I3(n7928), .O(n8737) );
  NAND3_GATE U770 ( .I1(n8330), .I2(n8716), .I3(n8734), .O(n8739) );
  AND3_GATE U771 ( .I1(n7931), .I2(n7932), .I3(n7938), .O(n8721) );
  NAND3_GATE U772 ( .I1(n8328), .I2(n8700), .I3(n8718), .O(n8723) );
  AND_GATE U773 ( .I1(n7949), .I2(n7948), .O(n8705) );
  AND_GATE U774 ( .I1(n8815), .I2(n8814), .O(n9622) );
  NAND3_GATE U775 ( .I1(n9219), .I2(n9601), .I3(n9619), .O(n9624) );
  NAND3_GATE U776 ( .I1(n10113), .I2(n9661), .I3(n9660), .O(n15334) );
  AND3_GATE U777 ( .I1(n6567), .I2(n6568), .I3(n6569), .O(n7188) );
  AND_GATE U778 ( .I1(n15099), .I2(n14817), .O(n15077) );
  NAND3_GATE U779 ( .I1(n11126), .I2(n11127), .I3(n11133), .O(n11586) );
  NAND4_GATE U780 ( .I1(n10491), .I2(n10493), .I3(n9672), .I4(n9671), .O(
        n15338) );
  AND3_GATE U781 ( .I1(n11031), .I2(n11032), .I3(n11033), .O(n11797) );
  AND3_GATE U782 ( .I1(n13142), .I2(n13143), .I3(n13141), .O(n13164) );
  NAND3_GATE U783 ( .I1(n10159), .I2(n10152), .I3(n10153), .O(n10881) );
  AND_GATE U784 ( .I1(n14400), .I2(n14399), .O(n14839) );
  NAND3_GATE U785 ( .I1(n13939), .I2(n13940), .I3(n13946), .O(n14080) );
  NAND4_GATE U786 ( .I1(n14432), .I2(n13623), .I3(n13624), .I4(n13625), .O(
        n14424) );
  AND3_GATE U787 ( .I1(n6698), .I2(n6699), .I3(n6700), .O(n7353) );
  AND3_GATE U788 ( .I1(n14499), .I2(n14500), .I3(n14501), .O(n14956) );
  NAND3_GATE U789 ( .I1(n14964), .I2(n14851), .I3(n14946), .O(n14862) );
  AND3_GATE U790 ( .I1(n14496), .I2(n14498), .I3(n14404), .O(n14855) );
  NAND5_GATE U791 ( .I1(n13981), .I2(n13221), .I3(n13222), .I4(n13976), .I5(
        n13217), .O(n13986) );
  NAND3_GATE U792 ( .I1(n13896), .I2(n13897), .I3(n13903), .O(n14118) );
  NAND3_GATE U793 ( .I1(n13951), .I2(n13952), .I3(n13548), .O(n13634) );
  NAND3_GATE U794 ( .I1(n14034), .I2(n13990), .I3(n14424), .O(n14040) );
  NAND3_GATE U795 ( .I1(n6100), .I2(n6101), .I3(n6115), .O(n6958) );
  AND_GATE U796 ( .I1(n8324), .I2(n8667), .O(n8688) );
  AND3_GATE U797 ( .I1(n11329), .I2(n11330), .I3(n11490), .O(n11477) );
  NAND3_GATE U798 ( .I1(n8081), .I2(n8082), .I3(n8089), .O(n8411) );
  AND_GATE U799 ( .I1(n2911), .I2(n2910), .O(n2915) );
  AND_GATE U800 ( .I1(n4819), .I2(n4820), .O(n5525) );
  NAND5_GATE U801 ( .I1(n7682), .I2(n7684), .I3(n7380), .I4(n7381), .I5(n7382), 
        .O(n8258) );
  AND_GATE U802 ( .I1(n12746), .I2(n12745), .O(n13159) );
  NAND3_GATE U803 ( .I1(n462), .I2(n13162), .I3(n13158), .O(n13166) );
  AND3_GATE U804 ( .I1(n8851), .I2(n8852), .I3(n8861), .O(n630) );
  AND_GATE U805 ( .I1(n10107), .I2(n10450), .O(n10464) );
  NAND3_GATE U806 ( .I1(n8851), .I2(n8852), .I3(n8861), .O(n9564) );
  NAND3_GATE U807 ( .I1(n5203), .I2(n5204), .I3(n5210), .O(n5996) );
  AND_GATE U808 ( .I1(n7971), .I2(n7970), .O(n8672) );
  NAND5_GATE U809 ( .I1(n503), .I2(n10463), .I3(n9690), .I4(n9691), .I5(n9692), 
        .O(n10504) );
  INV_GATE U810 ( .I1(n10506), .O(n503) );
  AND3_GATE U811 ( .I1(n11913), .I2(n11792), .I3(n11914), .O(n12207) );
  NAND3_GATE U812 ( .I1(n12216), .I2(n12217), .I3(n12369), .O(n12361) );
  NAND3_GATE U813 ( .I1(n12300), .I2(n12306), .I3(n12299), .O(n12312) );
  NAND3_GATE U814 ( .I1(n8394), .I2(n8393), .I3(n8588), .O(n8952) );
  NAND_GATE U815 ( .I1(n10925), .I2(n10926), .O(n11435) );
  NAND3_GATE U816 ( .I1(n10458), .I2(n1208), .I3(n1209), .O(n10459) );
  NAND3_GATE U817 ( .I1(n10459), .I2(n10460), .I3(n10523), .O(n10980) );
  AND3_GATE U818 ( .I1(n13216), .I2(n13213), .I3(n13128), .O(n13204) );
  NAND_GATE U819 ( .I1(n10097), .I2(n10098), .O(n10433) );
  NAND4_GATE U820 ( .I1(n504), .I2(n8955), .I3(n8959), .I4(n8958), .O(n9269)
         );
  INV_GATE U821 ( .I1(n9817), .O(n504) );
  NAND3_GATE U822 ( .I1(n10990), .I2(n11437), .I3(n11434), .O(n11445) );
  NAND4_GATE U823 ( .I1(n10461), .I2(n10459), .I3(n10460), .I4(n10523), .O(
        n10977) );
  AND3_GATE U824 ( .I1(n10462), .I2(n10522), .I3(n10521), .O(n10514) );
  AND_GATE U825 ( .I1(n8804), .I2(n8803), .O(n9638) );
  NAND3_GATE U826 ( .I1(n9221), .I2(n9617), .I3(n9635), .O(n9640) );
  NAND4_GATE U827 ( .I1(n14001), .I2(n14034), .I3(n13990), .I4(n14424), .O(
        n14038) );
  AND_GATE U828 ( .I1(n11432), .I2(n11431), .O(n11449) );
  AND_GATE U829 ( .I1(n10931), .I2(n10932), .O(n11362) );
  NAND3_GATE U830 ( .I1(n7715), .I2(n7714), .I3(n8013), .O(n8002) );
  NAND3_GATE U831 ( .I1(n10461), .I2(n10525), .I3(n10524), .O(n10976) );
  AND3_GATE U832 ( .I1(n8391), .I2(n8390), .I3(n8392), .O(n9161) );
  NAND5_GATE U833 ( .I1(n14376), .I2(n555), .I3(n554), .I4(n536), .I5(n535), 
        .O(n14081) );
  NAND3_GATE U834 ( .I1(n14001), .I2(n14033), .I3(n604), .O(n14037) );
  AND3_GATE U835 ( .I1(n9734), .I2(n9726), .I3(n9727), .O(n10434) );
  AND3_GATE U836 ( .I1(n8406), .I2(n8407), .I3(n8408), .O(n9139) );
  NAND3_GATE U837 ( .I1(n11355), .I2(n11416), .I3(n11413), .O(n11420) );
  NAND3_GATE U838 ( .I1(n2784), .I2(n2951), .I3(n2783), .O(n2960) );
  AND3_GATE U839 ( .I1(n12312), .I2(n12734), .I3(n12311), .O(n1213) );
  NAND4_GATE U840 ( .I1(n5356), .I2(n4847), .I3(n5359), .I4(n5366), .O(n5550)
         );
  NAND3_GATE U841 ( .I1(n11093), .I2(n11094), .I3(n11100), .O(n11563) );
  AND3_GATE U842 ( .I1(n9193), .I2(n9194), .I3(n9195), .O(n9505) );
  NAND3_GATE U843 ( .I1(n9503), .I2(n9509), .I3(n9792), .O(n9780) );
  AND3_GATE U844 ( .I1(n9793), .I2(n9794), .I3(n9795), .O(n10123) );
  NAND3_GATE U845 ( .I1(n10339), .I2(n10340), .I3(n10346), .O(n10705) );
  NAND3_GATE U846 ( .I1(n10491), .I2(n10488), .I3(n15338), .O(n10496) );
  NAND3_GATE U847 ( .I1(n13953), .I2(n13954), .I3(n13960), .O(n14066) );
  NAND3_GATE U848 ( .I1(n13537), .I2(n13538), .I3(n13544), .O(n13645) );
  NAND3_GATE U849 ( .I1(n13074), .I2(n13075), .I3(n13081), .O(n13258) );
  NAND3_GATE U850 ( .I1(n8986), .I2(n8987), .I3(n8993), .O(n9445) );
  AND3_GATE U851 ( .I1(n9499), .I2(n9500), .I3(n9802), .O(n10068) );
  AND3_GATE U852 ( .I1(n8943), .I2(n8944), .I3(n8945), .O(n9494) );
  NAND3_GATE U853 ( .I1(n14859), .I2(n841), .I3(n840), .O(n14860) );
  AND_GATE U854 ( .I1(n15070), .I2(n14821), .O(n15048) );
  AND3_GATE U855 ( .I1(n14871), .I2(n14872), .I3(n14873), .O(n14932) );
  NAND4_GATE U856 ( .I1(n12768), .I2(n12356), .I3(n12355), .I4(n12357), .O(
        n12772) );
  OR3_GATE U857 ( .I1(n13558), .I2(n13991), .I3(n13200), .O(n13996) );
  AND3_GATE U858 ( .I1(n9249), .I2(n9250), .I3(n9251), .O(n10067) );
  NAND3_GATE U859 ( .I1(n11008), .I2(n10914), .I3(n678), .O(n1235) );
  NAND3_GATE U860 ( .I1(n13178), .I2(n12750), .I3(n13185), .O(n13189) );
  AND3_GATE U861 ( .I1(n13627), .I2(n13629), .I3(n13552), .O(n13978) );
  AND3_GATE U862 ( .I1(n13988), .I2(n14047), .I3(n14049), .O(n14429) );
  NAND3_GATE U863 ( .I1(n7204), .I2(n6704), .I3(n7202), .O(n7206) );
  NAND3_GATE U864 ( .I1(n11552), .I2(n11553), .I3(n11559), .O(n11950) );
  NAND3_GATE U865 ( .I1(n11936), .I2(n11937), .I3(n11946), .O(n12409) );
  AND_GATE U866 ( .I1(n13996), .I2(n13564), .O(n13612) );
  AND3_GATE U867 ( .I1(n1305), .I2(n14453), .I3(n15365), .O(\A2[32] ) );
  NAND3_GATE U868 ( .I1(n6597), .I2(n6594), .I3(n6595), .O(n6601) );
  AND3_GATE U869 ( .I1(n9829), .I2(n9830), .I3(n9841), .O(n1328) );
  NAND3_GATE U870 ( .I1(n12795), .I2(n12780), .I3(n12781), .O(n13205) );
  AND3_GATE U871 ( .I1(n7540), .I2(n7326), .I3(n7541), .O(n917) );
  NAND3_GATE U872 ( .I1(n5270), .I2(n5271), .I3(n5277), .O(n5622) );
  NAND3_GATE U873 ( .I1(n10696), .I2(n10697), .I3(n10703), .O(n11102) );
  AND_GATE U874 ( .I1(n9672), .I2(n9671), .O(n10487) );
  OR_GATE U875 ( .I1(n8399), .I2(n772), .O(n8404) );
  NAND3_GATE U876 ( .I1(n11449), .I2(n12235), .I3(n12231), .O(n12242) );
  AND_GATE U877 ( .I1(A[0]), .I2(A[1]), .O(n1196) );
  AND_GATE U878 ( .I1(n1858), .I2(n1859), .O(n1297) );
  AND_GATE U879 ( .I1(n6377), .I2(n6376), .O(n6680) );
  AND_GATE U880 ( .I1(n5424), .I2(n5425), .O(n5682) );
  NAND3_GATE U881 ( .I1(n11915), .I2(n11916), .I3(n11922), .O(n12680) );
  NAND3_GATE U882 ( .I1(n3552), .I2(n3553), .I3(n3059), .O(n818) );
  NAND3_GATE U883 ( .I1(n6505), .I2(n6511), .I3(n6504), .O(n6801) );
  NAND5_GATE U884 ( .I1(n10672), .I2(n10200), .I3(n10202), .I4(n10675), .I5(
        n10201), .O(n10682) );
  NAND3_GATE U885 ( .I1(n12250), .I2(n12249), .I3(n12266), .O(n12274) );
  AND3_GATE U886 ( .I1(n15356), .I2(n12281), .I3(n12280), .O(\A2[36] ) );
  NAND3_GATE U887 ( .I1(n7988), .I2(n7989), .I3(n8001), .O(n8642) );
  AND3_GATE U888 ( .I1(n8616), .I2(n8311), .I3(n8312), .O(n8343) );
  NAND3_GATE U889 ( .I1(n8340), .I2(n8339), .I3(n8628), .O(n8893) );
  NAND3_GATE U890 ( .I1(n9695), .I2(n9696), .I3(n9705), .O(n10456) );
  NAND4_GATE U891 ( .I1(n1220), .I2(n11854), .I3(n11406), .I4(n11405), .O(
        n15354) );
  NAND3_GATE U892 ( .I1(n7703), .I2(n7708), .I3(n8042), .O(n8046) );
  NAND3_GATE U893 ( .I1(n504), .I2(n9274), .I3(n9822), .O(n9809) );
  AND3_GATE U894 ( .I1(n8034), .I2(n7713), .I3(n8031), .O(n8015) );
  AND_GATE U895 ( .I1(n9208), .I2(n9209), .O(n9551) );
  AND3_GATE U896 ( .I1(n9543), .I2(n9724), .I3(n9732), .O(n9711) );
  AND3_GATE U897 ( .I1(n11365), .I2(n11366), .I3(n11388), .O(n11379) );
  NAND3_GATE U898 ( .I1(n7112), .I2(n7113), .I3(n7119), .O(n7734) );
  AND_GATE U899 ( .I1(n2009), .I2(n2010), .O(n1193) );
  NAND3_GATE U900 ( .I1(n10590), .I2(n10599), .I3(n10591), .O(n11003) );
  NAND5_GATE U901 ( .I1(n262), .I2(n5357), .I3(n1151), .I4(n5368), .I5(n5381), 
        .O(n5549) );
  AND3_GATE U902 ( .I1(n5370), .I2(n5549), .I3(n5550), .O(n5810) );
  AND3_GATE U903 ( .I1(n10581), .I2(n10579), .I3(n10580), .O(n10997) );
  AND_GATE U904 ( .I1(n7677), .I2(n7676), .O(n8065) );
  AND3_GATE U905 ( .I1(n11868), .I2(n11835), .I3(n11836), .O(n12293) );
  AND_GATE U906 ( .I1(n5396), .I2(n5395), .O(n5772) );
  NAND3_GATE U907 ( .I1(n8064), .I2(n8068), .I3(n8378), .O(n8384) );
  AND3_GATE U908 ( .I1(n8266), .I2(n8267), .I3(n8268), .O(n8365) );
  AND3_GATE U909 ( .I1(n8356), .I2(n8355), .I3(n8357), .O(n9172) );
  NAND3_GATE U910 ( .I1(n10381), .I2(n10385), .I3(n10640), .O(n10631) );
  NAND3_GATE U911 ( .I1(n4822), .I2(n4821), .I3(n5516), .O(n5524) );
  AND_GATE U912 ( .I1(n2948), .I2(n2949), .O(n3645) );
  NAND3_GATE U913 ( .I1(n11079), .I2(n11080), .I3(n11090), .O(n11541) );
  NAND3_GATE U914 ( .I1(n8877), .I2(n8878), .I3(n8890), .O(n9538) );
  NAND3_GATE U915 ( .I1(n8455), .I2(n8456), .I3(n8462), .O(n9093) );
  NAND3_GATE U916 ( .I1(n8053), .I2(n8061), .I3(n8054), .O(n8608) );
  AND_GATE U917 ( .I1(n15042), .I2(n14825), .O(n15021) );
  NAND3_GATE U918 ( .I1(n7921), .I2(n7922), .I3(n7928), .O(n8734) );
  NAND3_GATE U919 ( .I1(n7931), .I2(n7932), .I3(n7938), .O(n8718) );
  NAND3_GATE U920 ( .I1(n10205), .I2(n10206), .I3(n10212), .O(n10849) );
  NAND3_GATE U921 ( .I1(n4399), .I2(n4400), .I3(n4406), .O(n4922) );
  NAND3_GATE U922 ( .I1(n4389), .I2(n4390), .I3(n4396), .O(n4938) );
  NAND3_GATE U923 ( .I1(n5310), .I2(n5311), .I3(n5324), .O(n5834) );
  AND_GATE U924 ( .I1(n10160), .I2(n10159), .O(n505) );
  AND3_GATE U925 ( .I1(n13557), .I2(n13620), .I3(n13621), .O(n506) );
  AND3_GATE U926 ( .I1(n12394), .I2(n12183), .I3(n12393), .O(n507) );
  AND_GATE U927 ( .I1(n10846), .I2(n10352), .O(n508) );
  OR_GATE U928 ( .I1(n1032), .I2(n511), .O(n509) );
  AND_GATE U929 ( .I1(n509), .I2(n510), .O(n10191) );
  OR_GATE U930 ( .I1(n10195), .I2(n10353), .O(n510) );
  OR_GATE U931 ( .I1(n10354), .I2(n10195), .O(n511) );
  AND_GATE U932 ( .I1(n13139), .I2(n13173), .O(n512) );
  AND_GATE U933 ( .I1(n9544), .I2(n9211), .O(n513) );
  AND3_GATE U934 ( .I1(n13566), .I2(n13565), .I3(n13610), .O(n514) );
  NAND_GATE U935 ( .I1(n10361), .I2(n517), .O(n515) );
  AND_GATE U936 ( .I1(n515), .I2(n516), .O(n10683) );
  OR_GATE U937 ( .I1(n10689), .I2(n10364), .O(n516) );
  AND_GATE U938 ( .I1(n10362), .I2(n10365), .O(n517) );
  NAND_GATE U939 ( .I1(n6388), .I2(n6387), .O(n518) );
  AND3_GATE U940 ( .I1(n8995), .I2(n519), .I3(n8994), .O(n768) );
  NAND_GATE U941 ( .I1(n8999), .I2(n8998), .O(n519) );
  AND_GATE U942 ( .I1(n520), .I2(n521), .O(n14879) );
  OR_GATE U943 ( .I1(n14886), .I2(n14478), .O(n521) );
  AND_GATE U944 ( .I1(n12162), .I2(n12161), .O(n522) );
  OR_GATE U945 ( .I1(n9139), .I2(n9149), .O(n9144) );
  AND3_GATE U946 ( .I1(n13138), .I2(n12761), .I3(n13137), .O(n523) );
  NOR_GATE U947 ( .I1(n1355), .I2(n1047), .O(n524) );
  AND_GATE U948 ( .I1(n12358), .I2(n12219), .O(n525) );
  AND_GATE U949 ( .I1(n7644), .I2(n7643), .O(n526) );
  AND_GATE U950 ( .I1(n6388), .I2(n6387), .O(n527) );
  NAND_GATE U951 ( .I1(n1311), .I2(n531), .O(n529) );
  AND_GATE U952 ( .I1(n529), .I2(n530), .O(n4470) );
  OR_GATE U953 ( .I1(n4600), .I2(n4468), .O(n530) );
  AND_GATE U954 ( .I1(n4590), .I2(n4608), .O(n531) );
  NAND_GATE U955 ( .I1(n12424), .I2(n534), .O(n532) );
  AND_GATE U956 ( .I1(n532), .I2(n533), .O(n13057) );
  OR_GATE U957 ( .I1(n13063), .I2(n12427), .O(n533) );
  AND_GATE U958 ( .I1(n12425), .I2(n12642), .O(n534) );
  NAND_GATE U959 ( .I1(n13665), .I2(n537), .O(n535) );
  OR_GATE U960 ( .I1(n14381), .I2(n13668), .O(n536) );
  AND_GATE U961 ( .I1(n13666), .I2(n13936), .O(n537) );
  NAND_GATE U962 ( .I1(n9611), .I2(n540), .O(n538) );
  AND_GATE U963 ( .I1(n538), .I2(n539), .O(n9662) );
  OR_GATE U964 ( .I1(n9668), .I2(n9614), .O(n539) );
  AND_GATE U965 ( .I1(n9612), .I2(n9615), .O(n540) );
  AND_GATE U966 ( .I1(n5844), .I2(n5566), .O(n541) );
  NAND_GATE U967 ( .I1(n13274), .I2(n544), .O(n542) );
  AND_GATE U968 ( .I1(n542), .I2(n543), .O(n13923) );
  OR_GATE U969 ( .I1(n13929), .I2(n13277), .O(n543) );
  AND_GATE U970 ( .I1(n13275), .I2(n13519), .O(n544) );
  AND3_GATE U971 ( .I1(n5306), .I2(n5305), .I3(n5304), .O(n545) );
  NAND_GATE U972 ( .I1(n8678), .I2(n548), .O(n546) );
  AND_GATE U973 ( .I1(n546), .I2(n547), .O(n8838) );
  OR_GATE U974 ( .I1(n8844), .I2(n8681), .O(n547) );
  AND_GATE U975 ( .I1(n8679), .I2(n8682), .O(n548) );
  NOR_GATE U976 ( .I1(n3889), .I2(n3888), .O(n549) );
  AND_GATE U977 ( .I1(n12654), .I2(n12653), .O(n550) );
  AND_GATE U978 ( .I1(n7700), .I2(n7699), .O(n551) );
  AND_GATE U979 ( .I1(n9873), .I2(n9872), .O(n552) );
  AND_GATE U980 ( .I1(n6629), .I2(n6628), .O(n553) );
  NAND_GATE U981 ( .I1(n13665), .I2(n557), .O(n554) );
  OR_GATE U982 ( .I1(n556), .I2(n13668), .O(n555) );
  INV_GATE U983 ( .I1(n14380), .O(n556) );
  AND_GATE U984 ( .I1(n13666), .I2(n14380), .O(n557) );
  NAND_GATE U985 ( .I1(n8742), .I2(n560), .O(n558) );
  AND_GATE U986 ( .I1(n558), .I2(n559), .O(n8794) );
  OR_GATE U987 ( .I1(n8800), .I2(n8745), .O(n559) );
  AND_GATE U988 ( .I1(n8743), .I2(n8746), .O(n560) );
  NAND_GATE U989 ( .I1(n8726), .I2(n563), .O(n561) );
  AND_GATE U990 ( .I1(n561), .I2(n562), .O(n8805) );
  OR_GATE U991 ( .I1(n8811), .I2(n8729), .O(n562) );
  AND_GATE U992 ( .I1(n8727), .I2(n8730), .O(n563) );
  AND_GATE U993 ( .I1(n5267), .I2(n5266), .O(n564) );
  AND_GATE U994 ( .I1(n10037), .I2(n10036), .O(n565) );
  AND3_GATE U995 ( .I1(n10172), .I2(n10177), .I3(n10176), .O(n566) );
  AND3_GATE U996 ( .I1(n10168), .I2(n10034), .I3(n10170), .O(n567) );
  AND3_GATE U997 ( .I1(n14002), .I2(n14032), .I3(n14035), .O(n568) );
  AND_GATE U998 ( .I1(n10098), .I2(n10097), .O(n569) );
  NAND_GATE U999 ( .I1(n9627), .I2(n572), .O(n570) );
  AND_GATE U1000 ( .I1(n570), .I2(n571), .O(n9651) );
  OR_GATE U1001 ( .I1(n9657), .I2(n9630), .O(n571) );
  AND_GATE U1002 ( .I1(n9628), .I2(n9631), .O(n572) );
  AND3_GATE U1003 ( .I1(n2946), .I2(n2945), .I3(n2944), .O(n573) );
  AND_GATE U1004 ( .I1(n4839), .I2(n4838), .O(n574) );
  AND_GATE U1005 ( .I1(B[31]), .I2(B[30]), .O(n1192) );
  AND_GATE U1006 ( .I1(n6584), .I2(n6583), .O(n575) );
  AND_GATE U1007 ( .I1(n10045), .I2(n10044), .O(n576) );
  NAND_GATE U1008 ( .I1(n12787), .I2(n579), .O(n577) );
  AND_GATE U1009 ( .I1(n577), .I2(n578), .O(n12694) );
  OR_GATE U1010 ( .I1(n12786), .I2(n12782), .O(n578) );
  AND_GATE U1011 ( .I1(n12785), .I2(n12778), .O(n579) );
  NAND_GATE U1012 ( .I1(n4431), .I2(n582), .O(n580) );
  AND_GATE U1013 ( .I1(n580), .I2(n581), .O(n4408) );
  OR_GATE U1014 ( .I1(n4418), .I2(n3960), .O(n581) );
  AND_GATE U1015 ( .I1(n4425), .I2(n3968), .O(n582) );
  AND_GATE U1016 ( .I1(n5278), .I2(n5277), .O(n583) );
  AND_GATE U1017 ( .I1(n3976), .I2(n3975), .O(n584) );
  AND_GATE U1018 ( .I1(n10929), .I2(n10928), .O(n585) );
  NAND_GATE U1019 ( .I1(n586), .I2(n8096), .O(n8094) );
  NOR_GATE U1020 ( .I1(n8099), .I2(n8095), .O(n586) );
  NAND_GATE U1021 ( .I1(n5444), .I2(n587), .O(n613) );
  NOR_GATE U1022 ( .I1(n5443), .I2(n614), .O(n587) );
  AND_GATE U1023 ( .I1(n9535), .I2(n9539), .O(n588) );
  AND_GATE U1024 ( .I1(n11449), .I2(n12231), .O(n589) );
  AND_GATE U1025 ( .I1(n8305), .I2(n8304), .O(n590) );
  AND3_GATE U1026 ( .I1(n11908), .I2(n11809), .I3(n11907), .O(n591) );
  AND_GATE U1027 ( .I1(n14027), .I2(n14006), .O(n592) );
  AND_GATE U1028 ( .I1(n12242), .I2(n11842), .O(n593) );
  AND3_GATE U1029 ( .I1(n10430), .I2(n10429), .I3(n10555), .O(n594) );
  AND3_GATE U1030 ( .I1(n5636), .I2(n5544), .I3(n5543), .O(n595) );
  AND_GATE U1031 ( .I1(n7414), .I2(n7413), .O(n596) );
  AND_GATE U1032 ( .I1(n7704), .I2(n7443), .O(n597) );
  NAND_GATE U1033 ( .I1(n14877), .I2(n598), .O(n14891) );
  AND_GATE U1034 ( .I1(n13986), .I2(n13985), .O(n599) );
  NAND3_GATE U1035 ( .I1(n4628), .I2(n4627), .I3(n4626), .O(n600) );
  AND_GATE U1036 ( .I1(n14466), .I2(n14442), .O(n601) );
  AND_GATE U1037 ( .I1(n11346), .I2(n11345), .O(n602) );
  AND3_GATE U1038 ( .I1(n10150), .I2(n10149), .I3(n10148), .O(n603) );
  AND_GATE U1039 ( .I1(n14000), .I2(n13999), .O(n604) );
  AND_GATE U1040 ( .I1(n11538), .I2(n11537), .O(n605) );
  AND_GATE U1041 ( .I1(n12744), .I2(n12743), .O(n606) );
  AND_GATE U1042 ( .I1(n7561), .I2(n7560), .O(n607) );
  OR_GATE U1043 ( .I1(n3901), .I2(n1304), .O(n608) );
  AND_GATE U1044 ( .I1(n4605), .I2(n4604), .O(n609) );
  OR_GATE U1045 ( .I1(n1397), .I2(B[30]), .O(n1933) );
  AND_GATE U1046 ( .I1(n3584), .I2(n3583), .O(n610) );
  AND_GATE U1047 ( .I1(n12772), .I2(n12696), .O(n611) );
  OR_GATE U1048 ( .I1(n5444), .I2(n615), .O(n612) );
  AND_GATE U1049 ( .I1(n612), .I2(n613), .O(n5447) );
  INV_GATE U1050 ( .I1(n5719), .O(n614) );
  OR_GATE U1051 ( .I1(n714), .I2(n614), .O(n615) );
  AND_GATE U1052 ( .I1(n3714), .I2(n3713), .O(n616) );
  AND_GATE U1053 ( .I1(n8826), .I2(n8825), .O(n617) );
  NAND_GATE U1054 ( .I1(n6816), .I2(n6515), .O(n618) );
  NOR_GATE U1055 ( .I1(n5384), .I2(n5388), .O(n619) );
  AND_GATE U1056 ( .I1(n861), .I2(n3661), .O(n620) );
  AND3_GATE U1057 ( .I1(n10543), .I2(n10542), .I3(n10541), .O(n621) );
  AND_GATE U1058 ( .I1(n11845), .I2(n11844), .O(n622) );
  AND_GATE U1059 ( .I1(n11427), .I2(n11426), .O(n623) );
  AND_GATE U1060 ( .I1(n12706), .I2(n12705), .O(n624) );
  AND_GATE U1061 ( .I1(n11933), .I2(n11932), .O(n625) );
  AND3_GATE U1062 ( .I1(n14870), .I2(n14868), .I3(n14421), .O(n626) );
  AND3_GATE U1063 ( .I1(n11934), .I2(n11758), .I3(n11935), .O(n627) );
  AND_GATE U1064 ( .I1(n14491), .I2(n14490), .O(n628) );
  AND_GATE U1065 ( .I1(n11947), .I2(n11946), .O(n629) );
  AND_GATE U1066 ( .I1(n6779), .I2(n6778), .O(n631) );
  INV_GATE U1067 ( .I1(n631), .O(n7141) );
  AND3_GATE U1068 ( .I1(n9286), .I2(n9125), .I3(n9285), .O(n632) );
  OR_GATE U1069 ( .I1(n632), .I2(n9470), .O(n9472) );
  NOR_GATE U1070 ( .I1(n10850), .I2(n695), .O(n696) );
  AND_GATE U1071 ( .I1(n9338), .I2(n9337), .O(n633) );
  INV_GATE U1072 ( .I1(n633), .O(n9973) );
  OR_GATE U1073 ( .I1(n467), .I2(n523), .O(n13192) );
  AND_GATE U1074 ( .I1(n4840), .I2(n4844), .O(n634) );
  INV_GATE U1075 ( .I1(n634), .O(n5377) );
  NAND_GATE U1076 ( .I1(n11120), .I2(n638), .O(n635) );
  AND_GATE U1077 ( .I1(n635), .I2(n636), .O(n11728) );
  OR_GATE U1078 ( .I1(n637), .I2(n11122), .O(n636) );
  INV_GATE U1079 ( .I1(n11123), .O(n637) );
  AND_GATE U1080 ( .I1(n11121), .I2(n11123), .O(n638) );
  NAND_GATE U1081 ( .I1(n10231), .I2(n641), .O(n639) );
  AND_GATE U1082 ( .I1(n639), .I2(n640), .O(n10234) );
  OR_GATE U1083 ( .I1(n10229), .I2(n10232), .O(n640) );
  AND_GATE U1084 ( .I1(n10230), .I2(n10233), .O(n641) );
  NAND_GATE U1085 ( .I1(n642), .I2(n12617), .O(n12616) );
  NOR_GATE U1086 ( .I1(n12618), .I2(n12619), .O(n642) );
  NAND_GATE U1087 ( .I1(n643), .I2(n8131), .O(n8130) );
  NOR_GATE U1088 ( .I1(n8133), .I2(n8132), .O(n643) );
  AND_GATE U1089 ( .I1(n14355), .I2(n14354), .O(n644) );
  NAND_GATE U1090 ( .I1(n14862), .I2(n14950), .O(n645) );
  NAND_GATE U1091 ( .I1(n645), .I2(n646), .O(n14874) );
  AND_GATE U1092 ( .I1(n14831), .I2(n15001), .O(n647) );
  AND_GATE U1093 ( .I1(n14576), .I2(n14575), .O(n648) );
  AND_GATE U1094 ( .I1(n7290), .I2(n7289), .O(n649) );
  OR_GATE U1095 ( .I1(n14107), .I2(n14106), .O(n14109) );
  NAND_GATE U1096 ( .I1(n13637), .I2(n440), .O(n650) );
  AND_GATE U1097 ( .I1(n650), .I2(n438), .O(n14057) );
  NAND_GATE U1098 ( .I1(n651), .I2(n9321), .O(n9320) );
  NOR_GATE U1099 ( .I1(n9323), .I2(n9322), .O(n651) );
  NAND3_GATE U1100 ( .I1(n13964), .I2(n14058), .I3(n14061), .O(n652) );
  OR_GATE U1101 ( .I1(n5), .I2(n9713), .O(n9708) );
  NOR3_GATE U1102 ( .I1(n6472), .I2(n595), .I3(n6473), .O(n653) );
  NAND_GATE U1103 ( .I1(n654), .I2(n8842), .O(n8841) );
  NOR_GATE U1104 ( .I1(n8844), .I2(n8843), .O(n654) );
  NAND_GATE U1105 ( .I1(n655), .I2(n7965), .O(n7964) );
  NOR_GATE U1106 ( .I1(n7967), .I2(n7966), .O(n655) );
  NAND_GATE U1107 ( .I1(n6812), .I2(n658), .O(n656) );
  OR_GATE U1108 ( .I1(n6815), .I2(n6811), .O(n657) );
  AND_GATE U1109 ( .I1(n6813), .I2(n6823), .O(n658) );
  NAND_GATE U1110 ( .I1(n4881), .I2(n5314), .O(n659) );
  NAND_GATE U1111 ( .I1(n659), .I2(n660), .O(n5311) );
  AND_GATE U1112 ( .I1(n661), .I2(n4882), .O(n660) );
  INV_GATE U1113 ( .I1(n5320), .O(n661) );
  AND_GATE U1114 ( .I1(n9572), .I2(n9215), .O(n662) );
  AND_GATE U1115 ( .I1(n2024), .I2(n1879), .O(n663) );
  NAND_GATE U1116 ( .I1(n6786), .I2(n6501), .O(n664) );
  AND_GATE U1117 ( .I1(n14018), .I2(n14017), .O(n665) );
  NAND_GATE U1118 ( .I1(n1234), .I2(n667), .O(n11010) );
  AND_GATE U1119 ( .I1(n1235), .I2(n11009), .O(n667) );
  AND_GATE U1120 ( .I1(n11021), .I2(n11020), .O(n668) );
  NAND3_GATE U1121 ( .I1(n10624), .I2(n10400), .I3(n10610), .O(n669) );
  AND3_GATE U1122 ( .I1(n9806), .I2(n9805), .I3(n9804), .O(n670) );
  AND_GATE U1123 ( .I1(n9269), .I2(n9157), .O(n671) );
  AND3_GATE U1124 ( .I1(n9268), .I2(n9267), .I3(n9266), .O(n672) );
  AND3_GATE U1125 ( .I1(n8078), .I2(n8077), .I3(n8076), .O(n673) );
  AND3_GATE U1126 ( .I1(n6417), .I2(n6416), .I3(n6415), .O(n674) );
  AND3_GATE U1127 ( .I1(n4789), .I2(n4788), .I3(n5480), .O(n675) );
  AND_GATE U1128 ( .I1(n4546), .I2(n4545), .O(n676) );
  AND_GATE U1129 ( .I1(n11872), .I2(n11871), .O(n677) );
  AND3_GATE U1130 ( .I1(n10624), .I2(n10400), .I3(n10610), .O(n678) );
  AND_GATE U1131 ( .I1(n7394), .I2(n7393), .O(n679) );
  INV_GATE U1132 ( .I1(n679), .O(n7501) );
  AND_GATE U1133 ( .I1(n9661), .I2(n9660), .O(n680) );
  OR_GATE U1134 ( .I1(n8659), .I2(n791), .O(n8660) );
  AND3_GATE U1135 ( .I1(n5308), .I2(n5307), .I3(n4883), .O(n681) );
  INV_GATE U1136 ( .I1(n681), .O(n5298) );
  AND_GATE U1137 ( .I1(n682), .I2(n683), .O(n14084) );
  INV_GATE U1138 ( .I1(n14083), .O(n684) );
  OR_GATE U1139 ( .I1(n10849), .I2(n685), .O(n694) );
  NAND_GATE U1140 ( .I1(n10850), .I2(n10852), .O(n685) );
  AND3_GATE U1141 ( .I1(n11754), .I2(n12153), .I3(n12152), .O(n686) );
  INV_GATE U1142 ( .I1(n686), .O(n11952) );
  NAND_GATE U1143 ( .I1(n522), .I2(n689), .O(n687) );
  AND_GATE U1144 ( .I1(n687), .I2(n688), .O(n12424) );
  AND_GATE U1145 ( .I1(n12421), .I2(n12423), .O(n689) );
  NAND_GATE U1146 ( .I1(n9093), .I2(n692), .O(n690) );
  AND_GATE U1147 ( .I1(n690), .I2(n691), .O(n9099) );
  OR_GATE U1148 ( .I1(n9094), .I2(n9096), .O(n691) );
  AND_GATE U1149 ( .I1(n768), .I2(n9098), .O(n692) );
  NAND_GATE U1150 ( .I1(n10849), .I2(n696), .O(n693) );
  AND_GATE U1151 ( .I1(n693), .I2(n694), .O(n10853) );
  INV_GATE U1152 ( .I1(n10852), .O(n695) );
  NAND_GATE U1153 ( .I1(n13270), .I2(n699), .O(n697) );
  AND_GATE U1154 ( .I1(n697), .I2(n698), .O(n13274) );
  OR_GATE U1155 ( .I1(n13269), .I2(n13272), .O(n698) );
  AND_GATE U1156 ( .I1(n13271), .I2(n13273), .O(n699) );
  NAND_GATE U1157 ( .I1(n6257), .I2(n702), .O(n700) );
  AND_GATE U1158 ( .I1(n700), .I2(n701), .O(n6264) );
  OR_GATE U1159 ( .I1(n6259), .I2(n6252), .O(n701) );
  AND_GATE U1160 ( .I1(n6251), .I2(n5829), .O(n702) );
  NAND_GATE U1161 ( .I1(n5332), .I2(n705), .O(n703) );
  AND_GATE U1162 ( .I1(n703), .I2(n704), .O(n5338) );
  OR_GATE U1163 ( .I1(n5335), .I2(n5328), .O(n704) );
  AND_GATE U1164 ( .I1(n5327), .I2(n4871), .O(n705) );
  NOR_GATE U1165 ( .I1(n4603), .I2(n4602), .O(n706) );
  AND_GATE U1166 ( .I1(n7446), .I2(n7445), .O(n707) );
  AND3_GATE U1167 ( .I1(n6268), .I2(n6267), .I3(n6266), .O(n708) );
  AND3_GATE U1168 ( .I1(n5342), .I2(n5341), .I3(n5340), .O(n709) );
  AND_GATE U1169 ( .I1(n4646), .I2(n4645), .O(n710) );
  NAND3_GATE U1170 ( .I1(n7163), .I2(n7162), .I3(n7161), .O(n711) );
  AND3_GATE U1171 ( .I1(n3666), .I2(n3665), .I3(n3809), .O(n712) );
  AND_GATE U1172 ( .I1(n5733), .I2(n5737), .O(n713) );
  INV_GATE U1173 ( .I1(n713), .O(n6297) );
  OR_GATE U1174 ( .I1(n1361), .I2(n5736), .O(n5738) );
  OR_GATE U1175 ( .I1(n714), .I2(n5444), .O(n5446) );
  INV_GATE U1176 ( .I1(n5443), .O(n714) );
  NAND_GATE U1177 ( .I1(n9448), .I2(n717), .O(n715) );
  AND_GATE U1178 ( .I1(n715), .I2(n716), .O(n9451) );
  OR_GATE U1179 ( .I1(n9446), .I2(n9449), .O(n716) );
  AND_GATE U1180 ( .I1(n9447), .I2(n9450), .O(n717) );
  NAND_GATE U1181 ( .I1(n718), .I2(n6334), .O(n6330) );
  NOR_GATE U1182 ( .I1(n6338), .I2(n6333), .O(n718) );
  AND3_GATE U1183 ( .I1(n11551), .I2(n11280), .I3(n11550), .O(n719) );
  NAND_GATE U1184 ( .I1(n169), .I2(n722), .O(n720) );
  AND_GATE U1185 ( .I1(n720), .I2(n721), .O(n6320) );
  OR_GATE U1186 ( .I1(n6316), .I2(n6315), .O(n721) );
  AND_GATE U1187 ( .I1(n6323), .I2(n6319), .O(n722) );
  NAND_GATE U1188 ( .I1(n723), .I2(n14394), .O(n14393) );
  NAND_GATE U1189 ( .I1(n724), .I2(n11532), .O(n11531) );
  NOR_GATE U1190 ( .I1(n11534), .I2(n11533), .O(n724) );
  NAND_GATE U1191 ( .I1(n10679), .I2(n728), .O(n725) );
  AND_GATE U1192 ( .I1(n725), .I2(n726), .O(n11081) );
  OR_GATE U1193 ( .I1(n727), .I2(n10681), .O(n726) );
  INV_GATE U1194 ( .I1(n10682), .O(n727) );
  AND_GATE U1195 ( .I1(n10680), .I2(n10682), .O(n728) );
  OR_GATE U1196 ( .I1(n874), .I2(n732), .O(n729) );
  AND_GATE U1197 ( .I1(n729), .I2(n730), .O(n8554) );
  OR_GATE U1198 ( .I1(n731), .I2(n8551), .O(n730) );
  INV_GATE U1199 ( .I1(n8553), .O(n731) );
  OR_GATE U1200 ( .I1(n8550), .I2(n731), .O(n732) );
  AND3_GATE U1201 ( .I1(n7163), .I2(n7162), .I3(n7161), .O(n733) );
  AND3_GATE U1202 ( .I1(n13548), .I2(n13952), .I3(n13951), .O(n734) );
  OR3_GATE U1203 ( .I1(n735), .I2(n6399), .I3(n6398), .O(n6396) );
  INV_GATE U1204 ( .I1(n6391), .O(n735) );
  AND_GATE U1205 ( .I1(n12291), .I2(n289), .O(n12718) );
  AND_GATE U1206 ( .I1(n9747), .I2(n9746), .O(n736) );
  AND3_GATE U1207 ( .I1(n8931), .I2(n8930), .I3(n8614), .O(n737) );
  AND3_GATE U1208 ( .I1(n10561), .I2(n10560), .I3(n10559), .O(n738) );
  AND_GATE U1209 ( .I1(n12246), .I2(n12245), .O(n739) );
  AND_GATE U1210 ( .I1(n4630), .I2(n4629), .O(n740) );
  INV_GATE U1211 ( .I1(n740), .O(n4860) );
  AND3_GATE U1212 ( .I1(n9825), .I2(n9824), .I3(n9823), .O(n741) );
  AND_GATE U1213 ( .I1(n12337), .I2(n12222), .O(n742) );
  AND_GATE U1214 ( .I1(n10382), .I2(n10050), .O(n743) );
  AND_GATE U1215 ( .I1(n3592), .I2(n3593), .O(n744) );
  NAND_GATE U1216 ( .I1(n12751), .I2(n12752), .O(n745) );
  AND3_GATE U1217 ( .I1(n8452), .I2(n8451), .I3(n8450), .O(n746) );
  OR3_GATE U1218 ( .I1(n747), .I2(n748), .I3(n8886), .O(n8889) );
  INV_GATE U1219 ( .I1(n8884), .O(n747) );
  INV_GATE U1220 ( .I1(n8883), .O(n748) );
  OR_GATE U1221 ( .I1(n733), .I2(n7480), .O(n7476) );
  NAND_GATE U1222 ( .I1(n2904), .I2(n2903), .O(n749) );
  OR_GATE U1223 ( .I1(n11003), .I2(n154), .O(n11005) );
  OR_GATE U1224 ( .I1(n1256), .I2(n7685), .O(n7686) );
  OR3_GATE U1225 ( .I1(n576), .I2(n10158), .I3(n10154), .O(n10153) );
  OR3_GATE U1226 ( .I1(n750), .I2(n2979), .I3(n2970), .O(n2981) );
  INV_GATE U1227 ( .I1(n2976), .O(n750) );
  OR3_GATE U1228 ( .I1(n751), .I2(n2963), .I3(n2960), .O(n2958) );
  INV_GATE U1229 ( .I1(n2954), .O(n751) );
  OR_GATE U1230 ( .I1(n7574), .I2(n7573), .O(n7576) );
  OR_GATE U1231 ( .I1(n633), .I2(n9975), .O(n9977) );
  AND3_GATE U1232 ( .I1(n10843), .I2(n11250), .I3(n11249), .O(n752) );
  INV_GATE U1233 ( .I1(n752), .O(n11104) );
  NOR_GATE U1234 ( .I1(n6774), .I2(n6773), .O(n753) );
  INV_GATE U1235 ( .I1(n753), .O(n6768) );
  NAND_GATE U1236 ( .I1(n10457), .I2(n754), .O(n1209) );
  AND_GATE U1237 ( .I1(n10456), .I2(n10455), .O(n754) );
  AND3_GATE U1238 ( .I1(n9476), .I2(n9826), .I3(n9827), .O(n755) );
  INV_GATE U1239 ( .I1(n755), .O(n10038) );
  AND_GATE U1240 ( .I1(n5563), .I2(n5562), .O(n756) );
  INV_GATE U1241 ( .I1(n756), .O(n5832) );
  OR_GATE U1242 ( .I1(n4440), .I2(n757), .O(n4443) );
  INV_GATE U1243 ( .I1(n4439), .O(n757) );
  NAND_GATE U1244 ( .I1(n9160), .I2(n760), .O(n758) );
  AND_GATE U1245 ( .I1(n758), .I2(n759), .O(n9259) );
  OR_GATE U1246 ( .I1(n9158), .I2(n9163), .O(n759) );
  AND_GATE U1247 ( .I1(n9161), .I2(n9258), .O(n760) );
  NAND_GATE U1248 ( .I1(n4793), .I2(n763), .O(n761) );
  AND_GATE U1249 ( .I1(n761), .I2(n762), .O(n5389) );
  OR_GATE U1250 ( .I1(n4790), .I2(n4795), .O(n762) );
  AND_GATE U1251 ( .I1(n4792), .I2(n5399), .O(n763) );
  NAND_GATE U1252 ( .I1(n5772), .I2(n5771), .O(n764) );
  AND_GATE U1253 ( .I1(n11333), .I2(n11332), .O(n765) );
  AND3_GATE U1254 ( .I1(n7219), .I2(n7218), .I3(n7217), .O(n766) );
  AND3_GATE U1255 ( .I1(n3627), .I2(n3626), .I3(n3625), .O(n767) );
  INV_GATE U1256 ( .I1(n768), .O(n9095) );
  AND_GATE U1257 ( .I1(n9004), .I2(n9003), .O(n769) );
  INV_GATE U1258 ( .I1(n769), .O(n9427) );
  AND3_GATE U1259 ( .I1(n8404), .I2(n8248), .I3(n8403), .O(n770) );
  NAND_GATE U1260 ( .I1(n771), .I2(n7544), .O(n7543) );
  NOR_GATE U1261 ( .I1(n7546), .I2(n7545), .O(n771) );
  AND_GATE U1262 ( .I1(n8418), .I2(n8227), .O(n772) );
  INV_GATE U1263 ( .I1(n772), .O(n8402) );
  NAND_GATE U1264 ( .I1(n10487), .I2(n775), .O(n773) );
  AND_GATE U1265 ( .I1(n773), .I2(n774), .O(n10495) );
  OR_GATE U1266 ( .I1(n10491), .I2(n10488), .O(n774) );
  AND_GATE U1267 ( .I1(n10493), .I2(n15336), .O(n775) );
  NAND_GATE U1268 ( .I1(n776), .I2(n8820), .O(n8819) );
  NOR_GATE U1269 ( .I1(n8822), .I2(n8821), .O(n776) );
  NAND_GATE U1270 ( .I1(n777), .I2(n7943), .O(n7942) );
  NOR_GATE U1271 ( .I1(n7945), .I2(n7944), .O(n777) );
  AND_GATE U1272 ( .I1(n6220), .I2(n6219), .O(n778) );
  OR_GATE U1273 ( .I1(n801), .I2(n793), .O(n779) );
  AND3_GATE U1274 ( .I1(n3573), .I2(n3572), .I3(n3571), .O(n780) );
  NAND_GATE U1275 ( .I1(n2996), .I2(n2812), .O(n781) );
  NOR_GATE U1276 ( .I1(n13135), .I2(n12758), .O(n920) );
  AND_GATE U1277 ( .I1(n10421), .I2(n10095), .O(n782) );
  OR3_GATE U1278 ( .I1(n783), .I2(n5507), .I3(n5505), .O(n5509) );
  INV_GATE U1279 ( .I1(n5502), .O(n783) );
  NOR_GATE U1280 ( .I1(n5788), .I2(n5787), .O(n784) );
  AND_GATE U1281 ( .I1(n6422), .I2(n6421), .O(n785) );
  INV_GATE U1282 ( .I1(n785), .O(n6553) );
  OR_GATE U1283 ( .I1(n1290), .I2(n786), .O(n6716) );
  AND_GATE U1284 ( .I1(n7187), .I2(n7190), .O(n786) );
  AND_GATE U1285 ( .I1(n14823), .I2(n15054), .O(n787) );
  INV_GATE U1286 ( .I1(n787), .O(n15033) );
  AND3_GATE U1287 ( .I1(n5296), .I2(n5568), .I3(n5567), .O(n788) );
  INV_GATE U1288 ( .I1(n788), .O(n5853) );
  AND_GATE U1289 ( .I1(n6816), .I2(n6515), .O(n789) );
  AND_GATE U1290 ( .I1(n6496), .I2(n6495), .O(n790) );
  INV_GATE U1291 ( .I1(n790), .O(n6771) );
  AND_GATE U1292 ( .I1(n8321), .I2(n8320), .O(n791) );
  AND_GATE U1293 ( .I1(n10926), .I2(n10925), .O(n792) );
  OR_GATE U1294 ( .I1(n824), .I2(n6801), .O(n6802) );
  NOR_GATE U1295 ( .I1(n801), .I2(n793), .O(n872) );
  AND_GATE U1296 ( .I1(n5832), .I2(n5564), .O(n793) );
  AND_GATE U1297 ( .I1(n5750), .I2(n5749), .O(n794) );
  AND_GATE U1298 ( .I1(n795), .I2(n796), .O(n1972) );
  OR_GATE U1299 ( .I1(n797), .I2(n1880), .O(n796) );
  INV_GATE U1300 ( .I1(n1981), .O(n797) );
  AND_GATE U1301 ( .I1(n5899), .I2(n5581), .O(n798) );
  AND_GATE U1302 ( .I1(n3542), .I2(n3541), .O(n799) );
  AND3_GATE U1303 ( .I1(n2110), .I2(n2109), .I3(n2111), .O(n800) );
  NOR_GATE U1304 ( .I1(n5834), .I2(n5831), .O(n801) );
  NAND3_GATE U1305 ( .I1(n3899), .I2(n3898), .I3(n3900), .O(n802) );
  OR_GATE U1306 ( .I1(n9538), .I2(n176), .O(n9540) );
  OR_GATE U1307 ( .I1(n3809), .I2(n3817), .O(n4582) );
  AND_GATE U1308 ( .I1(n805), .I2(n1310), .O(n803) );
  AND_GATE U1309 ( .I1(n1980), .I2(n1979), .O(n804) );
  INV_GATE U1310 ( .I1(n804), .O(n2720) );
  AND3_GATE U1311 ( .I1(n3054), .I2(n3051), .I3(n3548), .O(n805) );
  OR_GATE U1312 ( .I1(n799), .I2(n3981), .O(n3979) );
  AND3_GATE U1313 ( .I1(n9777), .I2(n9776), .I3(n9775), .O(n806) );
  AND_GATE U1314 ( .I1(n8299), .I2(n8298), .O(n807) );
  OR_GATE U1315 ( .I1(n1053), .I2(n810), .O(n808) );
  OR_GATE U1316 ( .I1(n1415), .I2(n8291), .O(n809) );
  OR_GATE U1317 ( .I1(n1360), .I2(n1415), .O(n810) );
  AND_GATE U1318 ( .I1(n5531), .I2(n5530), .O(n811) );
  OR_GATE U1319 ( .I1(n5646), .I2(n819), .O(n812) );
  AND3_GATE U1320 ( .I1(n4577), .I2(n4576), .I3(n4575), .O(n813) );
  AND3_GATE U1321 ( .I1(n3652), .I2(n3651), .I3(n3650), .O(n814) );
  AND3_GATE U1322 ( .I1(n8606), .I2(n8605), .I3(n9191), .O(n815) );
  AND3_GATE U1323 ( .I1(n6550), .I2(n6549), .I3(n6548), .O(n816) );
  AND_GATE U1324 ( .I1(n6431), .I2(n6430), .O(n817) );
  INV_GATE U1325 ( .I1(n818), .O(n1310) );
  NOR_GATE U1326 ( .I1(n5646), .I2(n819), .O(n1241) );
  INV_GATE U1327 ( .I1(n6458), .O(n819) );
  NOR_GATE U1328 ( .I1(n3863), .I2(n3862), .O(n820) );
  AND_GATE U1329 ( .I1(n10471), .I2(n10110), .O(n821) );
  INV_GATE U1330 ( .I1(n821), .O(n10493) );
  OR_GATE U1331 ( .I1(n1309), .I2(n3049), .O(n3042) );
  AND3_GATE U1332 ( .I1(n8941), .I2(n8595), .I3(n8940), .O(n822) );
  INV_GATE U1333 ( .I1(n822), .O(n9171) );
  AND_GATE U1334 ( .I1(n5772), .I2(n5771), .O(n823) );
  OR_GATE U1335 ( .I1(n10477), .I2(n1242), .O(n10478) );
  AND_GATE U1336 ( .I1(n6786), .I2(n6501), .O(n824) );
  OR_GATE U1337 ( .I1(n788), .I2(n5857), .O(n5851) );
  AND3_GATE U1338 ( .I1(n10129), .I2(n10082), .I3(n10128), .O(n825) );
  INV_GATE U1339 ( .I1(n825), .O(n10124) );
  AND_GATE U1340 ( .I1(n11000), .I2(n11004), .O(n826) );
  AND_GATE U1341 ( .I1(n6491), .I2(n6490), .O(n827) );
  INV_GATE U1342 ( .I1(n827), .O(n7423) );
  AND_GATE U1343 ( .I1(n14829), .I2(n15015), .O(n828) );
  INV_GATE U1344 ( .I1(n828), .O(n14994) );
  NAND_GATE U1345 ( .I1(n829), .I2(n5283), .O(n5282) );
  NOR_GATE U1346 ( .I1(n5285), .I2(n5284), .O(n829) );
  AND_GATE U1347 ( .I1(n8837), .I2(n8836), .O(n830) );
  AND_GATE U1348 ( .I1(n7960), .I2(n7959), .O(n831) );
  AND_GATE U1349 ( .I1(n7098), .I2(n7097), .O(n832) );
  NAND_GATE U1350 ( .I1(n8694), .I2(n835), .O(n833) );
  AND_GATE U1351 ( .I1(n833), .I2(n834), .O(n8827) );
  OR_GATE U1352 ( .I1(n8833), .I2(n8697), .O(n834) );
  AND_GATE U1353 ( .I1(n8695), .I2(n8698), .O(n835) );
  NAND_GATE U1354 ( .I1(n7766), .I2(n838), .O(n836) );
  AND_GATE U1355 ( .I1(n836), .I2(n837), .O(n7950) );
  OR_GATE U1356 ( .I1(n7956), .I2(n7769), .O(n837) );
  AND_GATE U1357 ( .I1(n7767), .I2(n7770), .O(n838) );
  AND_GATE U1358 ( .I1(n2972), .I2(n2808), .O(n839) );
  INV_GATE U1359 ( .I1(n839), .O(n2991) );
  OR_GATE U1360 ( .I1(n7503), .I2(n679), .O(n7498) );
  NAND_GATE U1361 ( .I1(n14855), .I2(n842), .O(n840) );
  OR_GATE U1362 ( .I1(n14854), .I2(n14857), .O(n841) );
  AND_GATE U1363 ( .I1(n1319), .I2(n14858), .O(n842) );
  NAND_GATE U1364 ( .I1(n843), .I2(n10008), .O(n10007) );
  NOR_GATE U1365 ( .I1(n10010), .I2(n10009), .O(n843) );
  AND3_GATE U1366 ( .I1(n9312), .I2(n9108), .I3(n9307), .O(n844) );
  INV_GATE U1367 ( .I1(n844), .O(n9303) );
  NAND_GATE U1368 ( .I1(n9576), .I2(n847), .O(n845) );
  OR_GATE U1369 ( .I1(n9574), .I2(n9579), .O(n846) );
  AND_GATE U1370 ( .I1(n9575), .I2(n9580), .O(n847) );
  NAND_GATE U1371 ( .I1(n4905), .I2(n850), .O(n848) );
  AND_GATE U1372 ( .I1(n848), .I2(n849), .O(n4910) );
  OR_GATE U1373 ( .I1(n4903), .I2(n4908), .O(n849) );
  AND_GATE U1374 ( .I1(n4904), .I2(n4909), .O(n850) );
  NAND_GATE U1375 ( .I1(n788), .I2(n853), .O(n851) );
  AND_GATE U1376 ( .I1(n851), .I2(n852), .O(n5865) );
  OR_GATE U1377 ( .I1(n5855), .I2(n5851), .O(n852) );
  AND_GATE U1378 ( .I1(n5857), .I2(n5864), .O(n853) );
  NOR_GATE U1379 ( .I1(n4503), .I2(n4549), .O(n854) );
  INV_GATE U1380 ( .I1(n854), .O(n4793) );
  OR3_GATE U1381 ( .I1(n855), .I2(n6429), .I3(n5792), .O(n6432) );
  INV_GATE U1382 ( .I1(n5793), .O(n855) );
  AND3_GATE U1383 ( .I1(n4628), .I2(n4627), .I3(n4626), .O(n856) );
  AND3_GATE U1384 ( .I1(n10198), .I2(n10016), .I3(n10191), .O(n857) );
  INV_GATE U1385 ( .I1(n857), .O(n10187) );
  OR_GATE U1386 ( .I1(n10194), .I2(n10199), .O(n10197) );
  AND_GATE U1387 ( .I1(n7134), .I2(n7133), .O(n858) );
  OR_GATE U1388 ( .I1(n8184), .I2(n859), .O(n8188) );
  INV_GATE U1389 ( .I1(n8186), .O(n859) );
  AND3_GATE U1390 ( .I1(n10204), .I2(n10003), .I3(n10203), .O(n860) );
  INV_GATE U1391 ( .I1(n860), .O(n10356) );
  AND_GATE U1392 ( .I1(n2904), .I2(n2903), .O(n861) );
  AND3_GATE U1393 ( .I1(n13964), .I2(n14058), .I3(n14061), .O(n862) );
  NAND_GATE U1394 ( .I1(n863), .I2(n6210), .O(n6218) );
  INV_GATE U1395 ( .I1(n6215), .O(n863) );
  AND_GATE U1396 ( .I1(n864), .I2(n865), .O(n11580) );
  NAND_GATE U1397 ( .I1(n866), .I2(n13912), .O(n13911) );
  NOR_GATE U1398 ( .I1(n13913), .I2(n13914), .O(n866) );
  NAND_GATE U1399 ( .I1(n867), .I2(n9332), .O(n9331) );
  NOR_GATE U1400 ( .I1(n9334), .I2(n9333), .O(n867) );
  NAND_GATE U1401 ( .I1(n14832), .I2(n870), .O(n868) );
  AND_GATE U1402 ( .I1(n868), .I2(n869), .O(n14975) );
  AND_GATE U1403 ( .I1(n14981), .I2(n14968), .O(n870) );
  OR3_GATE U1404 ( .I1(n871), .I2(n3006), .I3(n2997), .O(n3003) );
  INV_GATE U1405 ( .I1(n2999), .O(n871) );
  AND_GATE U1406 ( .I1(n2996), .I2(n2812), .O(n873) );
  OR_GATE U1407 ( .I1(n875), .I2(n5291), .O(n5571) );
  INV_GATE U1408 ( .I1(n5290), .O(n875) );
  AND_GATE U1409 ( .I1(n877), .I2(n9231), .O(n876) );
  INV_GATE U1410 ( .I1(n9764), .O(n877) );
  OR_GATE U1411 ( .I1(n874), .I2(n8550), .O(n8552) );
  OR_GATE U1412 ( .I1(n10594), .I2(n878), .O(n10583) );
  INV_GATE U1413 ( .I1(n10598), .O(n878) );
  OR_GATE U1414 ( .I1(n9271), .I2(n9270), .O(n9273) );
  OR_GATE U1415 ( .I1(n8909), .I2(n8905), .O(n9201) );
  OR_GATE U1416 ( .I1(n10382), .I2(n10379), .O(n10640) );
  OR_GATE U1417 ( .I1(n10051), .I2(n10054), .O(n10140) );
  OR_GATE U1418 ( .I1(n8306), .I2(n8307), .O(n8309) );
  OR_GATE U1419 ( .I1(n10391), .I2(n879), .O(n10613) );
  INV_GATE U1420 ( .I1(n10395), .O(n879) );
  OR_GATE U1421 ( .I1(n11308), .I2(n11306), .O(n11507) );
  OR_GATE U1422 ( .I1(n8395), .I2(n770), .O(n8588) );
  OR_GATE U1423 ( .I1(n9302), .I2(n844), .O(n9462) );
  OR_GATE U1424 ( .I1(n8023), .I2(n880), .O(n8027) );
  INV_GATE U1425 ( .I1(n8024), .O(n880) );
  INV_GATE U1426 ( .I1(n14062), .O(n881) );
  OR_GATE U1427 ( .I1(n12297), .I2(n882), .O(n12227) );
  INV_GATE U1428 ( .I1(n12300), .O(n882) );
  OR_GATE U1429 ( .I1(n11460), .I2(n883), .O(n11451) );
  INV_GATE U1430 ( .I1(n11455), .O(n883) );
  OR_GATE U1431 ( .I1(n9482), .I2(n9483), .O(n9490) );
  OR_GATE U1432 ( .I1(n884), .I2(n8842), .O(n8845) );
  INV_GATE U1433 ( .I1(n8843), .O(n884) );
  OR_GATE U1434 ( .I1(n885), .I2(n7965), .O(n7968) );
  INV_GATE U1435 ( .I1(n7966), .O(n885) );
  OR_GATE U1436 ( .I1(n886), .I2(n7954), .O(n7957) );
  INV_GATE U1437 ( .I1(n7955), .O(n886) );
  OR_GATE U1438 ( .I1(n9), .I2(n8831), .O(n8834) );
  OR_GATE U1439 ( .I1(n887), .I2(n7943), .O(n7946) );
  INV_GATE U1440 ( .I1(n7944), .O(n887) );
  OR_GATE U1441 ( .I1(n9740), .I2(n9741), .O(n9743) );
  OR_GATE U1442 ( .I1(n888), .I2(n8820), .O(n8823) );
  INV_GATE U1443 ( .I1(n8821), .O(n888) );
  OR_GATE U1444 ( .I1(n889), .I2(n9679), .O(n9674) );
  INV_GATE U1445 ( .I1(n9676), .O(n889) );
  OR_GATE U1446 ( .I1(n890), .I2(n9666), .O(n9669) );
  INV_GATE U1447 ( .I1(n9667), .O(n890) );
  OR_GATE U1448 ( .I1(n184), .I2(n7173), .O(n7175) );
  OR_GATE U1449 ( .I1(n891), .I2(n14852), .O(n14861) );
  INV_GATE U1450 ( .I1(n14856), .O(n891) );
  OR_GATE U1451 ( .I1(n11857), .I2(n892), .O(n12300) );
  INV_GATE U1452 ( .I1(n12296), .O(n892) );
  OR_GATE U1453 ( .I1(n7240), .I2(n1359), .O(n7242) );
  OR_GATE U1454 ( .I1(n11548), .I2(n893), .O(n11940) );
  INV_GATE U1455 ( .I1(n11549), .O(n893) );
  OR_GATE U1456 ( .I1(n13627), .I2(n13626), .O(n13972) );
  OR_GATE U1457 ( .I1(n10681), .I2(n727), .O(n11084) );
  OR_GATE U1458 ( .I1(n12759), .I2(n13133), .O(n13138) );
  OR_GATE U1459 ( .I1(n9724), .I2(n9725), .O(n9734) );
  OR_GATE U1460 ( .I1(n8953), .I2(n8951), .O(n8958) );
  OR_GATE U1461 ( .I1(n894), .I2(n11385), .O(n11387) );
  INV_GATE U1462 ( .I1(n11393), .O(n894) );
  OR_GATE U1463 ( .I1(n12358), .I2(n895), .O(n12782) );
  INV_GATE U1464 ( .I1(n12361), .O(n895) );
  OR_GATE U1465 ( .I1(n10912), .I2(n678), .O(n11011) );
  OR_GATE U1466 ( .I1(n896), .I2(n7992), .O(n7995) );
  INV_GATE U1467 ( .I1(n7993), .O(n896) );
  OR_GATE U1468 ( .I1(n11539), .I2(n719), .O(n11549) );
  OR_GATE U1469 ( .I1(n336), .I2(n13106), .O(n13108) );
  OR_GATE U1470 ( .I1(n568), .I2(n14022), .O(n14026) );
  OR_GATE U1471 ( .I1(n897), .I2(n10933), .O(n10940) );
  INV_GATE U1472 ( .I1(n10934), .O(n897) );
  OR_GATE U1473 ( .I1(n514), .I2(n13592), .O(n13596) );
  OR_GATE U1474 ( .I1(n13608), .I2(n230), .O(n13602) );
  OR_GATE U1475 ( .I1(n12337), .I2(n1232), .O(n12756) );
  OR_GATE U1476 ( .I1(n13631), .I2(n734), .O(n13640) );
  OR_GATE U1477 ( .I1(n10071), .I2(n898), .O(n10075) );
  INV_GATE U1478 ( .I1(n10072), .O(n898) );
  OR_GATE U1479 ( .I1(n899), .I2(n9831), .O(n9837) );
  INV_GATE U1480 ( .I1(n9832), .O(n899) );
  OR_GATE U1481 ( .I1(n10654), .I2(n279), .O(n10647) );
  OR_GATE U1482 ( .I1(n11062), .I2(n900), .O(n10871) );
  INV_GATE U1483 ( .I1(n11071), .O(n900) );
  OR_GATE U1484 ( .I1(n901), .I2(n8879), .O(n8884) );
  INV_GATE U1485 ( .I1(n8880), .O(n901) );
  OR_GATE U1486 ( .I1(n80), .I2(n8809), .O(n8812) );
  OR_GATE U1487 ( .I1(n902), .I2(n9655), .O(n9658) );
  INV_GATE U1488 ( .I1(n9656), .O(n902) );
  OR_GATE U1489 ( .I1(n11055), .I2(n11047), .O(n11057) );
  OR_GATE U1490 ( .I1(n8418), .I2(n8410), .O(n8420) );
  OR_GATE U1491 ( .I1(n11101), .I2(n752), .O(n11111) );
  OR_GATE U1492 ( .I1(n903), .I2(n14539), .O(n14551) );
  INV_GATE U1493 ( .I1(n14543), .O(n903) );
  OR_GATE U1494 ( .I1(n9467), .I2(n9470), .O(n9832) );
  OR_GATE U1495 ( .I1(n904), .I2(n7933), .O(n7936) );
  INV_GATE U1496 ( .I1(n7934), .O(n904) );
  OR_GATE U1497 ( .I1(n905), .I2(n7923), .O(n7926) );
  INV_GATE U1498 ( .I1(n7924), .O(n905) );
  OR_GATE U1499 ( .I1(n95), .I2(n8798), .O(n8801) );
  OR_GATE U1500 ( .I1(n906), .I2(n12830), .O(n12842) );
  INV_GATE U1501 ( .I1(n12834), .O(n906) );
  OR_GATE U1502 ( .I1(n907), .I2(n11960), .O(n11970) );
  INV_GATE U1503 ( .I1(n11964), .O(n907) );
  OR_GATE U1504 ( .I1(n13088), .I2(n908), .O(n13099) );
  INV_GATE U1505 ( .I1(n13092), .O(n908) );
  OR_GATE U1506 ( .I1(n909), .I2(n13669), .O(n13679) );
  INV_GATE U1507 ( .I1(n13672), .O(n909) );
  OR_GATE U1508 ( .I1(n12186), .I2(n910), .O(n12198) );
  INV_GATE U1509 ( .I1(n12190), .O(n910) );
  OR_GATE U1510 ( .I1(n911), .I2(n7912), .O(n7915) );
  INV_GATE U1511 ( .I1(n7913), .O(n911) );
  OR_GATE U1512 ( .I1(n912), .I2(n8787), .O(n8790) );
  INV_GATE U1513 ( .I1(n8788), .O(n912) );
  OR_GATE U1514 ( .I1(n913), .I2(n7901), .O(n7904) );
  INV_GATE U1515 ( .I1(n7902), .O(n913) );
  OR_GATE U1516 ( .I1(n914), .I2(n7890), .O(n7893) );
  INV_GATE U1517 ( .I1(n7891), .O(n914) );
  OR_GATE U1518 ( .I1(n9228), .I2(n14), .O(n9755) );
  OR_GATE U1519 ( .I1(n8616), .I2(n590), .O(n8917) );
  OR_GATE U1520 ( .I1(n6950), .I2(n6944), .O(n7003) );
  OR_GATE U1521 ( .I1(n7030), .I2(n282), .O(n7856) );
  AND_GATE U1522 ( .I1(n11838), .I2(n11837), .O(n915) );
  OR_GATE U1523 ( .I1(n9269), .I2(n9270), .O(n9822) );
  OR_GATE U1524 ( .I1(n10180), .I2(n10181), .O(n10186) );
  AND_GATE U1525 ( .I1(n9504), .I2(n9780), .O(n916) );
  OR_GATE U1526 ( .I1(n7605), .I2(n917), .O(n8104) );
  AND_GATE U1527 ( .I1(n12302), .I2(n12227), .O(n918) );
  AND_GATE U1528 ( .I1(n8629), .I2(n8893), .O(n919) );
  OR_GATE U1529 ( .I1(n9299), .I2(n9459), .O(n9302) );
  OR_GATE U1530 ( .I1(n6753), .I2(n827), .O(n7422) );
  OR_GATE U1531 ( .I1(n9232), .I2(n921), .O(n9230) );
  INV_GATE U1532 ( .I1(n9233), .O(n921) );
  OR_GATE U1533 ( .I1(n12354), .I2(n525), .O(n12349) );
  OR_GATE U1534 ( .I1(n922), .I2(n11909), .O(n11903) );
  INV_GATE U1535 ( .I1(n11906), .O(n922) );
  OR_GATE U1536 ( .I1(n13955), .I2(n365), .O(n13958) );
  OR_GATE U1537 ( .I1(n13539), .I2(n923), .O(n13542) );
  INV_GATE U1538 ( .I1(n13540), .O(n923) );
  OR_GATE U1539 ( .I1(n188), .I2(n11494), .O(n11496) );
  OR_GATE U1540 ( .I1(n116), .I2(n12800), .O(n12803) );
  OR_GATE U1541 ( .I1(n13076), .I2(n360), .O(n13079) );
  OR_GATE U1542 ( .I1(n924), .I2(n12397), .O(n12400) );
  INV_GATE U1543 ( .I1(n12398), .O(n924) );
  OR_GATE U1544 ( .I1(n13941), .I2(n361), .O(n13944) );
  OR_GATE U1545 ( .I1(n14394), .I2(n418), .O(n14397) );
  OR_GATE U1546 ( .I1(n925), .I2(n7103), .O(n7106) );
  INV_GATE U1547 ( .I1(n7104), .O(n925) );
  OR_GATE U1548 ( .I1(n926), .I2(n7092), .O(n7095) );
  INV_GATE U1549 ( .I1(n7093), .O(n926) );
  OR_GATE U1550 ( .I1(n13525), .I2(n927), .O(n13528) );
  INV_GATE U1551 ( .I1(n13526), .O(n927) );
  OR_GATE U1552 ( .I1(n928), .I2(n11532), .O(n11535) );
  INV_GATE U1553 ( .I1(n11533), .O(n928) );
  OR_GATE U1554 ( .I1(n12648), .I2(n929), .O(n12651) );
  INV_GATE U1555 ( .I1(n12649), .O(n929) );
  OR_GATE U1556 ( .I1(n13912), .I2(n930), .O(n13915) );
  INV_GATE U1557 ( .I1(n13913), .O(n930) );
  OR_GATE U1558 ( .I1(n8939), .I2(n931), .O(n8937) );
  INV_GATE U1559 ( .I1(n8942), .O(n931) );
  OR_GATE U1560 ( .I1(n13047), .I2(n932), .O(n13050) );
  INV_GATE U1561 ( .I1(n13048), .O(n932) );
  OR_GATE U1562 ( .I1(n933), .I2(n11554), .O(n11557) );
  INV_GATE U1563 ( .I1(n11555), .O(n933) );
  OR_GATE U1564 ( .I1(n14556), .I2(n934), .O(n14559) );
  INV_GATE U1565 ( .I1(n14557), .O(n934) );
  OR_GATE U1566 ( .I1(n10664), .I2(n170), .O(n10662) );
  OR_GATE U1567 ( .I1(n12141), .I2(n935), .O(n12144) );
  INV_GATE U1568 ( .I1(n12142), .O(n935) );
  OR_GATE U1569 ( .I1(n936), .I2(n9803), .O(n9798) );
  INV_GATE U1570 ( .I1(n9796), .O(n936) );
  OR_GATE U1571 ( .I1(n7672), .I2(n937), .O(n7674) );
  INV_GATE U1572 ( .I1(n7671), .O(n937) );
  OR_GATE U1573 ( .I1(n7403), .I2(n7402), .O(n7405) );
  OR_GATE U1574 ( .I1(n508), .I2(n10687), .O(n10690) );
  OR_GATE U1575 ( .I1(n8349), .I2(n8350), .O(n8352) );
  OR_GATE U1576 ( .I1(n11253), .I2(n938), .O(n11256) );
  INV_GATE U1577 ( .I1(n11254), .O(n938) );
  OR_GATE U1578 ( .I1(n14497), .I2(n435), .O(n14493) );
  OR_GATE U1579 ( .I1(n173), .I2(n8096), .O(n8098) );
  OR_GATE U1580 ( .I1(n939), .I2(n7536), .O(n7530) );
  INV_GATE U1581 ( .I1(n7533), .O(n939) );
  OR_GATE U1582 ( .I1(n9308), .I2(n940), .O(n9310) );
  INV_GATE U1583 ( .I1(n9313), .O(n940) );
  OR_GATE U1584 ( .I1(n941), .I2(n9844), .O(n9845) );
  INV_GATE U1585 ( .I1(n9849), .O(n941) );
  OR_GATE U1586 ( .I1(n7620), .I2(n189), .O(n7622) );
  OR_GATE U1587 ( .I1(n942), .I2(n8988), .O(n8991) );
  INV_GATE U1588 ( .I1(n8989), .O(n942) );
  OR_GATE U1589 ( .I1(n943), .I2(n10008), .O(n10011) );
  INV_GATE U1590 ( .I1(n10009), .O(n943) );
  OR_GATE U1591 ( .I1(n944), .I2(n9332), .O(n9335) );
  INV_GATE U1592 ( .I1(n9333), .O(n944) );
  OR_GATE U1593 ( .I1(n945), .I2(n10341), .O(n10344) );
  INV_GATE U1594 ( .I1(n10342), .O(n945) );
  OR_GATE U1595 ( .I1(n9261), .I2(n9262), .O(n9263) );
  NOR_GATE U1596 ( .I1(n946), .I2(n1291), .O(n12751) );
  AND_GATE U1597 ( .I1(n12336), .I2(n742), .O(n946) );
  NOR_GATE U1598 ( .I1(n11849), .I2(n479), .O(\A2[38] ) );
  AND_GATE U1599 ( .I1(n11503), .I2(n11505), .O(n947) );
  OR_GATE U1600 ( .I1(n452), .I2(n13197), .O(n13559) );
  OR_GATE U1601 ( .I1(n7658), .I2(n7659), .O(n8233) );
  OR_GATE U1602 ( .I1(n10465), .I2(n948), .O(n10467) );
  INV_GATE U1603 ( .I1(n10463), .O(n948) );
  OR_GATE U1604 ( .I1(n9093), .I2(n9098), .O(n9091) );
  AND_GATE U1605 ( .I1(n9750), .I2(n9752), .O(n949) );
  OR_GATE U1606 ( .I1(n6833), .I2(n789), .O(n6842) );
  OR_GATE U1607 ( .I1(n6816), .I2(n6812), .O(n6826) );
  AND_GATE U1608 ( .I1(n9164), .I2(n9260), .O(n950) );
  AND_GATE U1609 ( .I1(n6463), .I2(n6462), .O(n951) );
  OR_GATE U1610 ( .I1(n8946), .I2(n8947), .O(n8959) );
  AND_GATE U1611 ( .I1(n7687), .I2(n8262), .O(n952) );
  OR_GATE U1612 ( .I1(n953), .I2(n7146), .O(n7150) );
  INV_GATE U1613 ( .I1(n7147), .O(n953) );
  OR_GATE U1614 ( .I1(n14543), .I2(n14542), .O(n14545) );
  OR_GATE U1615 ( .I1(n13228), .I2(n13227), .O(n13229) );
  OR_GATE U1616 ( .I1(n12372), .I2(n12373), .O(n12376) );
  OR_GATE U1617 ( .I1(n954), .I2(n11015), .O(n11017) );
  INV_GATE U1618 ( .I1(n11016), .O(n954) );
  OR_GATE U1619 ( .I1(n232), .I2(n11917), .O(n11919) );
  OR_GATE U1620 ( .I1(n955), .I2(n10132), .O(n10134) );
  INV_GATE U1621 ( .I1(n10133), .O(n955) );
  OR_GATE U1622 ( .I1(n956), .I2(n11927), .O(n11930) );
  INV_GATE U1623 ( .I1(n11928), .O(n956) );
  OR_GATE U1624 ( .I1(n13927), .I2(n49), .O(n13930) );
  OR_GATE U1625 ( .I1(n957), .I2(n11514), .O(n11509) );
  INV_GATE U1626 ( .I1(n11511), .O(n957) );
  OR_GATE U1627 ( .I1(n14379), .I2(n556), .O(n14382) );
  OR_GATE U1628 ( .I1(n242), .I2(n10605), .O(n10600) );
  OR_GATE U1629 ( .I1(n958), .I2(n7081), .O(n7084) );
  INV_GATE U1630 ( .I1(n7082), .O(n958) );
  OR_GATE U1631 ( .I1(n959), .I2(n7114), .O(n7117) );
  INV_GATE U1632 ( .I1(n7115), .O(n959) );
  OR_GATE U1633 ( .I1(n13061), .I2(n960), .O(n13064) );
  INV_GATE U1634 ( .I1(n13062), .O(n960) );
  OR_GATE U1635 ( .I1(n13619), .I2(n401), .O(n13617) );
  OR_GATE U1636 ( .I1(n12156), .I2(n961), .O(n12159) );
  INV_GATE U1637 ( .I1(n12157), .O(n961) );
  OR_GATE U1638 ( .I1(n14349), .I2(n962), .O(n14352) );
  INV_GATE U1639 ( .I1(n14350), .O(n962) );
  OR_GATE U1640 ( .I1(n13494), .I2(n963), .O(n13497) );
  INV_GATE U1641 ( .I1(n13495), .O(n963) );
  OR_GATE U1642 ( .I1(n14046), .I2(n599), .O(n14045) );
  OR_GATE U1643 ( .I1(n12617), .I2(n964), .O(n12620) );
  INV_GATE U1644 ( .I1(n12618), .O(n964) );
  OR_GATE U1645 ( .I1(n965), .I2(n11095), .O(n11098) );
  INV_GATE U1646 ( .I1(n11096), .O(n965) );
  OR_GATE U1647 ( .I1(n14532), .I2(n966), .O(n14535) );
  INV_GATE U1648 ( .I1(n14533), .O(n966) );
  OR_GATE U1649 ( .I1(n10040), .I2(n755), .O(n10042) );
  OR_GATE U1650 ( .I1(n967), .I2(n9281), .O(n9275) );
  INV_GATE U1651 ( .I1(n9278), .O(n967) );
  OR_GATE U1652 ( .I1(n592), .I2(n14449), .O(n14452) );
  OR_GATE U1653 ( .I1(n11728), .I2(n968), .O(n11731) );
  INV_GATE U1654 ( .I1(n11729), .O(n968) );
  OR_GATE U1655 ( .I1(n969), .I2(n10207), .O(n10210) );
  INV_GATE U1656 ( .I1(n10208), .O(n969) );
  OR_GATE U1657 ( .I1(n970), .I2(n8457), .O(n8460) );
  INV_GATE U1658 ( .I1(n8458), .O(n970) );
  OR_GATE U1659 ( .I1(n971), .I2(n9321), .O(n9324) );
  INV_GATE U1660 ( .I1(n9322), .O(n971) );
  OR_GATE U1661 ( .I1(n14012), .I2(n972), .O(n14014) );
  INV_GATE U1662 ( .I1(n14016), .O(n972) );
  OR_GATE U1663 ( .I1(n14457), .I2(n601), .O(n14459) );
  OR_GATE U1664 ( .I1(n10982), .I2(n973), .O(n10985) );
  INV_GATE U1665 ( .I1(n10984), .O(n973) );
  OR_GATE U1666 ( .I1(n493), .I2(n11381), .O(n11375) );
  OR_GATE U1667 ( .I1(n14869), .I2(n441), .O(n14865) );
  OR_GATE U1668 ( .I1(n974), .I2(n9878), .O(n9881) );
  INV_GATE U1669 ( .I1(n9879), .O(n974) );
  OR_GATE U1670 ( .I1(n10722), .I2(n975), .O(n10725) );
  INV_GATE U1671 ( .I1(n10723), .O(n975) );
  OR_GATE U1672 ( .I1(n6592), .I2(n976), .O(n6586) );
  INV_GATE U1673 ( .I1(n6595), .O(n976) );
  OR_GATE U1674 ( .I1(n9560), .I2(n513), .O(n9701) );
  OR_GATE U1675 ( .I1(n680), .I2(n10113), .O(n10114) );
  OR_GATE U1676 ( .I1(n8369), .I2(n977), .O(n8367) );
  INV_GATE U1677 ( .I1(n8373), .O(n977) );
  AND_GATE U1678 ( .I1(n13140), .I2(n13175), .O(n978) );
  OR_GATE U1679 ( .I1(n6881), .I2(n979), .O(n6891) );
  INV_GATE U1680 ( .I1(n6882), .O(n979) );
  OR_GATE U1681 ( .I1(n6898), .I2(n980), .O(n6908) );
  INV_GATE U1682 ( .I1(n6899), .O(n980) );
  OR_GATE U1683 ( .I1(n6850), .I2(n6847), .O(n6858) );
  OR_GATE U1684 ( .I1(n6915), .I2(n981), .O(n6925) );
  INV_GATE U1685 ( .I1(n6916), .O(n981) );
  OR_GATE U1686 ( .I1(n769), .I2(n9429), .O(n9431) );
  OR_GATE U1687 ( .I1(n6973), .I2(n6972), .O(n6975) );
  OR_GATE U1688 ( .I1(n13672), .I2(n50), .O(n13674) );
  OR_GATE U1689 ( .I1(n12834), .I2(n12833), .O(n12836) );
  OR_GATE U1690 ( .I1(n6932), .I2(n982), .O(n6942) );
  INV_GATE U1691 ( .I1(n6933), .O(n982) );
  OR_GATE U1692 ( .I1(n983), .I2(n7048), .O(n7051) );
  INV_GATE U1693 ( .I1(n7049), .O(n983) );
  OR_GATE U1694 ( .I1(n14506), .I2(n984), .O(n14509) );
  INV_GATE U1695 ( .I1(n14507), .O(n984) );
  OR_GATE U1696 ( .I1(n10698), .I2(n985), .O(n10701) );
  INV_GATE U1697 ( .I1(n10699), .O(n985) );
  OR_GATE U1698 ( .I1(n986), .I2(n9867), .O(n9870) );
  INV_GATE U1699 ( .I1(n9868), .O(n986) );
  OR_GATE U1700 ( .I1(n2589), .I2(n987), .O(n2590) );
  INV_GATE U1701 ( .I1(n2588), .O(n987) );
  OR_GATE U1702 ( .I1(n2575), .I2(n988), .O(n2576) );
  INV_GATE U1703 ( .I1(n2574), .O(n988) );
  OR_GATE U1704 ( .I1(n8655), .I2(n791), .O(n8857) );
  AND_GATE U1705 ( .I1(n7168), .I2(n7169), .O(n989) );
  AND_GATE U1706 ( .I1(n8275), .I2(n8277), .O(n990) );
  AND_GATE U1707 ( .I1(n6397), .I2(n6396), .O(n991) );
  OR_GATE U1708 ( .I1(n89), .I2(n7070), .O(n7073) );
  OR_GATE U1709 ( .I1(n992), .I2(n7059), .O(n7062) );
  INV_GATE U1710 ( .I1(n7060), .O(n992) );
  OR_GATE U1711 ( .I1(n13898), .I2(n993), .O(n13901) );
  INV_GATE U1712 ( .I1(n13899), .O(n993) );
  OR_GATE U1713 ( .I1(n13032), .I2(n994), .O(n13035) );
  INV_GATE U1714 ( .I1(n13033), .O(n994) );
  OR_GATE U1715 ( .I1(n14581), .I2(n995), .O(n14584) );
  INV_GATE U1716 ( .I1(n14582), .O(n995) );
  OR_GATE U1717 ( .I1(n12127), .I2(n996), .O(n12130) );
  INV_GATE U1718 ( .I1(n12128), .O(n996) );
  OR_GATE U1719 ( .I1(n10242), .I2(n997), .O(n10245) );
  INV_GATE U1720 ( .I1(n10243), .O(n997) );
  OR_GATE U1721 ( .I1(n11128), .I2(n998), .O(n11131) );
  INV_GATE U1722 ( .I1(n11129), .O(n998) );
  OR_GATE U1723 ( .I1(n2561), .I2(n999), .O(n2562) );
  INV_GATE U1724 ( .I1(n2560), .O(n999) );
  AND_GATE U1725 ( .I1(n8648), .I2(n8650), .O(n1000) );
  OR_GATE U1726 ( .I1(n6866), .I2(n6860), .O(n6874) );
  OR_GATE U1727 ( .I1(n14335), .I2(n1001), .O(n14338) );
  INV_GATE U1728 ( .I1(n14336), .O(n1001) );
  OR_GATE U1729 ( .I1(n13480), .I2(n1002), .O(n13483) );
  INV_GATE U1730 ( .I1(n13481), .O(n1002) );
  OR_GATE U1731 ( .I1(n12602), .I2(n1003), .O(n12605) );
  INV_GATE U1732 ( .I1(n12603), .O(n1003) );
  OR_GATE U1733 ( .I1(n10747), .I2(n1004), .O(n10750) );
  INV_GATE U1734 ( .I1(n10748), .O(n1004) );
  OR_GATE U1735 ( .I1(n11602), .I2(n1005), .O(n11605) );
  INV_GATE U1736 ( .I1(n11603), .O(n1005) );
  OR_GATE U1737 ( .I1(n13884), .I2(n1006), .O(n13887) );
  INV_GATE U1738 ( .I1(n13885), .O(n1006) );
  OR_GATE U1739 ( .I1(n13017), .I2(n1007), .O(n13020) );
  INV_GATE U1740 ( .I1(n13018), .O(n1007) );
  OR_GATE U1741 ( .I1(n14607), .I2(n1008), .O(n14610) );
  INV_GATE U1742 ( .I1(n14608), .O(n1008) );
  OR_GATE U1743 ( .I1(n11152), .I2(n1009), .O(n11155) );
  INV_GATE U1744 ( .I1(n11153), .O(n1009) );
  OR_GATE U1745 ( .I1(n12001), .I2(n1010), .O(n12004) );
  INV_GATE U1746 ( .I1(n12002), .O(n1010) );
  OR_GATE U1747 ( .I1(n9224), .I2(n284), .O(n15331) );
  OR_GATE U1748 ( .I1(n156), .I2(n6538), .O(n6539) );
  OR_GATE U1749 ( .I1(n14320), .I2(n1011), .O(n14323) );
  INV_GATE U1750 ( .I1(n14321), .O(n1011) );
  OR_GATE U1751 ( .I1(n13465), .I2(n1012), .O(n13468) );
  INV_GATE U1752 ( .I1(n13466), .O(n1012) );
  OR_GATE U1753 ( .I1(n10772), .I2(n1013), .O(n10775) );
  INV_GATE U1754 ( .I1(n10773), .O(n1013) );
  OR_GATE U1755 ( .I1(n11627), .I2(n1014), .O(n11630) );
  INV_GATE U1756 ( .I1(n11628), .O(n1014) );
  OR_GATE U1757 ( .I1(n12476), .I2(n1015), .O(n12479) );
  INV_GATE U1758 ( .I1(n12477), .O(n1015) );
  OR_GATE U1759 ( .I1(n7842), .I2(n7841), .O(n7844) );
  OR_GATE U1760 ( .I1(n8770), .I2(n8769), .O(n8772) );
  OR_GATE U1761 ( .I1(n13869), .I2(n1016), .O(n13872) );
  INV_GATE U1762 ( .I1(n13870), .O(n1016) );
  OR_GATE U1763 ( .I1(n14633), .I2(n1017), .O(n14636) );
  INV_GATE U1764 ( .I1(n14634), .O(n1017) );
  OR_GATE U1765 ( .I1(n12026), .I2(n1018), .O(n12029) );
  INV_GATE U1766 ( .I1(n12027), .O(n1018) );
  OR_GATE U1767 ( .I1(n12891), .I2(n1019), .O(n12894) );
  INV_GATE U1768 ( .I1(n12892), .O(n1019) );
  OR_GATE U1769 ( .I1(n8337), .I2(n285), .O(n15328) );
  OR_GATE U1770 ( .I1(n14305), .I2(n1020), .O(n14308) );
  INV_GATE U1771 ( .I1(n14306), .O(n1020) );
  OR_GATE U1772 ( .I1(n12501), .I2(n1021), .O(n12504) );
  INV_GATE U1773 ( .I1(n12502), .O(n1021) );
  OR_GATE U1774 ( .I1(n13339), .I2(n1022), .O(n13342) );
  INV_GATE U1775 ( .I1(n13340), .O(n1022) );
  OR_GATE U1776 ( .I1(n12916), .I2(n1023), .O(n12919) );
  INV_GATE U1777 ( .I1(n12917), .O(n1023) );
  OR_GATE U1778 ( .I1(n13743), .I2(n1024), .O(n13746) );
  INV_GATE U1779 ( .I1(n13744), .O(n1024) );
  OR_GATE U1780 ( .I1(n14659), .I2(n1025), .O(n14662) );
  INV_GATE U1781 ( .I1(n14660), .O(n1025) );
  OR_GATE U1782 ( .I1(n472), .I2(n7873), .O(n7875) );
  OR_GATE U1783 ( .I1(n13364), .I2(n1026), .O(n13367) );
  INV_GATE U1784 ( .I1(n13365), .O(n1026) );
  OR_GATE U1785 ( .I1(n14179), .I2(n1027), .O(n14182) );
  INV_GATE U1786 ( .I1(n14180), .O(n1027) );
  OR_GATE U1787 ( .I1(n13768), .I2(n1028), .O(n13771) );
  INV_GATE U1788 ( .I1(n13769), .O(n1028) );
  OR_GATE U1789 ( .I1(n14684), .I2(n1029), .O(n14687) );
  INV_GATE U1790 ( .I1(n14685), .O(n1029) );
  OR_GATE U1791 ( .I1(n14204), .I2(n1030), .O(n14207) );
  INV_GATE U1792 ( .I1(n14205), .O(n1030) );
  OR_GATE U1793 ( .I1(n14709), .I2(n1031), .O(n14712) );
  INV_GATE U1794 ( .I1(n14710), .O(n1031) );
  OR_GATE U1795 ( .I1(n471), .I2(n7474), .O(n7475) );
  OR_GATE U1796 ( .I1(n10354), .I2(n1032), .O(n10015) );
  AND_GATE U1797 ( .I1(n10360), .I2(n860), .O(n1032) );
  OR_GATE U1798 ( .I1(n6606), .I2(n6609), .O(n7331) );
  OR_GATE U1799 ( .I1(n6961), .I2(n6960), .O(n6963) );
  OR_GATE U1800 ( .I1(n6894), .I2(n6899), .O(n6896) );
  OR_GATE U1801 ( .I1(n9817), .I2(n1033), .O(n9818) );
  AND_GATE U1802 ( .I1(n9271), .I2(n9270), .O(n1033) );
  OR_GATE U1803 ( .I1(n6928), .I2(n6933), .O(n6930) );
  OR_GATE U1804 ( .I1(n6791), .I2(n6783), .O(n6786) );
  OR_GATE U1805 ( .I1(n3587), .I2(n1034), .O(n3710) );
  OR_GATE U1806 ( .I1(n3972), .I2(n1035), .O(n4411) );
  INV_GATE U1807 ( .I1(n3974), .O(n1035) );
  OR_GATE U1808 ( .I1(n3956), .I2(n1036), .O(n4423) );
  INV_GATE U1809 ( .I1(n3958), .O(n1036) );
  OR_GATE U1810 ( .I1(n5290), .I2(n5295), .O(n5567) );
  OR_GATE U1811 ( .I1(n1037), .I2(n4474), .O(n4467) );
  INV_GATE U1812 ( .I1(n4476), .O(n1037) );
  OR_GATE U1813 ( .I1(n6128), .I2(n283), .O(n6945) );
  OR_GATE U1814 ( .I1(n6911), .I2(n6916), .O(n6913) );
  OR_GATE U1815 ( .I1(n392), .I2(n5261), .O(n5264) );
  OR_GATE U1816 ( .I1(n397), .I2(n4391), .O(n4394) );
  OR_GATE U1817 ( .I1(n1038), .I2(n5272), .O(n5275) );
  INV_GATE U1818 ( .I1(n5273), .O(n1038) );
  OR_GATE U1819 ( .I1(n584), .I2(n4401), .O(n4404) );
  OR_GATE U1820 ( .I1(n1039), .I2(n5283), .O(n5286) );
  INV_GATE U1821 ( .I1(n5284), .O(n1039) );
  OR_GATE U1822 ( .I1(n1040), .I2(n6275), .O(n6270) );
  INV_GATE U1823 ( .I1(n6272), .O(n1040) );
  OR_GATE U1824 ( .I1(n3578), .I2(n235), .O(n3580) );
  OR_GATE U1825 ( .I1(n681), .I2(n5303), .O(n5300) );
  OR_GATE U1826 ( .I1(n2704), .I2(n2706), .O(n2702) );
  OR_GATE U1827 ( .I1(n1041), .I2(n7269), .O(n7264) );
  INV_GATE U1828 ( .I1(n7266), .O(n1041) );
  NAND_GATE U1829 ( .I1(n7608), .I2(n229), .O(n1346) );
  OR_GATE U1830 ( .I1(n7619), .I2(n1042), .O(n7623) );
  AND_GATE U1831 ( .I1(n7620), .I2(n189), .O(n1042) );
  OR_GATE U1832 ( .I1(n1043), .I2(n8467), .O(n8470) );
  INV_GATE U1833 ( .I1(n8468), .O(n1043) );
  OR_GATE U1834 ( .I1(n527), .I2(n6697), .O(n6693) );
  OR_GATE U1835 ( .I1(n14010), .I2(n1044), .O(n14013) );
  AND_GATE U1836 ( .I1(n14012), .I2(n14011), .O(n1044) );
  OR_GATE U1837 ( .I1(n1212), .I2(n1045), .O(n9229) );
  AND_GATE U1838 ( .I1(n9233), .I2(n9199), .O(n1045) );
  OR_GATE U1839 ( .I1(n1248), .I2(n1046), .O(n9814) );
  AND_GATE U1840 ( .I1(n10038), .I2(n9477), .O(n1046) );
  OR_GATE U1841 ( .I1(n1355), .I2(n1047), .O(n7526) );
  AND_GATE U1842 ( .I1(n7624), .I2(n7345), .O(n1047) );
  OR_GATE U1843 ( .I1(n1252), .I2(n1048), .O(n10468) );
  AND_GATE U1844 ( .I1(n10506), .I2(n10505), .O(n1048) );
  OR_GATE U1845 ( .I1(n1267), .I2(n1049), .O(n15359) );
  AND_GATE U1846 ( .I1(n14016), .I2(n13576), .O(n1049) );
  OR_GATE U1847 ( .I1(n1302), .I2(n1050), .O(n6722) );
  AND_GATE U1848 ( .I1(n7365), .I2(n208), .O(n1050) );
  OR3_GATE U1849 ( .I1(n1051), .I2(n1052), .I3(n8916), .O(n9202) );
  INV_GATE U1850 ( .I1(n8917), .O(n1051) );
  AND_GATE U1851 ( .I1(n8915), .I2(n8907), .O(n1052) );
  OR_GATE U1852 ( .I1(n1360), .I2(n1053), .O(n8290) );
  AND_GATE U1853 ( .I1(n8271), .I2(n8272), .O(n1053) );
  OR_GATE U1854 ( .I1(n5882), .I2(n1054), .O(n6213) );
  INV_GATE U1855 ( .I1(n5884), .O(n1054) );
  OR_GATE U1856 ( .I1(n6251), .I2(n1055), .O(n6256) );
  INV_GATE U1857 ( .I1(n6252), .O(n1055) );
  OR_GATE U1858 ( .I1(n5327), .I2(n1056), .O(n5331) );
  INV_GATE U1859 ( .I1(n5328), .O(n1056) );
  OR_GATE U1860 ( .I1(n1057), .I2(n5753), .O(n5757) );
  INV_GATE U1861 ( .I1(n5754), .O(n1057) );
  OR_GATE U1862 ( .I1(n1250), .I2(n1058), .O(n7744) );
  AND_GATE U1863 ( .I1(n7730), .I2(n7453), .O(n1058) );
  OR_GATE U1864 ( .I1(n11038), .I2(n11039), .O(n11042) );
  OR_GATE U1865 ( .I1(n1059), .I2(n5205), .O(n5208) );
  INV_GATE U1866 ( .I1(n5206), .O(n1059) );
  OR_GATE U1867 ( .I1(n4330), .I2(n1060), .O(n4333) );
  INV_GATE U1868 ( .I1(n4329), .O(n1060) );
  OR_GATE U1869 ( .I1(n10039), .I2(n1061), .O(n10043) );
  AND_GATE U1870 ( .I1(n10040), .I2(n755), .O(n1061) );
  OR_GATE U1871 ( .I1(n3526), .I2(n1062), .O(n3529) );
  INV_GATE U1872 ( .I1(n3525), .O(n1062) );
  OR_GATE U1873 ( .I1(n3482), .I2(n1063), .O(n3485) );
  INV_GATE U1874 ( .I1(n3481), .O(n1063) );
  OR_GATE U1875 ( .I1(n3493), .I2(n1064), .O(n3496) );
  INV_GATE U1876 ( .I1(n3492), .O(n1064) );
  OR_GATE U1877 ( .I1(n3504), .I2(n1065), .O(n3507) );
  INV_GATE U1878 ( .I1(n3503), .O(n1065) );
  OR_GATE U1879 ( .I1(n1066), .I2(n7544), .O(n7547) );
  INV_GATE U1880 ( .I1(n7545), .O(n1066) );
  OR_GATE U1881 ( .I1(n5730), .I2(n1067), .O(n5717) );
  INV_GATE U1882 ( .I1(n6589), .O(n1067) );
  OR_GATE U1883 ( .I1(n3515), .I2(n1068), .O(n3518) );
  INV_GATE U1884 ( .I1(n3514), .O(n1068) );
  OR3_GATE U1885 ( .I1(n10983), .I2(n1069), .I3(n1070), .O(n10987) );
  AND_GATE U1886 ( .I1(n973), .I2(n10978), .O(n1069) );
  AND4_GATE U1887 ( .I1(n10981), .I2(n10980), .I3(n973), .I4(n10979), .O(n1070) );
  OR_GATE U1888 ( .I1(n1071), .I2(n6991), .O(n6995) );
  INV_GATE U1889 ( .I1(n6992), .O(n1071) );
  OR_GATE U1890 ( .I1(n1072), .I2(n9009), .O(n9012) );
  INV_GATE U1891 ( .I1(n9010), .O(n1072) );
  OR_GATE U1892 ( .I1(n1353), .I2(n1073), .O(n9849) );
  AND_GATE U1893 ( .I1(n9856), .I2(n9457), .O(n1073) );
  OR3_GATE U1894 ( .I1(n1074), .I2(n10655), .I3(n279), .O(n10659) );
  AND_GATE U1895 ( .I1(n10654), .I2(n10646), .O(n1074) );
  OR_GATE U1896 ( .I1(n5216), .I2(n1075), .O(n5219) );
  INV_GATE U1897 ( .I1(n5215), .O(n1075) );
  OR_GATE U1898 ( .I1(n1076), .I2(n5226), .O(n5229) );
  INV_GATE U1899 ( .I1(n5227), .O(n1076) );
  OR_GATE U1900 ( .I1(n1077), .I2(n5250), .O(n5253) );
  INV_GATE U1901 ( .I1(n5251), .O(n1077) );
  OR_GATE U1902 ( .I1(n2669), .I2(n1078), .O(n2672) );
  INV_GATE U1903 ( .I1(n2668), .O(n1078) );
  OR_GATE U1904 ( .I1(n3471), .I2(n1079), .O(n3474) );
  INV_GATE U1905 ( .I1(n3470), .O(n1079) );
  OR_GATE U1906 ( .I1(n2658), .I2(n1080), .O(n2661) );
  INV_GATE U1907 ( .I1(n2657), .O(n1080) );
  OR_GATE U1908 ( .I1(n2647), .I2(n1081), .O(n2650) );
  INV_GATE U1909 ( .I1(n2646), .O(n1081) );
  OR_GATE U1910 ( .I1(n2636), .I2(n1082), .O(n2639) );
  INV_GATE U1911 ( .I1(n2635), .O(n1082) );
  OR_GATE U1912 ( .I1(n2625), .I2(n1083), .O(n2628) );
  INV_GATE U1913 ( .I1(n2624), .O(n1083) );
  OR_GATE U1914 ( .I1(n1255), .I2(n1084), .O(n8257) );
  AND_GATE U1915 ( .I1(n8254), .I2(n8253), .O(n1084) );
  OR_GATE U1916 ( .I1(n1301), .I2(n1085), .O(n9254) );
  AND_GATE U1917 ( .I1(n9258), .I2(n9257), .O(n1085) );
  OR_GATE U1918 ( .I1(n7587), .I2(n7588), .O(n7600) );
  OR_GATE U1919 ( .I1(n1086), .I2(n4318), .O(n4321) );
  INV_GATE U1920 ( .I1(n4319), .O(n1086) );
  OR_GATE U1921 ( .I1(n1087), .I2(n3448), .O(n3451) );
  INV_GATE U1922 ( .I1(n3449), .O(n1087) );
  OR_GATE U1923 ( .I1(n2576), .I2(n1088), .O(n2578) );
  INV_GATE U1924 ( .I1(n2577), .O(n1088) );
  OR_GATE U1925 ( .I1(n1089), .I2(n9343), .O(n9346) );
  INV_GATE U1926 ( .I1(n9344), .O(n1089) );
  OR_GATE U1927 ( .I1(n2614), .I2(n1090), .O(n2617) );
  INV_GATE U1928 ( .I1(n2613), .O(n1090) );
  OR_GATE U1929 ( .I1(n5916), .I2(n5911), .O(n5926) );
  OR_GATE U1930 ( .I1(n1091), .I2(n5194), .O(n5197) );
  INV_GATE U1931 ( .I1(n5195), .O(n1091) );
  OR_GATE U1932 ( .I1(n4307), .I2(n1092), .O(n4310) );
  INV_GATE U1933 ( .I1(n4308), .O(n1092) );
  OR_GATE U1934 ( .I1(n1093), .I2(n3437), .O(n3440) );
  INV_GATE U1935 ( .I1(n3438), .O(n1093) );
  OR_GATE U1936 ( .I1(n1094), .I2(n3459), .O(n3462) );
  INV_GATE U1937 ( .I1(n3460), .O(n1094) );
  OR_GATE U1938 ( .I1(n2590), .I2(n1095), .O(n2592) );
  INV_GATE U1939 ( .I1(n2591), .O(n1095) );
  OR_GATE U1940 ( .I1(n2603), .I2(n1096), .O(n2606) );
  INV_GATE U1941 ( .I1(n2602), .O(n1096) );
  OR_GATE U1942 ( .I1(n2562), .I2(n1097), .O(n2564) );
  INV_GATE U1943 ( .I1(n2563), .O(n1097) );
  OR_GATE U1944 ( .I1(n9958), .I2(n1098), .O(n9961) );
  INV_GATE U1945 ( .I1(n9959), .O(n1098) );
  OR_GATE U1946 ( .I1(n1099), .I2(n3426), .O(n3429) );
  INV_GATE U1947 ( .I1(n3427), .O(n1099) );
  OR_GATE U1948 ( .I1(n1100), .I2(n4296), .O(n4299) );
  INV_GATE U1949 ( .I1(n4297), .O(n1100) );
  OR_GATE U1950 ( .I1(n1101), .I2(n5183), .O(n5186) );
  INV_GATE U1951 ( .I1(n5184), .O(n1101) );
  OR_GATE U1952 ( .I1(n1102), .I2(n6092), .O(n6095) );
  INV_GATE U1953 ( .I1(n6093), .O(n1102) );
  OR_GATE U1954 ( .I1(n10268), .I2(n1103), .O(n10271) );
  INV_GATE U1955 ( .I1(n10269), .O(n1103) );
  OR_GATE U1956 ( .I1(n2550), .I2(n1104), .O(n2553) );
  INV_GATE U1957 ( .I1(n2549), .O(n1104) );
  OR_GATE U1958 ( .I1(n11177), .I2(n1105), .O(n11180) );
  INV_GATE U1959 ( .I1(n11178), .O(n1105) );
  OR_GATE U1960 ( .I1(n1106), .I2(n4285), .O(n4288) );
  INV_GATE U1961 ( .I1(n4286), .O(n1106) );
  OR_GATE U1962 ( .I1(n1107), .I2(n5172), .O(n5175) );
  INV_GATE U1963 ( .I1(n5173), .O(n1107) );
  OR_GATE U1964 ( .I1(n1108), .I2(n6081), .O(n6084) );
  INV_GATE U1965 ( .I1(n6082), .O(n1108) );
  OR_GATE U1966 ( .I1(n11652), .I2(n1109), .O(n11655) );
  INV_GATE U1967 ( .I1(n11653), .O(n1109) );
  OR_GATE U1968 ( .I1(n3752), .I2(n1110), .O(n3755) );
  INV_GATE U1969 ( .I1(n3751), .O(n1110) );
  OR_GATE U1970 ( .I1(n290), .I2(n15366), .O(n14895) );
  OR_GATE U1971 ( .I1(n1111), .I2(n4274), .O(n4277) );
  INV_GATE U1972 ( .I1(n4275), .O(n1111) );
  OR_GATE U1973 ( .I1(n2539), .I2(n1112), .O(n2542) );
  INV_GATE U1974 ( .I1(n2538), .O(n1112) );
  OR_GATE U1975 ( .I1(n12051), .I2(n1113), .O(n12054) );
  INV_GATE U1976 ( .I1(n12052), .O(n1113) );
  OR_GATE U1977 ( .I1(n1114), .I2(n5161), .O(n5164) );
  INV_GATE U1978 ( .I1(n5162), .O(n1114) );
  OR_GATE U1979 ( .I1(n14910), .I2(n348), .O(n14912) );
  OR_GATE U1980 ( .I1(n12526), .I2(n1115), .O(n12529) );
  INV_GATE U1981 ( .I1(n12527), .O(n1115) );
  OR_GATE U1982 ( .I1(n12941), .I2(n1116), .O(n12944) );
  INV_GATE U1983 ( .I1(n12942), .O(n1116) );
  OR_GATE U1984 ( .I1(n3416), .I2(n1117), .O(n3419) );
  INV_GATE U1985 ( .I1(n3415), .O(n1117) );
  OR_GATE U1986 ( .I1(n13389), .I2(n1118), .O(n13392) );
  INV_GATE U1987 ( .I1(n13390), .O(n1118) );
  OR_GATE U1988 ( .I1(n2528), .I2(n1119), .O(n2531) );
  INV_GATE U1989 ( .I1(n2527), .O(n1119) );
  OR_GATE U1990 ( .I1(n13793), .I2(n1120), .O(n13796) );
  INV_GATE U1991 ( .I1(n13794), .O(n1120) );
  OR_GATE U1992 ( .I1(n14229), .I2(n1121), .O(n14232) );
  INV_GATE U1993 ( .I1(n14230), .O(n1121) );
  OR_GATE U1994 ( .I1(n1122), .I2(n5150), .O(n5153) );
  INV_GATE U1995 ( .I1(n5151), .O(n1122) );
  OR_GATE U1996 ( .I1(n4264), .I2(n1123), .O(n4267) );
  INV_GATE U1997 ( .I1(n4263), .O(n1123) );
  OR_GATE U1998 ( .I1(n14734), .I2(n1124), .O(n14737) );
  INV_GATE U1999 ( .I1(n14735), .O(n1124) );
  OR_GATE U2000 ( .I1(n1125), .I2(n3405), .O(n3408) );
  INV_GATE U2001 ( .I1(n3404), .O(n1125) );
  OR_GATE U2002 ( .I1(n2517), .I2(n1126), .O(n2520) );
  INV_GATE U2003 ( .I1(n2516), .O(n1126) );
  OR_GATE U2004 ( .I1(n4253), .I2(n1127), .O(n4256) );
  INV_GATE U2005 ( .I1(n4252), .O(n1127) );
  OR_GATE U2006 ( .I1(n3394), .I2(n1128), .O(n3397) );
  INV_GATE U2007 ( .I1(n3393), .O(n1128) );
  OR_GATE U2008 ( .I1(n2506), .I2(n1129), .O(n2509) );
  INV_GATE U2009 ( .I1(n2505), .O(n1129) );
  OR_GATE U2010 ( .I1(n4242), .I2(n1130), .O(n4245) );
  INV_GATE U2011 ( .I1(n4241), .O(n1130) );
  OR_GATE U2012 ( .I1(n3383), .I2(n1131), .O(n3386) );
  INV_GATE U2013 ( .I1(n3382), .O(n1131) );
  OR_GATE U2014 ( .I1(n2857), .I2(n1132), .O(n2860) );
  INV_GATE U2015 ( .I1(n2856), .O(n1132) );
  OR_GATE U2016 ( .I1(n1133), .I2(n3371), .O(n3374) );
  INV_GATE U2017 ( .I1(n3372), .O(n1133) );
  OR_GATE U2018 ( .I1(n2495), .I2(n1134), .O(n2498) );
  INV_GATE U2019 ( .I1(n2494), .O(n1134) );
  OR_GATE U2020 ( .I1(n3361), .I2(n1135), .O(n3364) );
  INV_GATE U2021 ( .I1(n3360), .O(n1135) );
  OR_GATE U2022 ( .I1(n1136), .I2(n2484), .O(n2487) );
  INV_GATE U2023 ( .I1(n2483), .O(n1136) );
  OR_GATE U2024 ( .I1(n2473), .I2(n1137), .O(n2476) );
  INV_GATE U2025 ( .I1(n2472), .O(n1137) );
  OR_GATE U2026 ( .I1(n2462), .I2(n1138), .O(n2465) );
  INV_GATE U2027 ( .I1(n2461), .O(n1138) );
  OR_GATE U2028 ( .I1(n5814), .I2(n5820), .O(n5826) );
  AND_GATE U2029 ( .I1(n3677), .I2(n3676), .O(n1139) );
  OR_GATE U2030 ( .I1(n5980), .I2(n5985), .O(n5982) );
  OR_GATE U2031 ( .I1(n5946), .I2(n5951), .O(n5948) );
  OR_GATE U2032 ( .I1(n5929), .I2(n5934), .O(n5931) );
  OR_GATE U2033 ( .I1(n5844), .I2(n872), .O(n6224) );
  OR_GATE U2034 ( .I1(n3036), .I2(n1140), .O(n3035) );
  INV_GATE U2035 ( .I1(n3039), .O(n1140) );
  OR_GATE U2036 ( .I1(n5655), .I2(n5653), .O(n5784) );
  OR_GATE U2037 ( .I1(n215), .I2(n2905), .O(n2907) );
  AND_GATE U2038 ( .I1(n5538), .I2(n5539), .O(n1141) );
  AND_GATE U2039 ( .I1(n4561), .I2(n3895), .O(n1142) );
  AND_GATE U2040 ( .I1(n2800), .I2(n2801), .O(n1143) );
  OR_GATE U2041 ( .I1(n6232), .I2(n6233), .O(n6239) );
  OR_GATE U2042 ( .I1(n871), .I2(n2997), .O(n3005) );
  OR_GATE U2043 ( .I1(n3011), .I2(n873), .O(n3018) );
  OR_GATE U2044 ( .I1(n5997), .I2(n6002), .O(n5999) );
  OR_GATE U2045 ( .I1(n5963), .I2(n5968), .O(n5965) );
  OR_GATE U2046 ( .I1(n1144), .I2(n6199), .O(n6202) );
  INV_GATE U2047 ( .I1(n6200), .O(n1144) );
  OR_GATE U2048 ( .I1(n1145), .I2(n6166), .O(n6169) );
  INV_GATE U2049 ( .I1(n6167), .O(n1145) );
  OR_GATE U2050 ( .I1(n6156), .I2(n1146), .O(n6159) );
  INV_GATE U2051 ( .I1(n6155), .O(n1146) );
  OR_GATE U2052 ( .I1(n6145), .I2(n1147), .O(n6148) );
  INV_GATE U2053 ( .I1(n6144), .O(n1147) );
  OR_GATE U2054 ( .I1(n3537), .I2(n223), .O(n3540) );
  OR_GATE U2055 ( .I1(n6372), .I2(n6371), .O(n6374) );
  OR_GATE U2056 ( .I1(n6477), .I2(n6478), .O(n6480) );
  OR_GATE U2057 ( .I1(n6244), .I2(n1148), .O(n6243) );
  INV_GATE U2058 ( .I1(n6247), .O(n1148) );
  OR_GATE U2059 ( .I1(n3645), .I2(n3649), .O(n3643) );
  OR_GATE U2060 ( .I1(n277), .I2(n4833), .O(n4828) );
  OR_GATE U2061 ( .I1(n5696), .I2(n5695), .O(n5697) );
  OR_GATE U2062 ( .I1(n2735), .I2(n2734), .O(n2737) );
  OR_GATE U2063 ( .I1(n1149), .I2(n7555), .O(n7558) );
  INV_GATE U2064 ( .I1(n7556), .O(n1149) );
  OR_GATE U2065 ( .I1(n6411), .I2(n6410), .O(n6413) );
  OR_GATE U2066 ( .I1(n3027), .I2(n1150), .O(n3039) );
  OR_GATE U2067 ( .I1(n5034), .I2(n5033), .O(n5036) );
  OR_GATE U2068 ( .I1(n5625), .I2(n5621), .O(n5892) );
  AND_GATE U2069 ( .I1(n4849), .I2(n4848), .O(n1151) );
  OR_GATE U2070 ( .I1(n5856), .I2(n541), .O(n5868) );
  OR_GATE U2071 ( .I1(n3672), .I2(n3671), .O(n3680) );
  AND_GATE U2072 ( .I1(n3921), .I2(n3920), .O(n1152) );
  OR_GATE U2073 ( .I1(n4873), .I2(n4877), .O(n5314) );
  OR_GATE U2074 ( .I1(n4076), .I2(n4075), .O(n4078) );
  OR_GATE U2075 ( .I1(n4060), .I2(n4059), .O(n4062) );
  AND_GATE U2076 ( .I1(n2959), .I2(n2958), .O(n1153) );
  OR_GATE U2077 ( .I1(n4044), .I2(n4043), .O(n4046) );
  OR_GATE U2078 ( .I1(n3966), .I2(n3963), .O(n3974) );
  OR_GATE U2079 ( .I1(n4028), .I2(n4027), .O(n4030) );
  OR_GATE U2080 ( .I1(n4012), .I2(n4011), .O(n4014) );
  OR_GATE U2081 ( .I1(n3950), .I2(n3947), .O(n3958) );
  OR_GATE U2082 ( .I1(n2990), .I2(n839), .O(n3684) );
  AND_GATE U2083 ( .I1(n3812), .I2(n3813), .O(n1154) );
  OR_GATE U2084 ( .I1(n2996), .I2(n1155), .O(n3004) );
  INV_GATE U2085 ( .I1(n2997), .O(n1155) );
  AND_GATE U2086 ( .I1(n4594), .I2(n4593), .O(n1156) );
  AND_GATE U2087 ( .I1(n4787), .I2(n4786), .O(n1157) );
  OR_GATE U2088 ( .I1(n5878), .I2(n5875), .O(n5884) );
  OR_GATE U2089 ( .I1(n1158), .I2(n6188), .O(n6191) );
  INV_GATE U2090 ( .I1(n6189), .O(n1158) );
  OR_GATE U2091 ( .I1(n6134), .I2(n1159), .O(n6137) );
  INV_GATE U2092 ( .I1(n6133), .O(n1159) );
  OR_GATE U2093 ( .I1(n1160), .I2(n8131), .O(n8134) );
  INV_GATE U2094 ( .I1(n8132), .O(n1160) );
  OR_GATE U2095 ( .I1(n5899), .I2(n5895), .O(n5909) );
  OR_GATE U2096 ( .I1(n5002), .I2(n5001), .O(n5004) );
  OR_GATE U2097 ( .I1(n4706), .I2(n4705), .O(n4708) );
  OR_GATE U2098 ( .I1(n4984), .I2(n4983), .O(n4986) );
  OR_GATE U2099 ( .I1(n4968), .I2(n4967), .O(n4970) );
  OR_GATE U2100 ( .I1(n3048), .I2(n3044), .O(n3057) );
  OR_GATE U2101 ( .I1(n3098), .I2(n3097), .O(n3100) );
  OR_GATE U2102 ( .I1(n3114), .I2(n3113), .O(n3116) );
  OR_GATE U2103 ( .I1(n3130), .I2(n3129), .O(n3132) );
  OR_GATE U2104 ( .I1(n3146), .I2(n3145), .O(n3148) );
  AND_GATE U2105 ( .I1(n5779), .I2(n5778), .O(n1161) );
  AND_GATE U2106 ( .I1(n5509), .I2(n5508), .O(n1162) );
  OR_GATE U2107 ( .I1(n6001), .I2(n1163), .O(n6011) );
  INV_GATE U2108 ( .I1(n6002), .O(n1163) );
  OR_GATE U2109 ( .I1(n1164), .I2(n6177), .O(n6180) );
  INV_GATE U2110 ( .I1(n6178), .O(n1164) );
  AND_GATE U2111 ( .I1(n6433), .I2(n6432), .O(n1165) );
  OR_GATE U2112 ( .I1(n6017), .I2(n6016), .O(n6019) );
  OR_GATE U2113 ( .I1(n4092), .I2(n4091), .O(n4094) );
  OR_GATE U2114 ( .I1(n3162), .I2(n3161), .O(n3164) );
  OR_GATE U2115 ( .I1(n1166), .I2(n8478), .O(n8481) );
  INV_GATE U2116 ( .I1(n8479), .O(n1166) );
  OR_GATE U2117 ( .I1(n1167), .I2(n9020), .O(n9023) );
  INV_GATE U2118 ( .I1(n9021), .O(n1167) );
  OR_GATE U2119 ( .I1(n6013), .I2(n1168), .O(n6106) );
  INV_GATE U2120 ( .I1(n6016), .O(n1168) );
  OR_GATE U2121 ( .I1(n3229), .I2(n3228), .O(n3231) );
  OR_GATE U2122 ( .I1(n9393), .I2(n1169), .O(n9396) );
  INV_GATE U2123 ( .I1(n9394), .O(n1169) );
  OR_GATE U2124 ( .I1(n9943), .I2(n1170), .O(n9946) );
  INV_GATE U2125 ( .I1(n9944), .O(n1170) );
  OR_GATE U2126 ( .I1(n10294), .I2(n1171), .O(n10297) );
  INV_GATE U2127 ( .I1(n10295), .O(n1171) );
  OR_GATE U2128 ( .I1(n5084), .I2(n5083), .O(n5086) );
  OR_GATE U2129 ( .I1(n10797), .I2(n1172), .O(n10800) );
  INV_GATE U2130 ( .I1(n10798), .O(n1172) );
  OR_GATE U2131 ( .I1(n3245), .I2(n3244), .O(n3247) );
  OR_GATE U2132 ( .I1(n4160), .I2(n4159), .O(n4162) );
  OR_GATE U2133 ( .I1(n3261), .I2(n3260), .O(n3263) );
  OR_GATE U2134 ( .I1(n5117), .I2(n5116), .O(n5119) );
  OR_GATE U2135 ( .I1(n4176), .I2(n4175), .O(n4178) );
  OR_GATE U2136 ( .I1(n14933), .I2(n21), .O(n14935) );
  OR_GATE U2137 ( .I1(n2878), .I2(n2877), .O(n2880) );
  OR_GATE U2138 ( .I1(n5133), .I2(n5132), .O(n5135) );
  OR_GATE U2139 ( .I1(n4192), .I2(n4191), .O(n4194) );
  OR_GATE U2140 ( .I1(n3279), .I2(n3278), .O(n3281) );
  OR_GATE U2141 ( .I1(n286), .I2(n4699), .O(n4700) );
  OR_GATE U2142 ( .I1(n4208), .I2(n4207), .O(n4210) );
  OR_GATE U2143 ( .I1(n4224), .I2(n4223), .O(n4226) );
  OR_GATE U2144 ( .I1(n3311), .I2(n3310), .O(n3313) );
  OR_GATE U2145 ( .I1(n287), .I2(n3770), .O(n3771) );
  OR_GATE U2146 ( .I1(n3327), .I2(n3326), .O(n3329) );
  OR_GATE U2147 ( .I1(n3343), .I2(n3342), .O(n3345) );
  OR_GATE U2148 ( .I1(n288), .I2(n2871), .O(n2872) );
  OR_GATE U2149 ( .I1(n4540), .I2(n4539), .O(n4543) );
  OR3_GATE U2150 ( .I1(n1307), .I2(n2003), .I3(n2795), .O(n2742) );
  OR3_GATE U2151 ( .I1(n1173), .I2(n1174), .I3(n4736), .O(n4787) );
  INV_GATE U2152 ( .I1(n4737), .O(n1173) );
  AND_GATE U2153 ( .I1(n4735), .I2(n4729), .O(n1174) );
  OR_GATE U2154 ( .I1(n4766), .I2(n4765), .O(n4770) );
  OR3_GATE U2155 ( .I1(n1263), .I2(n3919), .I3(n3915), .O(n3920) );
  OR_GATE U2156 ( .I1(n4448), .I2(n1175), .O(n4450) );
  INV_GATE U2157 ( .I1(n4449), .O(n1175) );
  NAND3_GATE U2158 ( .I1(n5767), .I2(n5766), .I3(n823), .O(n5779) );
  OR_GATE U2159 ( .I1(n5412), .I2(n5413), .O(n5415) );
  OR_GATE U2160 ( .I1(n5665), .I2(n5664), .O(n5667) );
  OR_GATE U2161 ( .I1(n5694), .I2(n1176), .O(n5699) );
  AND_GATE U2162 ( .I1(n5696), .I2(n5695), .O(n1176) );
  OR_GATE U2163 ( .I1(n2938), .I2(n2939), .O(n2941) );
  OR_GATE U2164 ( .I1(n3619), .I2(n3620), .O(n3622) );
  OR_GATE U2165 ( .I1(n1351), .I2(n1177), .O(n5710) );
  AND_GATE U2166 ( .I1(n5700), .I2(n5441), .O(n1177) );
  OR_GATE U2167 ( .I1(n5992), .I2(n1178), .O(n5988) );
  INV_GATE U2168 ( .I1(n5994), .O(n1178) );
  OR_GATE U2169 ( .I1(n5941), .I2(n1179), .O(n5937) );
  INV_GATE U2170 ( .I1(n5943), .O(n1179) );
  OR_GATE U2171 ( .I1(n5688), .I2(n5681), .O(n6332) );
  OR_GATE U2172 ( .I1(n4742), .I2(n4752), .O(n5407) );
  OR3_GATE U2173 ( .I1(n3798), .I2(n1303), .I3(n3793), .O(n3800) );
  OR_GATE U2174 ( .I1(n5975), .I2(n1180), .O(n5971) );
  INV_GATE U2175 ( .I1(n5977), .O(n1180) );
  OR_GATE U2176 ( .I1(n5958), .I2(n1181), .O(n5954) );
  INV_GATE U2177 ( .I1(n5960), .O(n1181) );
  AND_GATE U2178 ( .I1(n3632), .I2(n3869), .O(n1182) );
  OR_GATE U2179 ( .I1(n11202), .I2(n1183), .O(n11205) );
  INV_GATE U2180 ( .I1(n11203), .O(n1183) );
  OR_GATE U2181 ( .I1(n11677), .I2(n1184), .O(n11680) );
  INV_GATE U2182 ( .I1(n11678), .O(n1184) );
  OR_GATE U2183 ( .I1(n12076), .I2(n1185), .O(n12079) );
  INV_GATE U2184 ( .I1(n12077), .O(n1185) );
  OR_GATE U2185 ( .I1(n12551), .I2(n1186), .O(n12554) );
  INV_GATE U2186 ( .I1(n12552), .O(n1186) );
  OR_GATE U2187 ( .I1(n12966), .I2(n1187), .O(n12969) );
  INV_GATE U2188 ( .I1(n12967), .O(n1187) );
  OR_GATE U2189 ( .I1(n13414), .I2(n1188), .O(n13417) );
  INV_GATE U2190 ( .I1(n13415), .O(n1188) );
  OR_GATE U2191 ( .I1(n13818), .I2(n1189), .O(n13821) );
  INV_GATE U2192 ( .I1(n13819), .O(n1189) );
  OR_GATE U2193 ( .I1(n14254), .I2(n1190), .O(n14257) );
  INV_GATE U2194 ( .I1(n14255), .O(n1190) );
  OR_GATE U2195 ( .I1(n14759), .I2(n1191), .O(n14762) );
  INV_GATE U2196 ( .I1(n14760), .O(n1191) );
  OR_GATE U2197 ( .I1(n1193), .I2(n2786), .O(n2789) );
  OR_GATE U2198 ( .I1(n6358), .I2(n6349), .O(n6621) );
  AND_GATE U2199 ( .I1(n2020), .I2(n2019), .O(n1194) );
  OR_GATE U2200 ( .I1(n11214), .I2(n11213), .O(n11216) );
  OR_GATE U2201 ( .I1(n11689), .I2(n11688), .O(n11691) );
  OR_GATE U2202 ( .I1(n12088), .I2(n12087), .O(n12090) );
  OR_GATE U2203 ( .I1(n12563), .I2(n12562), .O(n12565) );
  OR_GATE U2204 ( .I1(n12978), .I2(n12977), .O(n12980) );
  OR_GATE U2205 ( .I1(n13426), .I2(n13425), .O(n13428) );
  OR_GATE U2206 ( .I1(n13830), .I2(n13829), .O(n13832) );
  OR_GATE U2207 ( .I1(n14266), .I2(n14265), .O(n14268) );
  OR_GATE U2208 ( .I1(n14771), .I2(n14770), .O(n14773) );
  OR_GATE U2209 ( .I1(n1411), .I2(n1195), .O(n15138) );
  INV_GATE U2210 ( .I1(B[0]), .O(n1195) );
  OR_GATE U2211 ( .I1(n1415), .I2(n1195), .O(n15080) );
  OR_GATE U2212 ( .I1(n6351), .I2(n6359), .O(n6353) );
  OR_GATE U2213 ( .I1(A[29]), .I2(n1397), .O(n1932) );
  OR_GATE U2214 ( .I1(n1197), .I2(n9856), .O(n9858) );
  INV_GATE U2215 ( .I1(n9853), .O(n1197) );
  OR_GATE U2216 ( .I1(n860), .I2(n10354), .O(n10357) );
  OR_GATE U2217 ( .I1(n746), .I2(n8975), .O(n8976) );
  OR_GATE U2218 ( .I1(n1198), .I2(n9689), .O(n9684) );
  INV_GATE U2219 ( .I1(n9686), .O(n1198) );
  OR_GATE U2220 ( .I1(n9299), .I2(n844), .O(n9298) );
  OR_GATE U2221 ( .I1(n5431), .I2(n1199), .O(n5428) );
  INV_GATE U2222 ( .I1(n5436), .O(n1199) );
  AND3_GATE U2223 ( .I1(n8953), .I2(n8590), .I3(n8947), .O(n1200) );
  INV_GATE U2224 ( .I1(n1200), .O(n9160) );
  AND_GATE U2225 ( .I1(n13571), .I2(n13570), .O(n1201) );
  AND_GATE U2226 ( .I1(n11045), .I2(n11044), .O(n1202) );
  AND_GATE U2227 ( .I1(n9297), .I2(n9296), .O(n1203) );
  AND_GATE U2228 ( .I1(n8433), .I2(n8432), .O(n1204) );
  AND3_GATE U2229 ( .I1(n7529), .I2(n7528), .I3(n7527), .O(n1205) );
  AND3_GATE U2230 ( .I1(n5730), .I2(n5729), .I3(n5728), .O(n1206) );
  AND_GATE U2231 ( .I1(n7243), .I2(n7242), .O(n1207) );
  NAND_GATE U2232 ( .I1(n10454), .I2(n1210), .O(n1208) );
  AND_GATE U2233 ( .I1(n10453), .I2(n10457), .O(n1210) );
  NAND_GATE U2234 ( .I1(n1211), .I2(n7976), .O(n7975) );
  NOR_GATE U2235 ( .I1(n7980), .I2(n7978), .O(n1211) );
  OR_GATE U2236 ( .I1(n5360), .I2(n856), .O(n4851) );
  OR_GATE U2237 ( .I1(n10421), .I2(n15), .O(n10569) );
  NOR_GATE U2238 ( .I1(n9764), .I2(n9232), .O(n1212) );
  OR3_GATE U2239 ( .I1(n14450), .I2(n592), .I3(n14449), .O(n14447) );
  OR_GATE U2240 ( .I1(n6474), .I2(n653), .O(n6469) );
  OR_GATE U2241 ( .I1(n772), .I2(n8405), .O(n8400) );
  AND_GATE U2242 ( .I1(n7494), .I2(n7492), .O(n1214) );
  INV_GATE U2243 ( .I1(n1214), .O(n8283) );
  OR_GATE U2244 ( .I1(n260), .I2(n7491), .O(n7490) );
  NAND_GATE U2245 ( .I1(n15352), .I2(n1217), .O(n1215) );
  NAND_GATE U2246 ( .I1(n1215), .I2(n1216), .O(\A2[37] ) );
  OR_GATE U2247 ( .I1(n16), .I2(n15354), .O(n1216) );
  AND_GATE U2248 ( .I1(n15353), .I2(n15355), .O(n1217) );
  AND_GATE U2249 ( .I1(n1218), .I2(n1219), .O(n12255) );
  INV_GATE U2250 ( .I1(n15351), .O(n1220) );
  AND_GATE U2251 ( .I1(n10951), .I2(n10950), .O(n1221) );
  NAND_GATE U2252 ( .I1(n7479), .I2(n1224), .O(n1222) );
  AND_GATE U2253 ( .I1(n1222), .I2(n1223), .O(n8031) );
  OR_GATE U2254 ( .I1(n8030), .I2(n8024), .O(n1223) );
  AND_GATE U2255 ( .I1(n8023), .I2(n7712), .O(n1224) );
  NAND_GATE U2256 ( .I1(n9541), .I2(n1227), .O(n1225) );
  AND_GATE U2257 ( .I1(n1225), .I2(n1226), .O(n9732) );
  OR_GATE U2258 ( .I1(n9730), .I2(n9718), .O(n1226) );
  AND_GATE U2259 ( .I1(n9717), .I2(n9723), .O(n1227) );
  AND_GATE U2260 ( .I1(n5542), .I2(n5541), .O(n1228) );
  AND3_GATE U2261 ( .I1(n7331), .I2(n7330), .I3(n7329), .O(n1229) );
  NAND_GATE U2262 ( .I1(n11889), .I2(n1233), .O(n1230) );
  AND_GATE U2263 ( .I1(n1230), .I2(n1231), .O(n12222) );
  OR_GATE U2264 ( .I1(n1232), .I2(n12338), .O(n1231) );
  INV_GATE U2265 ( .I1(n12339), .O(n1232) );
  AND_GATE U2266 ( .I1(n11890), .I2(n12339), .O(n1233) );
  NAND_GATE U2267 ( .I1(n244), .I2(n1236), .O(n1234) );
  AND_GATE U2268 ( .I1(n1234), .I2(n1235), .O(n10916) );
  AND_GATE U2269 ( .I1(n669), .I2(n11008), .O(n1236) );
  NAND_GATE U2270 ( .I1(n1237), .I2(n9248), .O(n9250) );
  NOR_GATE U2271 ( .I1(n9244), .I2(n9245), .O(n1237) );
  AND_GATE U2272 ( .I1(n4809), .I2(n4808), .O(n1238) );
  AND_GATE U2273 ( .I1(n11488), .I2(n11487), .O(n1239) );
  AND3_GATE U2274 ( .I1(n7506), .I2(n7505), .I3(n7504), .O(n1240) );
  OR_GATE U2275 ( .I1(n2738), .I2(n2735), .O(n2730) );
  NOR_GATE U2276 ( .I1(n1269), .I2(n1243), .O(n1242) );
  INV_GATE U2277 ( .I1(n1242), .O(n10475) );
  AND_GATE U2278 ( .I1(n10463), .I2(n10108), .O(n1243) );
  NOR3_GATE U2279 ( .I1(n1363), .I2(n1245), .I3(n1246), .O(n1244) );
  INV_GATE U2280 ( .I1(n1244), .O(n5532) );
  AND3_GATE U2281 ( .I1(n5518), .I2(n5524), .I3(n5523), .O(n1245) );
  AND3_GATE U2282 ( .I1(n5522), .I2(n5524), .I3(n5523), .O(n1246) );
  AND3_GATE U2283 ( .I1(n6542), .I2(n6467), .I3(n6466), .O(n1247) );
  INV_GATE U2284 ( .I1(n1247), .O(n6742) );
  NOR_GATE U2285 ( .I1(n10040), .I2(n10039), .O(n1248) );
  OR_GATE U2286 ( .I1(n1249), .I2(n14469), .O(n14471) );
  AND3_GATE U2287 ( .I1(n14038), .I2(n14036), .I3(n14037), .O(n1249) );
  OR_GATE U2288 ( .I1(n858), .I2(n7723), .O(n7724) );
  NOR_GATE U2289 ( .I1(n7734), .I2(n7732), .O(n1250) );
  OR_GATE U2290 ( .I1(n10971), .I2(n1294), .O(n10970) );
  AND_GATE U2291 ( .I1(n10973), .I2(n10972), .O(n1251) );
  INV_GATE U2292 ( .I1(n1251), .O(n15345) );
  NOR_GATE U2293 ( .I1(n10506), .I2(n1253), .O(n1252) );
  AND_GATE U2294 ( .I1(n10465), .I2(n10464), .O(n1253) );
  OR_GATE U2295 ( .I1(n1254), .I2(n6725), .O(n6726) );
  INV_GATE U2296 ( .I1(n7376), .O(n1254) );
  OR3_GATE U2297 ( .I1(n8272), .I2(n1360), .I3(n8274), .O(n8277) );
  AND_GATE U2298 ( .I1(n7682), .I2(n7681), .O(n1255) );
  OR_GATE U2299 ( .I1(n6786), .I2(n1257), .O(n6794) );
  OR_GATE U2300 ( .I1(n17), .I2(n4888), .O(n4891) );
  AND3_GATE U2301 ( .I1(n7667), .I2(n7364), .I3(n7668), .O(n1256) );
  INV_GATE U2302 ( .I1(n1256), .O(n7684) );
  OR_GATE U2303 ( .I1(n3793), .I2(n1303), .O(n3797) );
  AND_GATE U2304 ( .I1(n6768), .I2(n6498), .O(n1257) );
  INV_GATE U2305 ( .I1(n1257), .O(n6787) );
  OR_GATE U2306 ( .I1(n6783), .I2(n1257), .O(n6782) );
  OR_GATE U2307 ( .I1(n780), .I2(n3933), .O(n3931) );
  OR_GATE U2308 ( .I1(n8074), .I2(n1258), .O(n8070) );
  INV_GATE U2309 ( .I1(n8073), .O(n1258) );
  AND3_GATE U2310 ( .I1(n10637), .I2(n10389), .I3(n10642), .O(n1259) );
  INV_GATE U2311 ( .I1(n1259), .O(n10902) );
  INV_GATE U2312 ( .I1(n14937), .O(n1260) );
  AND_GATE U2313 ( .I1(n8200), .I2(n8205), .O(n1261) );
  INV_GATE U2314 ( .I1(n1261), .O(n8437) );
  NOR_GATE U2315 ( .I1(n2976), .I2(n2971), .O(n1262) );
  INV_GATE U2316 ( .I1(n1262), .O(n2972) );
  OR_GATE U2317 ( .I1(n804), .I2(n2726), .O(n2721) );
  NOR_GATE U2318 ( .I1(n3703), .I2(n3702), .O(n1263) );
  AND_GATE U2319 ( .I1(n13233), .I2(n13232), .O(n1264) );
  INV_GATE U2320 ( .I1(n1264), .O(n13630) );
  OR_GATE U2321 ( .I1(n1265), .I2(n13584), .O(n13585) );
  INV_GATE U2322 ( .I1(n15359), .O(n1265) );
  AND3_GATE U2323 ( .I1(n12369), .I2(n12217), .I3(n12216), .O(n1266) );
  NOR_GATE U2324 ( .I1(n14012), .I2(n14010), .O(n1267) );
  OR_GATE U2325 ( .I1(n15365), .I2(n1308), .O(n14455) );
  OR_GATE U2326 ( .I1(n6507), .I2(n1268), .O(n6510) );
  AND_GATE U2327 ( .I1(n5868), .I2(n5867), .O(n1268) );
  INV_GATE U2328 ( .I1(n1268), .O(n6506) );
  NOR_GATE U2329 ( .I1(n10465), .I2(n10506), .O(n1269) );
  NAND_GATE U2330 ( .I1(n1316), .I2(n1317), .O(n1271) );
  AND_GATE U2331 ( .I1(n14968), .I2(n1350), .O(n1272) );
  NAND_GATE U2332 ( .I1(n1273), .I2(n14365), .O(n14363) );
  NOR_GATE U2333 ( .I1(n14366), .I2(n14367), .O(n1273) );
  NAND_GATE U2334 ( .I1(n1274), .I2(n13510), .O(n13508) );
  NOR_GATE U2335 ( .I1(n13511), .I2(n13512), .O(n1274) );
  NAND_GATE U2336 ( .I1(n1275), .I2(n12633), .O(n12631) );
  NOR_GATE U2337 ( .I1(n12634), .I2(n12635), .O(n1275) );
  NAND_GATE U2338 ( .I1(n1276), .I2(n11744), .O(n11742) );
  NOR_GATE U2339 ( .I1(n11745), .I2(n11746), .O(n1276) );
  NAND_GATE U2340 ( .I1(n1277), .I2(n8998), .O(n8997) );
  NOR_GATE U2341 ( .I1(n9000), .I2(n8999), .O(n1277) );
  NAND_GATE U2342 ( .I1(n1278), .I2(n8120), .O(n8118) );
  NOR_GATE U2343 ( .I1(n8122), .I2(n8121), .O(n1278) );
  NAND_GATE U2344 ( .I1(n1279), .I2(n7278), .O(n7276) );
  NOR_GATE U2345 ( .I1(n7280), .I2(n7279), .O(n1279) );
  AND_GATE U2346 ( .I1(n14833), .I2(n14989), .O(n1280) );
  AND_GATE U2347 ( .I1(n14827), .I2(n15027), .O(n1281) );
  AND_GATE U2348 ( .I1(n14551), .I2(n14550), .O(n1282) );
  AND_GATE U2349 ( .I1(n13679), .I2(n13678), .O(n1283) );
  AND_GATE U2350 ( .I1(n12842), .I2(n12841), .O(n1284) );
  AND_GATE U2351 ( .I1(n11970), .I2(n11969), .O(n1285) );
  AND_GATE U2352 ( .I1(n11111), .I2(n11110), .O(n1286) );
  AND_GATE U2353 ( .I1(n7600), .I2(n7599), .O(n1287) );
  AND_GATE U2354 ( .I1(n6651), .I2(n6650), .O(n1288) );
  OR_GATE U2355 ( .I1(n1289), .I2(n5358), .O(n5367) );
  INV_GATE U2356 ( .I1(n5359), .O(n1289) );
  AND3_GATE U2357 ( .I1(n7215), .I2(n6715), .I3(n7214), .O(n1290) );
  INV_GATE U2358 ( .I1(n1290), .O(n7189) );
  OR_GATE U2359 ( .I1(n8291), .I2(n1360), .O(n8279) );
  NOR3_GATE U2360 ( .I1(n1292), .I2(n1293), .I3(n12328), .O(n1291) );
  INV_GATE U2361 ( .I1(n12329), .O(n1292) );
  AND_GATE U2362 ( .I1(n12327), .I2(n12326), .O(n1293) );
  NOR_GATE U2363 ( .I1(n1356), .I2(n1295), .O(n1294) );
  INV_GATE U2364 ( .I1(n1294), .O(n10975) );
  AND_GATE U2365 ( .I1(n10984), .I2(n10955), .O(n1295) );
  OR_GATE U2366 ( .I1(n11849), .I2(n479), .O(n11851) );
  OR_GATE U2367 ( .I1(n3591), .I2(n3657), .O(n2969) );
  INV_GATE U2368 ( .I1(n1296), .O(n3964) );
  OR_GATE U2369 ( .I1(n1297), .I2(n2028), .O(n2037) );
  INV_GATE U2370 ( .I1(n14960), .O(n1298) );
  OR_GATE U2371 ( .I1(n1299), .I2(n8998), .O(n9001) );
  INV_GATE U2372 ( .I1(n8999), .O(n1299) );
  OR_GATE U2373 ( .I1(n7135), .I2(n631), .O(n7138) );
  OR_GATE U2374 ( .I1(n9093), .I2(n768), .O(n9096) );
  OR_GATE U2375 ( .I1(n10194), .I2(n10195), .O(n10198) );
  AND_GATE U2376 ( .I1(n11834), .I2(n11833), .O(n1300) );
  AND_GATE U2377 ( .I1(n9158), .I2(n9163), .O(n1301) );
  AND_GATE U2378 ( .I1(n1343), .I2(n6721), .O(n1302) );
  NOR_GATE U2379 ( .I1(n3712), .I2(n3711), .O(n1303) );
  AND3_GATE U2380 ( .I1(n3899), .I2(n3898), .I3(n3900), .O(n1304) );
  AND_GATE U2381 ( .I1(n1305), .I2(n14453), .O(n1308) );
  AND_GATE U2382 ( .I1(n14447), .I2(n14446), .O(n1305) );
  OR_GATE U2383 ( .I1(n10181), .I2(n857), .O(n10178) );
  OR_GATE U2384 ( .I1(n1306), .I2(n8965), .O(n8967) );
  INV_GATE U2385 ( .I1(n8966), .O(n1306) );
  AND3_GATE U2386 ( .I1(n1995), .I2(n1994), .I3(n1993), .O(n1307) );
  NOR_GATE U2387 ( .I1(n2686), .I2(n280), .O(n1309) );
  INV_GATE U2388 ( .I1(n1309), .O(n3045) );
  OR_GATE U2389 ( .I1(n3915), .I2(n1263), .O(n3918) );
  OR_GATE U2390 ( .I1(n6230), .I2(n6221), .O(n6238) );
  NOR_GATE U2391 ( .I1(n3901), .I2(n1304), .O(n1311) );
  OR4_GATE U2392 ( .I1(n1312), .I2(n2982), .I3(n3678), .I4(n3672), .O(n3677)
         );
  INV_GATE U2393 ( .I1(n3669), .O(n1312) );
  OR_GATE U2394 ( .I1(n20), .I2(n6543), .O(n6545) );
  NAND_GATE U2395 ( .I1(n9842), .I2(n1315), .O(n1313) );
  AND_GATE U2396 ( .I1(n1313), .I2(n1314), .O(n10654) );
  OR_GATE U2397 ( .I1(n10653), .I2(n567), .O(n1314) );
  AND_GATE U2398 ( .I1(n9841), .I2(n10164), .O(n1315) );
  NAND_GATE U2399 ( .I1(n14877), .I2(n1318), .O(n1316) );
  OR_GATE U2400 ( .I1(n425), .I2(n1342), .O(n1317) );
  OR_GATE U2401 ( .I1(n281), .I2(n14407), .O(n1319) );
  NAND_GATE U2402 ( .I1(n1332), .I2(n1322), .O(n1320) );
  AND_GATE U2403 ( .I1(n1320), .I2(n1321), .O(n5464) );
  OR_GATE U2404 ( .I1(n5455), .I2(n5454), .O(n1321) );
  AND_GATE U2405 ( .I1(n4782), .I2(n5462), .O(n1322) );
  AND_GATE U2406 ( .I1(n14861), .I2(n14860), .O(n1323) );
  AND_GATE U2407 ( .I1(n13244), .I2(n13243), .O(n1324) );
  AND_GATE U2408 ( .I1(n12392), .I2(n12391), .O(n1325) );
  AND3_GATE U2409 ( .I1(n11527), .I2(n11526), .I3(n11525), .O(n1326) );
  AND3_GATE U2410 ( .I1(n10660), .I2(n10659), .I3(n10658), .O(n1327) );
  AND_GATE U2411 ( .I1(n8090), .I2(n8089), .O(n1329) );
  AND_GATE U2412 ( .I1(n7231), .I2(n7230), .O(n1330) );
  AND_GATE U2413 ( .I1(n6573), .I2(n6571), .O(n1331) );
  AND_GATE U2414 ( .I1(n4777), .I2(n4778), .O(n1332) );
  NAND_GATE U2415 ( .I1(n13097), .I2(n1336), .O(n1334) );
  AND_GATE U2416 ( .I1(n1334), .I2(n1335), .O(n13234) );
  OR_GATE U2417 ( .I1(n13240), .I2(n13099), .O(n1335) );
  NAND_GATE U2418 ( .I1(n12195), .I2(n1339), .O(n1337) );
  AND_GATE U2419 ( .I1(n1337), .I2(n1338), .O(n12380) );
  OR_GATE U2420 ( .I1(n12388), .I2(n12198), .O(n1338) );
  AND_GATE U2421 ( .I1(n12196), .I2(n12199), .O(n1339) );
  AND_GATE U2422 ( .I1(n11058), .I2(n11057), .O(n1340) );
  AND_GATE U2423 ( .I1(n8421), .I2(n8420), .O(n1341) );
  INV_GATE U2424 ( .I1(n14914), .O(n1342) );
  AND3_GATE U2425 ( .I1(n6554), .I2(n6426), .I3(n6425), .O(n1343) );
  INV_GATE U2426 ( .I1(n1343), .O(n7365) );
  AND_GATE U2427 ( .I1(n7411), .I2(n7410), .O(n1344) );
  INV_GATE U2428 ( .I1(n1344), .O(n7693) );
  NAND_GATE U2429 ( .I1(n14893), .I2(n1271), .O(n14892) );
  NAND_GATE U2430 ( .I1(n7610), .I2(n1347), .O(n1345) );
  AND_GATE U2431 ( .I1(n1345), .I2(n1346), .O(n7612) );
  AND_GATE U2432 ( .I1(n7609), .I2(n7611), .O(n1347) );
  NAND_GATE U2433 ( .I1(n1348), .I2(n14379), .O(n14378) );
  NOR_GATE U2434 ( .I1(n14380), .I2(n14381), .O(n1348) );
  AND_GATE U2435 ( .I1(n306), .I2(n300), .O(n1349) );
  NAND_GATE U2436 ( .I1(n14833), .I2(n14989), .O(n1350) );
  NOR_GATE U2437 ( .I1(n5694), .I2(n5696), .O(n1351) );
  OR_GATE U2438 ( .I1(n1352), .I2(n5861), .O(n6507) );
  INV_GATE U2439 ( .I1(n5862), .O(n1352) );
  NOR_GATE U2440 ( .I1(n9860), .I2(n9853), .O(n1353) );
  AND_GATE U2441 ( .I1(n12751), .I2(n12752), .O(n1354) );
  NOR_GATE U2442 ( .I1(n7619), .I2(n7620), .O(n1355) );
  OR_GATE U2443 ( .I1(n11464), .I2(n11461), .O(n11837) );
  NOR_GATE U2444 ( .I1(n10982), .I2(n10983), .O(n1356) );
  NOR_GATE U2445 ( .I1(n281), .I2(n14407), .O(n1357) );
  AND3_GATE U2446 ( .I1(n7378), .I2(n6727), .I3(n6726), .O(n1358) );
  INV_GATE U2447 ( .I1(n1358), .O(n7387) );
  AND3_GATE U2448 ( .I1(n6687), .I2(n6686), .I3(n6685), .O(n1359) );
  INV_GATE U2449 ( .I1(n1359), .O(n7241) );
  AND3_GATE U2450 ( .I1(n8255), .I2(n7689), .I3(n7688), .O(n1360) );
  AND3_GATE U2451 ( .I1(n5705), .I2(n5449), .I3(n5713), .O(n1361) );
  INV_GATE U2452 ( .I1(n1361), .O(n5735) );
  AND_GATE U2453 ( .I1(n14538), .I2(n14537), .O(n1362) );
  INV_GATE U2454 ( .I1(n1362), .O(n15014) );
  AND_GATE U2455 ( .I1(n5518), .I2(n5522), .O(n1363) );
  INV_GATE U2456 ( .I1(B[1]), .O(n1364) );
  INV_GATE U2457 ( .I1(n1366), .O(n1365) );
  INV_GATE U2458 ( .I1(B[2]), .O(n1366) );
  INV_GATE U2459 ( .I1(B[3]), .O(n1367) );
  INV_GATE U2460 ( .I1(B[4]), .O(n1368) );
  INV_GATE U2461 ( .I1(B[5]), .O(n1369) );
  INV_GATE U2462 ( .I1(B[6]), .O(n1370) );
  INV_GATE U2463 ( .I1(B[7]), .O(n1371) );
  INV_GATE U2464 ( .I1(B[8]), .O(n1372) );
  INV_GATE U2465 ( .I1(B[9]), .O(n1373) );
  INV_GATE U2466 ( .I1(B[10]), .O(n1374) );
  INV_GATE U2467 ( .I1(B[11]), .O(n1375) );
  INV_GATE U2468 ( .I1(B[12]), .O(n1376) );
  INV_GATE U2469 ( .I1(B[13]), .O(n1377) );
  INV_GATE U2470 ( .I1(B[14]), .O(n1378) );
  INV_GATE U2471 ( .I1(n1380), .O(n1379) );
  INV_GATE U2472 ( .I1(B[15]), .O(n1380) );
  INV_GATE U2473 ( .I1(B[16]), .O(n1381) );
  INV_GATE U2474 ( .I1(n1383), .O(n1382) );
  INV_GATE U2475 ( .I1(B[17]), .O(n1383) );
  INV_GATE U2476 ( .I1(B[18]), .O(n1384) );
  INV_GATE U2477 ( .I1(B[19]), .O(n1385) );
  INV_GATE U2478 ( .I1(B[20]), .O(n1386) );
  INV_GATE U2479 ( .I1(B[21]), .O(n1387) );
  INV_GATE U2480 ( .I1(B[22]), .O(n1388) );
  INV_GATE U2481 ( .I1(B[23]), .O(n1389) );
  INV_GATE U2482 ( .I1(B[24]), .O(n1390) );
  INV_GATE U2483 ( .I1(B[25]), .O(n1391) );
  INV_GATE U2484 ( .I1(B[26]), .O(n1392) );
  INV_GATE U2485 ( .I1(B[27]), .O(n1393) );
  INV_GATE U2486 ( .I1(B[28]), .O(n1394) );
  INV_GATE U2487 ( .I1(B[29]), .O(n1395) );
  INV_GATE U2488 ( .I1(B[30]), .O(n1396) );
  INV_GATE U2489 ( .I1(B[31]), .O(n1397) );
  INV_GATE U2490 ( .I1(A[0]), .O(n1398) );
  INV_GATE U2491 ( .I1(A[1]), .O(n1399) );
  INV_GATE U2492 ( .I1(A[2]), .O(n1400) );
  INV_GATE U2493 ( .I1(A[3]), .O(n1401) );
  INV_GATE U2494 ( .I1(A[4]), .O(n1402) );
  INV_GATE U2495 ( .I1(A[5]), .O(n1403) );
  INV_GATE U2496 ( .I1(A[6]), .O(n1404) );
  INV_GATE U2497 ( .I1(A[7]), .O(n1405) );
  INV_GATE U2498 ( .I1(A[8]), .O(n1406) );
  INV_GATE U2499 ( .I1(A[9]), .O(n1407) );
  INV_GATE U2500 ( .I1(A[10]), .O(n1408) );
  INV_GATE U2501 ( .I1(A[11]), .O(n1409) );
  INV_GATE U2502 ( .I1(A[12]), .O(n1410) );
  INV_GATE U2503 ( .I1(A[13]), .O(n1411) );
  INV_GATE U2504 ( .I1(A[14]), .O(n1412) );
  INV_GATE U2505 ( .I1(A[15]), .O(n1413) );
  INV_GATE U2506 ( .I1(A[16]), .O(n1414) );
  INV_GATE U2507 ( .I1(A[17]), .O(n1415) );
  INV_GATE U2508 ( .I1(A[18]), .O(n1416) );
  INV_GATE U2509 ( .I1(A[19]), .O(n1417) );
  INV_GATE U2510 ( .I1(A[20]), .O(n1418) );
  INV_GATE U2511 ( .I1(A[21]), .O(n1419) );
  INV_GATE U2512 ( .I1(A[22]), .O(n1420) );
  INV_GATE U2513 ( .I1(A[23]), .O(n1421) );
  INV_GATE U2514 ( .I1(A[24]), .O(n1422) );
  INV_GATE U2515 ( .I1(A[25]), .O(n1423) );
  INV_GATE U2516 ( .I1(A[26]), .O(n1424) );
  INV_GATE U2517 ( .I1(A[27]), .O(n1425) );
  INV_GATE U2518 ( .I1(A[28]), .O(n1426) );
  INV_GATE U2519 ( .I1(A[29]), .O(n1427) );
  INV_GATE U2520 ( .I1(A[30]), .O(n1428) );
  INV_GATE U2521 ( .I1(A[31]), .O(n1429) );
  NAND_GATE U2522 ( .I1(n15379), .I2(n291), .O(n1431) );
  OR_GATE U2523 ( .I1(n291), .I2(n15379), .O(n1430) );
  NAND_GATE U2524 ( .I1(n1431), .I2(n1430), .O(PRODUCT[1]) );
  NAND3_GATE U2525 ( .I1(A[31]), .I2(A[30]), .I3(n1192), .O(n1518) );
  NAND3_GATE U2526 ( .I1(A[29]), .I2(A[30]), .I3(n1192), .O(n1515) );
  NAND3_GATE U2527 ( .I1(A[28]), .I2(A[29]), .I3(n1192), .O(n1512) );
  NAND3_GATE U2528 ( .I1(A[27]), .I2(A[28]), .I3(n1192), .O(n1509) );
  NAND3_GATE U2529 ( .I1(A[26]), .I2(A[27]), .I3(n1192), .O(n1506) );
  NAND3_GATE U2530 ( .I1(A[25]), .I2(A[26]), .I3(n1192), .O(n1503) );
  NAND3_GATE U2531 ( .I1(A[24]), .I2(A[25]), .I3(n1192), .O(n1500) );
  NAND3_GATE U2532 ( .I1(A[23]), .I2(A[24]), .I3(n1192), .O(n1497) );
  NAND3_GATE U2533 ( .I1(A[22]), .I2(A[23]), .I3(n1192), .O(n1494) );
  NAND3_GATE U2534 ( .I1(A[21]), .I2(A[22]), .I3(n1192), .O(n1491) );
  NAND3_GATE U2535 ( .I1(A[20]), .I2(A[21]), .I3(n1192), .O(n1488) );
  NAND3_GATE U2536 ( .I1(A[19]), .I2(A[20]), .I3(n1192), .O(n1485) );
  NAND3_GATE U2537 ( .I1(A[18]), .I2(A[19]), .I3(n1192), .O(n1482) );
  NAND3_GATE U2538 ( .I1(A[17]), .I2(A[18]), .I3(n1192), .O(n1479) );
  NAND3_GATE U2539 ( .I1(A[16]), .I2(A[17]), .I3(n1192), .O(n1476) );
  NAND3_GATE U2540 ( .I1(A[15]), .I2(A[16]), .I3(n1192), .O(n1473) );
  NAND3_GATE U2541 ( .I1(A[14]), .I2(A[15]), .I3(n1192), .O(n1470) );
  NAND3_GATE U2542 ( .I1(A[13]), .I2(A[14]), .I3(n1192), .O(n1467) );
  NAND3_GATE U2543 ( .I1(A[12]), .I2(A[13]), .I3(n1192), .O(n1464) );
  NAND3_GATE U2544 ( .I1(A[11]), .I2(A[12]), .I3(n1192), .O(n1461) );
  NAND3_GATE U2545 ( .I1(A[10]), .I2(A[11]), .I3(n1192), .O(n1458) );
  NAND3_GATE U2546 ( .I1(A[9]), .I2(A[10]), .I3(n1192), .O(n1455) );
  NAND3_GATE U2547 ( .I1(A[8]), .I2(A[9]), .I3(n1192), .O(n1452) );
  NAND3_GATE U2548 ( .I1(A[7]), .I2(A[8]), .I3(n1192), .O(n1449) );
  NAND3_GATE U2549 ( .I1(A[6]), .I2(A[7]), .I3(n1192), .O(n1446) );
  NAND3_GATE U2550 ( .I1(A[5]), .I2(A[6]), .I3(n1192), .O(n1443) );
  NAND3_GATE U2551 ( .I1(A[4]), .I2(A[5]), .I3(n1192), .O(n1440) );
  NAND3_GATE U2552 ( .I1(A[3]), .I2(A[4]), .I3(n1192), .O(n1437) );
  NAND3_GATE U2553 ( .I1(A[2]), .I2(A[3]), .I3(n1192), .O(n1434) );
  NAND_GATE U2554 ( .I1(n1192), .I2(n1196), .O(n1864) );
  NAND3_GATE U2555 ( .I1(A[2]), .I2(A[1]), .I3(n1192), .O(n1862) );
  NAND_GATE U2556 ( .I1(n1864), .I2(n1862), .O(n1857) );
  OR_GATE U2557 ( .I1(A[2]), .I2(A[3]), .O(n1432) );
  NAND_GATE U2558 ( .I1(n1857), .I2(n1432), .O(n1433) );
  NAND_GATE U2559 ( .I1(n1434), .I2(n1433), .O(n1845) );
  OR_GATE U2560 ( .I1(A[3]), .I2(A[4]), .O(n1435) );
  NAND_GATE U2561 ( .I1(n1845), .I2(n1435), .O(n1436) );
  NAND_GATE U2562 ( .I1(n1437), .I2(n1436), .O(n1833) );
  OR_GATE U2563 ( .I1(A[4]), .I2(A[5]), .O(n1438) );
  NAND_GATE U2564 ( .I1(n1833), .I2(n1438), .O(n1439) );
  NAND_GATE U2565 ( .I1(n1440), .I2(n1439), .O(n1821) );
  OR_GATE U2566 ( .I1(A[5]), .I2(A[6]), .O(n1441) );
  NAND_GATE U2567 ( .I1(n1821), .I2(n1441), .O(n1442) );
  NAND_GATE U2568 ( .I1(n1443), .I2(n1442), .O(n1809) );
  OR_GATE U2569 ( .I1(A[6]), .I2(A[7]), .O(n1444) );
  NAND_GATE U2570 ( .I1(n1809), .I2(n1444), .O(n1445) );
  NAND_GATE U2571 ( .I1(n1446), .I2(n1445), .O(n1797) );
  OR_GATE U2572 ( .I1(A[7]), .I2(A[8]), .O(n1447) );
  NAND_GATE U2573 ( .I1(n1797), .I2(n1447), .O(n1448) );
  NAND_GATE U2574 ( .I1(n1449), .I2(n1448), .O(n1785) );
  OR_GATE U2575 ( .I1(A[8]), .I2(A[9]), .O(n1450) );
  NAND_GATE U2576 ( .I1(n1785), .I2(n1450), .O(n1451) );
  NAND_GATE U2577 ( .I1(n1452), .I2(n1451), .O(n1773) );
  OR_GATE U2578 ( .I1(A[9]), .I2(A[10]), .O(n1453) );
  NAND_GATE U2579 ( .I1(n1773), .I2(n1453), .O(n1454) );
  NAND_GATE U2580 ( .I1(n1455), .I2(n1454), .O(n1761) );
  OR_GATE U2581 ( .I1(A[10]), .I2(A[11]), .O(n1456) );
  NAND_GATE U2582 ( .I1(n1761), .I2(n1456), .O(n1457) );
  NAND_GATE U2583 ( .I1(n1458), .I2(n1457), .O(n1749) );
  OR_GATE U2584 ( .I1(A[11]), .I2(A[12]), .O(n1459) );
  NAND_GATE U2585 ( .I1(n1749), .I2(n1459), .O(n1460) );
  NAND_GATE U2586 ( .I1(n1461), .I2(n1460), .O(n1737) );
  OR_GATE U2587 ( .I1(A[12]), .I2(A[13]), .O(n1462) );
  NAND_GATE U2588 ( .I1(n1737), .I2(n1462), .O(n1463) );
  NAND_GATE U2589 ( .I1(n1464), .I2(n1463), .O(n1725) );
  OR_GATE U2590 ( .I1(A[13]), .I2(A[14]), .O(n1465) );
  NAND_GATE U2591 ( .I1(n1725), .I2(n1465), .O(n1466) );
  NAND_GATE U2592 ( .I1(n1467), .I2(n1466), .O(n1713) );
  OR_GATE U2593 ( .I1(A[14]), .I2(A[15]), .O(n1468) );
  NAND_GATE U2594 ( .I1(n1713), .I2(n1468), .O(n1469) );
  NAND_GATE U2595 ( .I1(n1470), .I2(n1469), .O(n1701) );
  OR_GATE U2596 ( .I1(A[15]), .I2(A[16]), .O(n1471) );
  NAND_GATE U2597 ( .I1(n1701), .I2(n1471), .O(n1472) );
  NAND_GATE U2598 ( .I1(n1473), .I2(n1472), .O(n1689) );
  OR_GATE U2599 ( .I1(A[16]), .I2(A[17]), .O(n1474) );
  NAND_GATE U2600 ( .I1(n1689), .I2(n1474), .O(n1475) );
  NAND_GATE U2601 ( .I1(n1476), .I2(n1475), .O(n1677) );
  OR_GATE U2602 ( .I1(A[17]), .I2(A[18]), .O(n1477) );
  NAND_GATE U2603 ( .I1(n1677), .I2(n1477), .O(n1478) );
  NAND_GATE U2604 ( .I1(n1479), .I2(n1478), .O(n1665) );
  OR_GATE U2605 ( .I1(A[18]), .I2(A[19]), .O(n1480) );
  NAND_GATE U2606 ( .I1(n1665), .I2(n1480), .O(n1481) );
  NAND_GATE U2607 ( .I1(n1482), .I2(n1481), .O(n1653) );
  OR_GATE U2608 ( .I1(A[19]), .I2(A[20]), .O(n1483) );
  NAND_GATE U2609 ( .I1(n1653), .I2(n1483), .O(n1484) );
  NAND_GATE U2610 ( .I1(n1485), .I2(n1484), .O(n1641) );
  OR_GATE U2611 ( .I1(A[20]), .I2(A[21]), .O(n1486) );
  NAND_GATE U2612 ( .I1(n1641), .I2(n1486), .O(n1487) );
  NAND_GATE U2613 ( .I1(n1488), .I2(n1487), .O(n1629) );
  OR_GATE U2614 ( .I1(A[21]), .I2(A[22]), .O(n1489) );
  NAND_GATE U2615 ( .I1(n1629), .I2(n1489), .O(n1490) );
  NAND_GATE U2616 ( .I1(n1491), .I2(n1490), .O(n1617) );
  OR_GATE U2617 ( .I1(A[22]), .I2(A[23]), .O(n1492) );
  NAND_GATE U2618 ( .I1(n1617), .I2(n1492), .O(n1493) );
  NAND_GATE U2619 ( .I1(n1494), .I2(n1493), .O(n1605) );
  OR_GATE U2620 ( .I1(A[23]), .I2(A[24]), .O(n1495) );
  NAND_GATE U2621 ( .I1(n1605), .I2(n1495), .O(n1496) );
  NAND_GATE U2622 ( .I1(n1497), .I2(n1496), .O(n1593) );
  OR_GATE U2623 ( .I1(A[24]), .I2(A[25]), .O(n1498) );
  NAND_GATE U2624 ( .I1(n1593), .I2(n1498), .O(n1499) );
  NAND_GATE U2625 ( .I1(n1500), .I2(n1499), .O(n1581) );
  OR_GATE U2626 ( .I1(A[25]), .I2(A[26]), .O(n1501) );
  NAND_GATE U2627 ( .I1(n1581), .I2(n1501), .O(n1502) );
  NAND_GATE U2628 ( .I1(n1503), .I2(n1502), .O(n1569) );
  OR_GATE U2629 ( .I1(A[26]), .I2(A[27]), .O(n1504) );
  NAND_GATE U2630 ( .I1(n1569), .I2(n1504), .O(n1505) );
  NAND_GATE U2631 ( .I1(n1506), .I2(n1505), .O(n1557) );
  OR_GATE U2632 ( .I1(A[27]), .I2(A[28]), .O(n1507) );
  NAND_GATE U2633 ( .I1(n1557), .I2(n1507), .O(n1508) );
  NAND_GATE U2634 ( .I1(n1509), .I2(n1508), .O(n1940) );
  OR_GATE U2635 ( .I1(A[28]), .I2(A[29]), .O(n1510) );
  NAND_GATE U2636 ( .I1(n1940), .I2(n1510), .O(n1511) );
  NAND_GATE U2637 ( .I1(n1512), .I2(n1511), .O(n1545) );
  OR_GATE U2638 ( .I1(A[29]), .I2(A[30]), .O(n1513) );
  NAND_GATE U2639 ( .I1(n1545), .I2(n1513), .O(n1514) );
  NAND_GATE U2640 ( .I1(n1515), .I2(n1514), .O(n1533) );
  OR_GATE U2641 ( .I1(A[31]), .I2(A[30]), .O(n1516) );
  NAND_GATE U2642 ( .I1(n1533), .I2(n1516), .O(n1517) );
  NAND_GATE U2643 ( .I1(n1518), .I2(n1517), .O(n15305) );
  INV_GATE U2644 ( .I1(n15305), .O(n1519) );
  NAND_GATE U2645 ( .I1(A[31]), .I2(B[31]), .O(n1520) );
  NAND_GATE U2646 ( .I1(n1519), .I2(n1520), .O(n1523) );
  INV_GATE U2647 ( .I1(n1520), .O(n1521) );
  NAND_GATE U2648 ( .I1(n15305), .I2(n1521), .O(n1522) );
  AND_GATE U2649 ( .I1(n1523), .I2(n1522), .O(\A1[60] ) );
  INV_GATE U2650 ( .I1(n1533), .O(n1530) );
  NAND_GATE U2651 ( .I1(n1397), .I2(B[30]), .O(n1930) );
  NAND_GATE U2652 ( .I1(n1428), .I2(B[30]), .O(n1524) );
  NAND_GATE U2653 ( .I1(n1930), .I2(n1524), .O(n1525) );
  NAND_GATE U2654 ( .I1(A[31]), .I2(n1525), .O(n1529) );
  NAND_GATE U2655 ( .I1(n1429), .I2(B[31]), .O(n1526) );
  NAND_GATE U2656 ( .I1(n1933), .I2(n1526), .O(n1527) );
  NAND_GATE U2657 ( .I1(A[30]), .I2(n1527), .O(n1528) );
  NAND_GATE U2658 ( .I1(n1529), .I2(n1528), .O(n1531) );
  NAND_GATE U2659 ( .I1(n1530), .I2(n1531), .O(n1535) );
  INV_GATE U2660 ( .I1(n1531), .O(n1532) );
  NAND_GATE U2661 ( .I1(n1533), .I2(n1532), .O(n1534) );
  NAND_GATE U2662 ( .I1(n1535), .I2(n1534), .O(n15307) );
  INV_GATE U2663 ( .I1(n15307), .O(n1947) );
  NAND_GATE U2664 ( .I1(B[29]), .I2(A[31]), .O(n2448) );
  INV_GATE U2665 ( .I1(n2448), .O(n2441) );
  INV_GATE U2666 ( .I1(n1545), .O(n1542) );
  NAND_GATE U2667 ( .I1(n1427), .I2(B[30]), .O(n1536) );
  NAND_GATE U2668 ( .I1(n1930), .I2(n1536), .O(n1537) );
  NAND_GATE U2669 ( .I1(A[30]), .I2(n1537), .O(n1541) );
  NAND_GATE U2670 ( .I1(n1428), .I2(B[31]), .O(n1538) );
  NAND_GATE U2671 ( .I1(n1933), .I2(n1538), .O(n1539) );
  NAND_GATE U2672 ( .I1(A[29]), .I2(n1539), .O(n1540) );
  NAND_GATE U2673 ( .I1(n1541), .I2(n1540), .O(n1543) );
  NAND_GATE U2674 ( .I1(n1542), .I2(n1543), .O(n1547) );
  INV_GATE U2675 ( .I1(n1543), .O(n1544) );
  NAND_GATE U2676 ( .I1(n1545), .I2(n1544), .O(n1546) );
  NAND_GATE U2677 ( .I1(n1547), .I2(n1546), .O(n2443) );
  NAND_GATE U2678 ( .I1(n2441), .I2(n2443), .O(n2438) );
  NAND_GATE U2679 ( .I1(B[29]), .I2(A[30]), .O(n2431) );
  INV_GATE U2680 ( .I1(n2431), .O(n2424) );
  NAND_GATE U2681 ( .I1(B[29]), .I2(A[29]), .O(n2414) );
  INV_GATE U2682 ( .I1(n2414), .O(n2407) );
  INV_GATE U2683 ( .I1(n1557), .O(n1554) );
  NAND_GATE U2684 ( .I1(n1425), .I2(B[30]), .O(n1548) );
  NAND_GATE U2685 ( .I1(n1930), .I2(n1548), .O(n1549) );
  NAND_GATE U2686 ( .I1(A[28]), .I2(n1549), .O(n1553) );
  NAND_GATE U2687 ( .I1(n1426), .I2(B[31]), .O(n1550) );
  NAND_GATE U2688 ( .I1(n1933), .I2(n1550), .O(n1551) );
  NAND_GATE U2689 ( .I1(A[27]), .I2(n1551), .O(n1552) );
  NAND_GATE U2690 ( .I1(n1553), .I2(n1552), .O(n1555) );
  NAND_GATE U2691 ( .I1(n1554), .I2(n1555), .O(n1559) );
  INV_GATE U2692 ( .I1(n1555), .O(n1556) );
  NAND_GATE U2693 ( .I1(n1557), .I2(n1556), .O(n1558) );
  NAND_GATE U2694 ( .I1(n1559), .I2(n1558), .O(n2409) );
  NAND_GATE U2695 ( .I1(n2407), .I2(n2409), .O(n2404) );
  NAND_GATE U2696 ( .I1(B[29]), .I2(A[28]), .O(n1961) );
  INV_GATE U2697 ( .I1(n1961), .O(n1954) );
  INV_GATE U2698 ( .I1(n1569), .O(n1566) );
  NAND_GATE U2699 ( .I1(n1424), .I2(B[30]), .O(n1560) );
  NAND_GATE U2700 ( .I1(n1930), .I2(n1560), .O(n1561) );
  NAND_GATE U2701 ( .I1(A[27]), .I2(n1561), .O(n1565) );
  NAND_GATE U2702 ( .I1(n1425), .I2(B[31]), .O(n1562) );
  NAND_GATE U2703 ( .I1(n1933), .I2(n1562), .O(n1563) );
  NAND_GATE U2704 ( .I1(A[26]), .I2(n1563), .O(n1564) );
  NAND_GATE U2705 ( .I1(n1565), .I2(n1564), .O(n1567) );
  NAND_GATE U2706 ( .I1(n1566), .I2(n1567), .O(n1571) );
  INV_GATE U2707 ( .I1(n1567), .O(n1568) );
  NAND_GATE U2708 ( .I1(n1569), .I2(n1568), .O(n1570) );
  NAND_GATE U2709 ( .I1(n1571), .I2(n1570), .O(n1956) );
  NAND_GATE U2710 ( .I1(n1954), .I2(n1956), .O(n1951) );
  NAND_GATE U2711 ( .I1(B[29]), .I2(A[27]), .O(n2395) );
  INV_GATE U2712 ( .I1(n2395), .O(n2388) );
  INV_GATE U2713 ( .I1(n1581), .O(n1578) );
  NAND_GATE U2714 ( .I1(n1423), .I2(B[30]), .O(n1572) );
  NAND_GATE U2715 ( .I1(n1930), .I2(n1572), .O(n1573) );
  NAND_GATE U2716 ( .I1(A[26]), .I2(n1573), .O(n1577) );
  NAND_GATE U2717 ( .I1(n1424), .I2(B[31]), .O(n1574) );
  NAND_GATE U2718 ( .I1(n1933), .I2(n1574), .O(n1575) );
  NAND_GATE U2719 ( .I1(A[25]), .I2(n1575), .O(n1576) );
  NAND_GATE U2720 ( .I1(n1577), .I2(n1576), .O(n1579) );
  NAND_GATE U2721 ( .I1(n1578), .I2(n1579), .O(n1583) );
  INV_GATE U2722 ( .I1(n1579), .O(n1580) );
  NAND_GATE U2723 ( .I1(n1581), .I2(n1580), .O(n1582) );
  NAND_GATE U2724 ( .I1(n1583), .I2(n1582), .O(n2390) );
  NAND_GATE U2725 ( .I1(n2388), .I2(n2390), .O(n2385) );
  NAND_GATE U2726 ( .I1(B[29]), .I2(A[26]), .O(n2378) );
  INV_GATE U2727 ( .I1(n2378), .O(n2371) );
  INV_GATE U2728 ( .I1(n1593), .O(n1590) );
  NAND_GATE U2729 ( .I1(n1422), .I2(B[30]), .O(n1584) );
  NAND_GATE U2730 ( .I1(n1930), .I2(n1584), .O(n1585) );
  NAND_GATE U2731 ( .I1(A[25]), .I2(n1585), .O(n1589) );
  NAND_GATE U2732 ( .I1(n1423), .I2(B[31]), .O(n1586) );
  NAND_GATE U2733 ( .I1(n1933), .I2(n1586), .O(n1587) );
  NAND_GATE U2734 ( .I1(A[24]), .I2(n1587), .O(n1588) );
  NAND_GATE U2735 ( .I1(n1589), .I2(n1588), .O(n1591) );
  NAND_GATE U2736 ( .I1(n1590), .I2(n1591), .O(n1595) );
  INV_GATE U2737 ( .I1(n1591), .O(n1592) );
  NAND_GATE U2738 ( .I1(n1593), .I2(n1592), .O(n1594) );
  NAND_GATE U2739 ( .I1(n1595), .I2(n1594), .O(n2373) );
  NAND_GATE U2740 ( .I1(n2371), .I2(n2373), .O(n2368) );
  NAND_GATE U2741 ( .I1(B[29]), .I2(A[25]), .O(n2361) );
  INV_GATE U2742 ( .I1(n2361), .O(n2354) );
  INV_GATE U2743 ( .I1(n1605), .O(n1602) );
  NAND_GATE U2744 ( .I1(n1421), .I2(B[30]), .O(n1596) );
  NAND_GATE U2745 ( .I1(n1930), .I2(n1596), .O(n1597) );
  NAND_GATE U2746 ( .I1(A[24]), .I2(n1597), .O(n1601) );
  NAND_GATE U2747 ( .I1(n1422), .I2(B[31]), .O(n1598) );
  NAND_GATE U2748 ( .I1(n1933), .I2(n1598), .O(n1599) );
  NAND_GATE U2749 ( .I1(A[23]), .I2(n1599), .O(n1600) );
  NAND_GATE U2750 ( .I1(n1601), .I2(n1600), .O(n1603) );
  NAND_GATE U2751 ( .I1(n1602), .I2(n1603), .O(n1607) );
  INV_GATE U2752 ( .I1(n1603), .O(n1604) );
  NAND_GATE U2753 ( .I1(n1605), .I2(n1604), .O(n1606) );
  NAND_GATE U2754 ( .I1(n1607), .I2(n1606), .O(n2356) );
  NAND_GATE U2755 ( .I1(n2354), .I2(n2356), .O(n2351) );
  NAND_GATE U2756 ( .I1(B[29]), .I2(A[24]), .O(n2344) );
  INV_GATE U2757 ( .I1(n2344), .O(n2337) );
  INV_GATE U2758 ( .I1(n1617), .O(n1614) );
  NAND_GATE U2759 ( .I1(n1420), .I2(B[30]), .O(n1608) );
  NAND_GATE U2760 ( .I1(n1930), .I2(n1608), .O(n1609) );
  NAND_GATE U2761 ( .I1(A[23]), .I2(n1609), .O(n1613) );
  NAND_GATE U2762 ( .I1(n1421), .I2(B[31]), .O(n1610) );
  NAND_GATE U2763 ( .I1(n1933), .I2(n1610), .O(n1611) );
  NAND_GATE U2764 ( .I1(A[22]), .I2(n1611), .O(n1612) );
  NAND_GATE U2765 ( .I1(n1613), .I2(n1612), .O(n1615) );
  NAND_GATE U2766 ( .I1(n1614), .I2(n1615), .O(n1619) );
  INV_GATE U2767 ( .I1(n1615), .O(n1616) );
  NAND_GATE U2768 ( .I1(n1617), .I2(n1616), .O(n1618) );
  NAND_GATE U2769 ( .I1(n1619), .I2(n1618), .O(n2339) );
  NAND_GATE U2770 ( .I1(n2337), .I2(n2339), .O(n2334) );
  NAND_GATE U2771 ( .I1(B[29]), .I2(A[23]), .O(n2327) );
  INV_GATE U2772 ( .I1(n2327), .O(n2320) );
  INV_GATE U2773 ( .I1(n1629), .O(n1626) );
  NAND_GATE U2774 ( .I1(n1419), .I2(B[30]), .O(n1620) );
  NAND_GATE U2775 ( .I1(n1930), .I2(n1620), .O(n1621) );
  NAND_GATE U2776 ( .I1(A[22]), .I2(n1621), .O(n1625) );
  NAND_GATE U2777 ( .I1(n1420), .I2(B[31]), .O(n1622) );
  NAND_GATE U2778 ( .I1(n1933), .I2(n1622), .O(n1623) );
  NAND_GATE U2779 ( .I1(A[21]), .I2(n1623), .O(n1624) );
  NAND_GATE U2780 ( .I1(n1625), .I2(n1624), .O(n1627) );
  NAND_GATE U2781 ( .I1(n1626), .I2(n1627), .O(n1631) );
  INV_GATE U2782 ( .I1(n1627), .O(n1628) );
  NAND_GATE U2783 ( .I1(n1629), .I2(n1628), .O(n1630) );
  NAND_GATE U2784 ( .I1(n1631), .I2(n1630), .O(n2322) );
  NAND_GATE U2785 ( .I1(n2320), .I2(n2322), .O(n2317) );
  NAND_GATE U2786 ( .I1(B[29]), .I2(A[22]), .O(n2310) );
  INV_GATE U2787 ( .I1(n2310), .O(n2303) );
  INV_GATE U2788 ( .I1(n1641), .O(n1638) );
  NAND_GATE U2789 ( .I1(n1418), .I2(B[30]), .O(n1632) );
  NAND_GATE U2790 ( .I1(n1930), .I2(n1632), .O(n1633) );
  NAND_GATE U2791 ( .I1(A[21]), .I2(n1633), .O(n1637) );
  NAND_GATE U2792 ( .I1(n1419), .I2(B[31]), .O(n1634) );
  NAND_GATE U2793 ( .I1(n1933), .I2(n1634), .O(n1635) );
  NAND_GATE U2794 ( .I1(A[20]), .I2(n1635), .O(n1636) );
  NAND_GATE U2795 ( .I1(n1637), .I2(n1636), .O(n1639) );
  NAND_GATE U2796 ( .I1(n1638), .I2(n1639), .O(n1643) );
  INV_GATE U2797 ( .I1(n1639), .O(n1640) );
  NAND_GATE U2798 ( .I1(n1641), .I2(n1640), .O(n1642) );
  NAND_GATE U2799 ( .I1(n1643), .I2(n1642), .O(n2305) );
  NAND_GATE U2800 ( .I1(n2303), .I2(n2305), .O(n2300) );
  NAND_GATE U2801 ( .I1(B[29]), .I2(A[21]), .O(n2293) );
  INV_GATE U2802 ( .I1(n2293), .O(n2286) );
  INV_GATE U2803 ( .I1(n1653), .O(n1650) );
  NAND_GATE U2804 ( .I1(n1417), .I2(B[30]), .O(n1644) );
  NAND_GATE U2805 ( .I1(n1930), .I2(n1644), .O(n1645) );
  NAND_GATE U2806 ( .I1(A[20]), .I2(n1645), .O(n1649) );
  NAND_GATE U2807 ( .I1(n1418), .I2(B[31]), .O(n1646) );
  NAND_GATE U2808 ( .I1(n1933), .I2(n1646), .O(n1647) );
  NAND_GATE U2809 ( .I1(A[19]), .I2(n1647), .O(n1648) );
  NAND_GATE U2810 ( .I1(n1649), .I2(n1648), .O(n1651) );
  NAND_GATE U2811 ( .I1(n1650), .I2(n1651), .O(n1655) );
  INV_GATE U2812 ( .I1(n1651), .O(n1652) );
  NAND_GATE U2813 ( .I1(n1653), .I2(n1652), .O(n1654) );
  NAND_GATE U2814 ( .I1(n1655), .I2(n1654), .O(n2288) );
  NAND_GATE U2815 ( .I1(n2286), .I2(n2288), .O(n2283) );
  NAND_GATE U2816 ( .I1(B[29]), .I2(A[20]), .O(n2276) );
  INV_GATE U2817 ( .I1(n2276), .O(n2269) );
  INV_GATE U2818 ( .I1(n1665), .O(n1662) );
  NAND_GATE U2819 ( .I1(n1416), .I2(B[30]), .O(n1656) );
  NAND_GATE U2820 ( .I1(n1930), .I2(n1656), .O(n1657) );
  NAND_GATE U2821 ( .I1(A[19]), .I2(n1657), .O(n1661) );
  NAND_GATE U2822 ( .I1(n1417), .I2(B[31]), .O(n1658) );
  NAND_GATE U2823 ( .I1(n1933), .I2(n1658), .O(n1659) );
  NAND_GATE U2824 ( .I1(A[18]), .I2(n1659), .O(n1660) );
  NAND_GATE U2825 ( .I1(n1661), .I2(n1660), .O(n1663) );
  NAND_GATE U2826 ( .I1(n1662), .I2(n1663), .O(n1667) );
  INV_GATE U2827 ( .I1(n1663), .O(n1664) );
  NAND_GATE U2828 ( .I1(n1665), .I2(n1664), .O(n1666) );
  NAND_GATE U2829 ( .I1(n1667), .I2(n1666), .O(n2271) );
  NAND_GATE U2830 ( .I1(n2269), .I2(n2271), .O(n2266) );
  NAND_GATE U2831 ( .I1(B[29]), .I2(A[19]), .O(n2260) );
  INV_GATE U2832 ( .I1(n2260), .O(n2253) );
  INV_GATE U2833 ( .I1(n1677), .O(n1674) );
  NAND_GATE U2834 ( .I1(n1415), .I2(B[30]), .O(n1668) );
  NAND_GATE U2835 ( .I1(n1930), .I2(n1668), .O(n1669) );
  NAND_GATE U2836 ( .I1(A[18]), .I2(n1669), .O(n1673) );
  NAND_GATE U2837 ( .I1(n1416), .I2(B[31]), .O(n1670) );
  NAND_GATE U2838 ( .I1(n1933), .I2(n1670), .O(n1671) );
  NAND_GATE U2839 ( .I1(A[17]), .I2(n1671), .O(n1672) );
  NAND_GATE U2840 ( .I1(n1673), .I2(n1672), .O(n1675) );
  NAND_GATE U2841 ( .I1(n1674), .I2(n1675), .O(n1679) );
  INV_GATE U2842 ( .I1(n1675), .O(n1676) );
  NAND_GATE U2843 ( .I1(n1677), .I2(n1676), .O(n1678) );
  NAND_GATE U2844 ( .I1(n1679), .I2(n1678), .O(n2255) );
  NAND_GATE U2845 ( .I1(n2253), .I2(n2255), .O(n2250) );
  NAND_GATE U2846 ( .I1(B[29]), .I2(A[18]), .O(n2244) );
  INV_GATE U2847 ( .I1(n2244), .O(n2237) );
  INV_GATE U2848 ( .I1(n1689), .O(n1686) );
  NAND_GATE U2849 ( .I1(n1414), .I2(B[30]), .O(n1680) );
  NAND_GATE U2850 ( .I1(n1930), .I2(n1680), .O(n1681) );
  NAND_GATE U2851 ( .I1(A[17]), .I2(n1681), .O(n1685) );
  NAND_GATE U2852 ( .I1(n1415), .I2(B[31]), .O(n1682) );
  NAND_GATE U2853 ( .I1(n1933), .I2(n1682), .O(n1683) );
  NAND_GATE U2854 ( .I1(A[16]), .I2(n1683), .O(n1684) );
  NAND_GATE U2855 ( .I1(n1685), .I2(n1684), .O(n1687) );
  NAND_GATE U2856 ( .I1(n1686), .I2(n1687), .O(n1691) );
  INV_GATE U2857 ( .I1(n1687), .O(n1688) );
  NAND_GATE U2858 ( .I1(n1689), .I2(n1688), .O(n1690) );
  NAND_GATE U2859 ( .I1(n1691), .I2(n1690), .O(n2239) );
  NAND_GATE U2860 ( .I1(n2237), .I2(n2239), .O(n2234) );
  NAND_GATE U2861 ( .I1(B[29]), .I2(A[17]), .O(n2228) );
  INV_GATE U2862 ( .I1(n2228), .O(n2221) );
  INV_GATE U2863 ( .I1(n1701), .O(n1698) );
  NAND_GATE U2864 ( .I1(n1413), .I2(B[30]), .O(n1692) );
  NAND_GATE U2865 ( .I1(n1930), .I2(n1692), .O(n1693) );
  NAND_GATE U2866 ( .I1(A[16]), .I2(n1693), .O(n1697) );
  NAND_GATE U2867 ( .I1(n1414), .I2(B[31]), .O(n1694) );
  NAND_GATE U2868 ( .I1(n1933), .I2(n1694), .O(n1695) );
  NAND_GATE U2869 ( .I1(A[15]), .I2(n1695), .O(n1696) );
  NAND_GATE U2870 ( .I1(n1697), .I2(n1696), .O(n1699) );
  NAND_GATE U2871 ( .I1(n1698), .I2(n1699), .O(n1703) );
  INV_GATE U2872 ( .I1(n1699), .O(n1700) );
  NAND_GATE U2873 ( .I1(n1701), .I2(n1700), .O(n1702) );
  NAND_GATE U2874 ( .I1(n1703), .I2(n1702), .O(n2223) );
  NAND_GATE U2875 ( .I1(n2221), .I2(n2223), .O(n2218) );
  NAND_GATE U2876 ( .I1(B[29]), .I2(A[16]), .O(n2211) );
  INV_GATE U2877 ( .I1(n2211), .O(n2204) );
  INV_GATE U2878 ( .I1(n1713), .O(n1710) );
  NAND_GATE U2879 ( .I1(n1412), .I2(B[30]), .O(n1704) );
  NAND_GATE U2880 ( .I1(n1930), .I2(n1704), .O(n1705) );
  NAND_GATE U2881 ( .I1(A[15]), .I2(n1705), .O(n1709) );
  NAND_GATE U2882 ( .I1(n1413), .I2(B[31]), .O(n1706) );
  NAND_GATE U2883 ( .I1(n1933), .I2(n1706), .O(n1707) );
  NAND_GATE U2884 ( .I1(A[14]), .I2(n1707), .O(n1708) );
  NAND_GATE U2885 ( .I1(n1709), .I2(n1708), .O(n1711) );
  NAND_GATE U2886 ( .I1(n1710), .I2(n1711), .O(n1715) );
  INV_GATE U2887 ( .I1(n1711), .O(n1712) );
  NAND_GATE U2888 ( .I1(n1713), .I2(n1712), .O(n1714) );
  NAND_GATE U2889 ( .I1(n1715), .I2(n1714), .O(n2206) );
  NAND_GATE U2890 ( .I1(n2204), .I2(n2206), .O(n2201) );
  NAND_GATE U2891 ( .I1(B[29]), .I2(A[15]), .O(n2194) );
  INV_GATE U2892 ( .I1(n2194), .O(n2187) );
  INV_GATE U2893 ( .I1(n1725), .O(n1722) );
  NAND_GATE U2894 ( .I1(n1411), .I2(B[30]), .O(n1716) );
  NAND_GATE U2895 ( .I1(n1930), .I2(n1716), .O(n1717) );
  NAND_GATE U2896 ( .I1(A[14]), .I2(n1717), .O(n1721) );
  NAND_GATE U2897 ( .I1(n1412), .I2(B[31]), .O(n1718) );
  NAND_GATE U2898 ( .I1(n1933), .I2(n1718), .O(n1719) );
  NAND_GATE U2899 ( .I1(A[13]), .I2(n1719), .O(n1720) );
  NAND_GATE U2900 ( .I1(n1721), .I2(n1720), .O(n1723) );
  NAND_GATE U2901 ( .I1(n1722), .I2(n1723), .O(n1727) );
  INV_GATE U2902 ( .I1(n1723), .O(n1724) );
  NAND_GATE U2903 ( .I1(n1725), .I2(n1724), .O(n1726) );
  NAND_GATE U2904 ( .I1(n1727), .I2(n1726), .O(n2189) );
  NAND_GATE U2905 ( .I1(n2187), .I2(n2189), .O(n2184) );
  NAND_GATE U2906 ( .I1(B[29]), .I2(A[14]), .O(n2177) );
  INV_GATE U2907 ( .I1(n2177), .O(n2170) );
  INV_GATE U2908 ( .I1(n1737), .O(n1734) );
  NAND_GATE U2909 ( .I1(n1410), .I2(B[30]), .O(n1728) );
  NAND_GATE U2910 ( .I1(n1930), .I2(n1728), .O(n1729) );
  NAND_GATE U2911 ( .I1(A[13]), .I2(n1729), .O(n1733) );
  NAND_GATE U2912 ( .I1(n1411), .I2(B[31]), .O(n1730) );
  NAND_GATE U2913 ( .I1(n1933), .I2(n1730), .O(n1731) );
  NAND_GATE U2914 ( .I1(A[12]), .I2(n1731), .O(n1732) );
  NAND_GATE U2915 ( .I1(n1733), .I2(n1732), .O(n1735) );
  NAND_GATE U2916 ( .I1(n1734), .I2(n1735), .O(n1739) );
  INV_GATE U2917 ( .I1(n1735), .O(n1736) );
  NAND_GATE U2918 ( .I1(n1737), .I2(n1736), .O(n1738) );
  NAND_GATE U2919 ( .I1(n1739), .I2(n1738), .O(n2172) );
  NAND_GATE U2920 ( .I1(n2170), .I2(n2172), .O(n2167) );
  NAND_GATE U2921 ( .I1(B[29]), .I2(A[13]), .O(n2160) );
  INV_GATE U2922 ( .I1(n2160), .O(n2153) );
  INV_GATE U2923 ( .I1(n1749), .O(n1746) );
  NAND_GATE U2924 ( .I1(n1409), .I2(B[30]), .O(n1740) );
  NAND_GATE U2925 ( .I1(n1930), .I2(n1740), .O(n1741) );
  NAND_GATE U2926 ( .I1(A[12]), .I2(n1741), .O(n1745) );
  NAND_GATE U2927 ( .I1(n1410), .I2(B[31]), .O(n1742) );
  NAND_GATE U2928 ( .I1(n1933), .I2(n1742), .O(n1743) );
  NAND_GATE U2929 ( .I1(A[11]), .I2(n1743), .O(n1744) );
  NAND_GATE U2930 ( .I1(n1745), .I2(n1744), .O(n1747) );
  NAND_GATE U2931 ( .I1(n1746), .I2(n1747), .O(n1751) );
  INV_GATE U2932 ( .I1(n1747), .O(n1748) );
  NAND_GATE U2933 ( .I1(n1749), .I2(n1748), .O(n1750) );
  NAND_GATE U2934 ( .I1(n1751), .I2(n1750), .O(n2155) );
  NAND_GATE U2935 ( .I1(n2153), .I2(n2155), .O(n2150) );
  NAND_GATE U2936 ( .I1(B[29]), .I2(A[12]), .O(n2143) );
  INV_GATE U2937 ( .I1(n2143), .O(n2136) );
  INV_GATE U2938 ( .I1(n1761), .O(n1758) );
  NAND_GATE U2939 ( .I1(n1408), .I2(B[30]), .O(n1752) );
  NAND_GATE U2940 ( .I1(n1930), .I2(n1752), .O(n1753) );
  NAND_GATE U2941 ( .I1(A[11]), .I2(n1753), .O(n1757) );
  NAND_GATE U2942 ( .I1(n1409), .I2(B[31]), .O(n1754) );
  NAND_GATE U2943 ( .I1(n1933), .I2(n1754), .O(n1755) );
  NAND_GATE U2944 ( .I1(A[10]), .I2(n1755), .O(n1756) );
  NAND_GATE U2945 ( .I1(n1757), .I2(n1756), .O(n1759) );
  NAND_GATE U2946 ( .I1(n1758), .I2(n1759), .O(n1763) );
  INV_GATE U2947 ( .I1(n1759), .O(n1760) );
  NAND_GATE U2948 ( .I1(n1761), .I2(n1760), .O(n1762) );
  NAND_GATE U2949 ( .I1(n1763), .I2(n1762), .O(n2138) );
  NAND_GATE U2950 ( .I1(n2136), .I2(n2138), .O(n2133) );
  NAND_GATE U2951 ( .I1(B[29]), .I2(A[11]), .O(n2126) );
  INV_GATE U2952 ( .I1(n2126), .O(n2119) );
  INV_GATE U2953 ( .I1(n1773), .O(n1770) );
  NAND_GATE U2954 ( .I1(n1407), .I2(B[30]), .O(n1764) );
  NAND_GATE U2955 ( .I1(n1930), .I2(n1764), .O(n1765) );
  NAND_GATE U2956 ( .I1(A[10]), .I2(n1765), .O(n1769) );
  NAND_GATE U2957 ( .I1(n1408), .I2(B[31]), .O(n1766) );
  NAND_GATE U2958 ( .I1(n1933), .I2(n1766), .O(n1767) );
  NAND_GATE U2959 ( .I1(A[9]), .I2(n1767), .O(n1768) );
  NAND_GATE U2960 ( .I1(n1769), .I2(n1768), .O(n1771) );
  NAND_GATE U2961 ( .I1(n1770), .I2(n1771), .O(n1775) );
  INV_GATE U2962 ( .I1(n1771), .O(n1772) );
  NAND_GATE U2963 ( .I1(n1773), .I2(n1772), .O(n1774) );
  NAND_GATE U2964 ( .I1(n1775), .I2(n1774), .O(n2121) );
  NAND_GATE U2965 ( .I1(n2119), .I2(n2121), .O(n2116) );
  NAND_GATE U2966 ( .I1(B[29]), .I2(A[10]), .O(n2104) );
  INV_GATE U2967 ( .I1(n2104), .O(n2097) );
  INV_GATE U2968 ( .I1(n1785), .O(n1782) );
  NAND_GATE U2969 ( .I1(n1406), .I2(B[30]), .O(n1776) );
  NAND_GATE U2970 ( .I1(n1930), .I2(n1776), .O(n1777) );
  NAND_GATE U2971 ( .I1(A[9]), .I2(n1777), .O(n1781) );
  NAND_GATE U2972 ( .I1(n1407), .I2(B[31]), .O(n1778) );
  NAND_GATE U2973 ( .I1(n1933), .I2(n1778), .O(n1779) );
  NAND_GATE U2974 ( .I1(A[8]), .I2(n1779), .O(n1780) );
  NAND_GATE U2975 ( .I1(n1781), .I2(n1780), .O(n1783) );
  NAND_GATE U2976 ( .I1(n1782), .I2(n1783), .O(n1787) );
  INV_GATE U2977 ( .I1(n1783), .O(n1784) );
  NAND_GATE U2978 ( .I1(n1785), .I2(n1784), .O(n1786) );
  NAND_GATE U2979 ( .I1(n1787), .I2(n1786), .O(n2099) );
  NAND_GATE U2980 ( .I1(n2097), .I2(n2099), .O(n2094) );
  NAND_GATE U2981 ( .I1(B[29]), .I2(A[9]), .O(n2089) );
  INV_GATE U2982 ( .I1(n2089), .O(n2082) );
  INV_GATE U2983 ( .I1(n1797), .O(n1794) );
  NAND_GATE U2984 ( .I1(n1405), .I2(B[30]), .O(n1788) );
  NAND_GATE U2985 ( .I1(n1930), .I2(n1788), .O(n1789) );
  NAND_GATE U2986 ( .I1(A[8]), .I2(n1789), .O(n1793) );
  NAND_GATE U2987 ( .I1(n1406), .I2(B[31]), .O(n1790) );
  NAND_GATE U2988 ( .I1(n1933), .I2(n1790), .O(n1791) );
  NAND_GATE U2989 ( .I1(A[7]), .I2(n1791), .O(n1792) );
  NAND_GATE U2990 ( .I1(n1793), .I2(n1792), .O(n1795) );
  NAND_GATE U2991 ( .I1(n1794), .I2(n1795), .O(n1799) );
  INV_GATE U2992 ( .I1(n1795), .O(n1796) );
  NAND_GATE U2993 ( .I1(n1797), .I2(n1796), .O(n1798) );
  NAND_GATE U2994 ( .I1(n1799), .I2(n1798), .O(n2084) );
  NAND_GATE U2995 ( .I1(n2082), .I2(n2084), .O(n2079) );
  NAND_GATE U2996 ( .I1(B[29]), .I2(A[8]), .O(n2072) );
  INV_GATE U2997 ( .I1(n2072), .O(n2066) );
  INV_GATE U2998 ( .I1(n1809), .O(n1806) );
  NAND_GATE U2999 ( .I1(n1404), .I2(B[30]), .O(n1800) );
  NAND_GATE U3000 ( .I1(n1930), .I2(n1800), .O(n1801) );
  NAND_GATE U3001 ( .I1(A[7]), .I2(n1801), .O(n1805) );
  NAND_GATE U3002 ( .I1(n1405), .I2(B[31]), .O(n1802) );
  NAND_GATE U3003 ( .I1(n1933), .I2(n1802), .O(n1803) );
  NAND_GATE U3004 ( .I1(A[6]), .I2(n1803), .O(n1804) );
  NAND_GATE U3005 ( .I1(n1805), .I2(n1804), .O(n1807) );
  NAND_GATE U3006 ( .I1(n1806), .I2(n1807), .O(n1811) );
  INV_GATE U3007 ( .I1(n1807), .O(n1808) );
  NAND_GATE U3008 ( .I1(n1809), .I2(n1808), .O(n1810) );
  NAND_GATE U3009 ( .I1(n1811), .I2(n1810), .O(n2067) );
  NAND_GATE U3010 ( .I1(n2066), .I2(n2067), .O(n2063) );
  NAND_GATE U3011 ( .I1(B[29]), .I2(A[7]), .O(n2056) );
  INV_GATE U3012 ( .I1(n2056), .O(n2049) );
  INV_GATE U3013 ( .I1(n1821), .O(n1818) );
  NAND_GATE U3014 ( .I1(n1403), .I2(B[30]), .O(n1812) );
  NAND_GATE U3015 ( .I1(n1930), .I2(n1812), .O(n1813) );
  NAND_GATE U3016 ( .I1(A[6]), .I2(n1813), .O(n1817) );
  NAND_GATE U3017 ( .I1(n1404), .I2(B[31]), .O(n1814) );
  NAND_GATE U3018 ( .I1(n1933), .I2(n1814), .O(n1815) );
  NAND_GATE U3019 ( .I1(A[5]), .I2(n1815), .O(n1816) );
  NAND_GATE U3020 ( .I1(n1817), .I2(n1816), .O(n1819) );
  NAND_GATE U3021 ( .I1(n1818), .I2(n1819), .O(n1823) );
  INV_GATE U3022 ( .I1(n1819), .O(n1820) );
  NAND_GATE U3023 ( .I1(n1821), .I2(n1820), .O(n1822) );
  NAND_GATE U3024 ( .I1(n1823), .I2(n1822), .O(n2051) );
  NAND_GATE U3025 ( .I1(n2049), .I2(n2051), .O(n2046) );
  NAND_GATE U3026 ( .I1(B[29]), .I2(A[6]), .O(n1976) );
  INV_GATE U3027 ( .I1(n1976), .O(n1969) );
  INV_GATE U3028 ( .I1(n1833), .O(n1830) );
  NAND_GATE U3029 ( .I1(n1402), .I2(B[30]), .O(n1824) );
  NAND_GATE U3030 ( .I1(n1930), .I2(n1824), .O(n1825) );
  NAND_GATE U3031 ( .I1(A[5]), .I2(n1825), .O(n1829) );
  NAND_GATE U3032 ( .I1(n1403), .I2(B[31]), .O(n1826) );
  NAND_GATE U3033 ( .I1(n1933), .I2(n1826), .O(n1827) );
  NAND_GATE U3034 ( .I1(A[4]), .I2(n1827), .O(n1828) );
  NAND_GATE U3035 ( .I1(n1829), .I2(n1828), .O(n1831) );
  NAND_GATE U3036 ( .I1(n1830), .I2(n1831), .O(n1835) );
  INV_GATE U3037 ( .I1(n1831), .O(n1832) );
  NAND_GATE U3038 ( .I1(n1833), .I2(n1832), .O(n1834) );
  NAND_GATE U3039 ( .I1(n1835), .I2(n1834), .O(n1971) );
  NAND_GATE U3040 ( .I1(n1969), .I2(n1971), .O(n1966) );
  NAND_GATE U3041 ( .I1(B[29]), .I2(A[5]), .O(n1988) );
  INV_GATE U3042 ( .I1(n1988), .O(n1982) );
  INV_GATE U3043 ( .I1(n1845), .O(n1842) );
  NAND_GATE U3044 ( .I1(n1401), .I2(B[30]), .O(n1836) );
  NAND_GATE U3045 ( .I1(n1930), .I2(n1836), .O(n1837) );
  NAND_GATE U3046 ( .I1(A[4]), .I2(n1837), .O(n1841) );
  NAND_GATE U3047 ( .I1(n1402), .I2(B[31]), .O(n1838) );
  NAND_GATE U3048 ( .I1(n1933), .I2(n1838), .O(n1839) );
  NAND_GATE U3049 ( .I1(A[3]), .I2(n1839), .O(n1840) );
  NAND_GATE U3050 ( .I1(n1841), .I2(n1840), .O(n1843) );
  NAND_GATE U3051 ( .I1(n1842), .I2(n1843), .O(n1847) );
  INV_GATE U3052 ( .I1(n1843), .O(n1844) );
  NAND_GATE U3053 ( .I1(n1845), .I2(n1844), .O(n1846) );
  NAND_GATE U3054 ( .I1(n1847), .I2(n1846), .O(n1985) );
  NAND_GATE U3055 ( .I1(n1982), .I2(n1985), .O(n1981) );
  NAND_GATE U3056 ( .I1(B[29]), .I2(A[4]), .O(n2035) );
  INV_GATE U3057 ( .I1(n2035), .O(n2034) );
  INV_GATE U3058 ( .I1(n1857), .O(n1854) );
  NAND_GATE U3059 ( .I1(n1400), .I2(B[30]), .O(n1848) );
  NAND_GATE U3060 ( .I1(n1930), .I2(n1848), .O(n1849) );
  NAND_GATE U3061 ( .I1(A[3]), .I2(n1849), .O(n1853) );
  NAND_GATE U3062 ( .I1(n1401), .I2(B[31]), .O(n1850) );
  NAND_GATE U3063 ( .I1(n1933), .I2(n1850), .O(n1851) );
  NAND_GATE U3064 ( .I1(A[2]), .I2(n1851), .O(n1852) );
  NAND_GATE U3065 ( .I1(n1853), .I2(n1852), .O(n1855) );
  NAND_GATE U3066 ( .I1(n1854), .I2(n1855), .O(n1859) );
  INV_GATE U3067 ( .I1(n1855), .O(n1856) );
  NAND_GATE U3068 ( .I1(n1857), .I2(n1856), .O(n1858) );
  NAND_GATE U3069 ( .I1(n1859), .I2(n1858), .O(n2029) );
  AND_GATE U3070 ( .I1(A[2]), .I2(B[30]), .O(n1861) );
  NAND_GATE U3071 ( .I1(B[31]), .I2(A[1]), .O(n1860) );
  NAND_GATE U3072 ( .I1(n1861), .I2(n1860), .O(n1870) );
  INV_GATE U3073 ( .I1(n1864), .O(n1863) );
  NAND_GATE U3074 ( .I1(n1863), .I2(n1862), .O(n1868) );
  NAND3_GATE U3075 ( .I1(B[31]), .I2(n1396), .I3(A[1]), .O(n1866) );
  NAND3_GATE U3076 ( .I1(B[31]), .I2(A[1]), .I3(n1400), .O(n1865) );
  NAND3_GATE U3077 ( .I1(n1866), .I2(n1865), .I3(n1864), .O(n1867) );
  NAND_GATE U3078 ( .I1(n1868), .I2(n1867), .O(n1869) );
  NAND_GATE U3079 ( .I1(n1870), .I2(n1869), .O(n1997) );
  NAND3_GATE U3080 ( .I1(B[29]), .I2(B[30]), .I3(n1196), .O(n2014) );
  INV_GATE U3081 ( .I1(n2014), .O(n2013) );
  NAND3_GATE U3082 ( .I1(B[30]), .I2(A[1]), .I3(n1397), .O(n1873) );
  NAND_GATE U3083 ( .I1(B[29]), .I2(A[2]), .O(n2011) );
  NAND_GATE U3084 ( .I1(n1873), .I2(n2011), .O(n1871) );
  NAND_GATE U3085 ( .I1(n2013), .I2(n1871), .O(n1877) );
  INV_GATE U3086 ( .I1(n2011), .O(n2018) );
  NAND3_GATE U3087 ( .I1(B[31]), .I2(n1399), .I3(A[0]), .O(n1875) );
  NAND3_GATE U3088 ( .I1(B[30]), .I2(A[1]), .I3(n1398), .O(n1874) );
  NAND3_GATE U3089 ( .I1(B[31]), .I2(n1396), .I3(A[0]), .O(n1872) );
  NAND4_GATE U3090 ( .I1(n1875), .I2(n1874), .I3(n1873), .I4(n1872), .O(n2012)
         );
  NAND_GATE U3091 ( .I1(n2018), .I2(n2012), .O(n1876) );
  NAND_GATE U3092 ( .I1(n1877), .I2(n1876), .O(n2000) );
  NAND_GATE U3093 ( .I1(n1997), .I2(n2000), .O(n2026) );
  NAND_GATE U3094 ( .I1(B[29]), .I2(A[3]), .O(n1993) );
  INV_GATE U3095 ( .I1(n1993), .O(n1998) );
  NAND_GATE U3096 ( .I1(n1998), .I2(n2000), .O(n2025) );
  NAND_GATE U3097 ( .I1(n1998), .I2(n1997), .O(n2027) );
  NAND3_GATE U3098 ( .I1(n2026), .I2(n2025), .I3(n2027), .O(n2028) );
  NAND_GATE U3099 ( .I1(n1858), .I2(n7), .O(n1878) );
  NAND_GATE U3100 ( .I1(n2028), .I2(n1878), .O(n1879) );
  NAND_GATE U3101 ( .I1(n2024), .I2(n1879), .O(n1986) );
  INV_GATE U3102 ( .I1(n1985), .O(n1987) );
  NAND_GATE U3103 ( .I1(n1988), .I2(n1987), .O(n1880) );
  NAND_GATE U3104 ( .I1(n1986), .I2(n1880), .O(n1970) );
  INV_GATE U3105 ( .I1(n1971), .O(n1973) );
  NAND_GATE U3106 ( .I1(n1976), .I2(n1973), .O(n1881) );
  NAND_GATE U3107 ( .I1(n1972), .I2(n1881), .O(n1882) );
  NAND_GATE U3108 ( .I1(n1966), .I2(n1882), .O(n2052) );
  INV_GATE U3109 ( .I1(n2051), .O(n2053) );
  NAND_GATE U3110 ( .I1(n2056), .I2(n2053), .O(n1883) );
  NAND_GATE U3111 ( .I1(n2052), .I2(n1883), .O(n1884) );
  NAND_GATE U3112 ( .I1(n2046), .I2(n1884), .O(n2068) );
  INV_GATE U3113 ( .I1(n2067), .O(n2069) );
  NAND_GATE U3114 ( .I1(n2072), .I2(n2069), .O(n1885) );
  NAND_GATE U3115 ( .I1(n2068), .I2(n1885), .O(n1886) );
  NAND_GATE U3116 ( .I1(n2063), .I2(n1886), .O(n2085) );
  INV_GATE U3117 ( .I1(n2084), .O(n2086) );
  NAND_GATE U3118 ( .I1(n2089), .I2(n2086), .O(n1887) );
  NAND_GATE U3119 ( .I1(n2085), .I2(n1887), .O(n1888) );
  NAND_GATE U3120 ( .I1(n2079), .I2(n1888), .O(n2100) );
  INV_GATE U3121 ( .I1(n2099), .O(n2101) );
  NAND_GATE U3122 ( .I1(n2104), .I2(n2101), .O(n1889) );
  NAND_GATE U3123 ( .I1(n2100), .I2(n1889), .O(n1890) );
  NAND_GATE U3124 ( .I1(n2094), .I2(n1890), .O(n2122) );
  INV_GATE U3125 ( .I1(n2121), .O(n2123) );
  NAND_GATE U3126 ( .I1(n2126), .I2(n2123), .O(n1891) );
  NAND_GATE U3127 ( .I1(n2122), .I2(n1891), .O(n1892) );
  NAND_GATE U3128 ( .I1(n2116), .I2(n1892), .O(n2139) );
  INV_GATE U3129 ( .I1(n2138), .O(n2140) );
  NAND_GATE U3130 ( .I1(n2143), .I2(n2140), .O(n1893) );
  NAND_GATE U3131 ( .I1(n2139), .I2(n1893), .O(n1894) );
  NAND_GATE U3132 ( .I1(n2133), .I2(n1894), .O(n2156) );
  INV_GATE U3133 ( .I1(n2155), .O(n2157) );
  NAND_GATE U3134 ( .I1(n2160), .I2(n2157), .O(n1895) );
  NAND_GATE U3135 ( .I1(n2156), .I2(n1895), .O(n1896) );
  NAND_GATE U3136 ( .I1(n2150), .I2(n1896), .O(n2173) );
  INV_GATE U3137 ( .I1(n2172), .O(n2174) );
  NAND_GATE U3138 ( .I1(n2177), .I2(n2174), .O(n1897) );
  NAND_GATE U3139 ( .I1(n2173), .I2(n1897), .O(n1898) );
  NAND_GATE U3140 ( .I1(n2167), .I2(n1898), .O(n2190) );
  INV_GATE U3141 ( .I1(n2189), .O(n2191) );
  NAND_GATE U3142 ( .I1(n2194), .I2(n2191), .O(n1899) );
  NAND_GATE U3143 ( .I1(n2190), .I2(n1899), .O(n1900) );
  NAND_GATE U3144 ( .I1(n2184), .I2(n1900), .O(n2207) );
  INV_GATE U3145 ( .I1(n2206), .O(n2208) );
  NAND_GATE U3146 ( .I1(n2211), .I2(n2208), .O(n1901) );
  NAND_GATE U3147 ( .I1(n2207), .I2(n1901), .O(n1902) );
  NAND_GATE U3148 ( .I1(n2201), .I2(n1902), .O(n2224) );
  INV_GATE U3149 ( .I1(n2223), .O(n2225) );
  NAND_GATE U3150 ( .I1(n2228), .I2(n2225), .O(n1903) );
  NAND_GATE U3151 ( .I1(n2224), .I2(n1903), .O(n1904) );
  NAND_GATE U3152 ( .I1(n2218), .I2(n1904), .O(n2240) );
  INV_GATE U3153 ( .I1(n2239), .O(n2241) );
  NAND_GATE U3154 ( .I1(n2244), .I2(n2241), .O(n1905) );
  NAND_GATE U3155 ( .I1(n2240), .I2(n1905), .O(n1906) );
  NAND_GATE U3156 ( .I1(n2234), .I2(n1906), .O(n2256) );
  INV_GATE U3157 ( .I1(n2255), .O(n2257) );
  NAND_GATE U3158 ( .I1(n2260), .I2(n2257), .O(n1907) );
  NAND_GATE U3159 ( .I1(n2256), .I2(n1907), .O(n1908) );
  NAND_GATE U3160 ( .I1(n2250), .I2(n1908), .O(n2272) );
  INV_GATE U3161 ( .I1(n2271), .O(n2273) );
  NAND_GATE U3162 ( .I1(n2276), .I2(n2273), .O(n1909) );
  NAND_GATE U3163 ( .I1(n2272), .I2(n1909), .O(n1910) );
  NAND_GATE U3164 ( .I1(n2266), .I2(n1910), .O(n2289) );
  INV_GATE U3165 ( .I1(n2288), .O(n2290) );
  NAND_GATE U3166 ( .I1(n2293), .I2(n2290), .O(n1911) );
  NAND_GATE U3167 ( .I1(n2289), .I2(n1911), .O(n1912) );
  NAND_GATE U3168 ( .I1(n2283), .I2(n1912), .O(n2306) );
  INV_GATE U3169 ( .I1(n2305), .O(n2307) );
  NAND_GATE U3170 ( .I1(n2310), .I2(n2307), .O(n1913) );
  NAND_GATE U3171 ( .I1(n2306), .I2(n1913), .O(n1914) );
  NAND_GATE U3172 ( .I1(n2300), .I2(n1914), .O(n2323) );
  INV_GATE U3173 ( .I1(n2322), .O(n2324) );
  NAND_GATE U3174 ( .I1(n2327), .I2(n2324), .O(n1915) );
  NAND_GATE U3175 ( .I1(n2323), .I2(n1915), .O(n1916) );
  NAND_GATE U3176 ( .I1(n2317), .I2(n1916), .O(n2340) );
  INV_GATE U3177 ( .I1(n2339), .O(n2341) );
  NAND_GATE U3178 ( .I1(n2344), .I2(n2341), .O(n1917) );
  NAND_GATE U3179 ( .I1(n2340), .I2(n1917), .O(n1918) );
  NAND_GATE U3180 ( .I1(n2334), .I2(n1918), .O(n2357) );
  INV_GATE U3181 ( .I1(n2356), .O(n2358) );
  NAND_GATE U3182 ( .I1(n2361), .I2(n2358), .O(n1919) );
  NAND_GATE U3183 ( .I1(n2357), .I2(n1919), .O(n1920) );
  NAND_GATE U3184 ( .I1(n2351), .I2(n1920), .O(n2374) );
  INV_GATE U3185 ( .I1(n2373), .O(n2375) );
  NAND_GATE U3186 ( .I1(n2378), .I2(n2375), .O(n1921) );
  NAND_GATE U3187 ( .I1(n2374), .I2(n1921), .O(n1922) );
  NAND_GATE U3188 ( .I1(n2368), .I2(n1922), .O(n2391) );
  INV_GATE U3189 ( .I1(n2390), .O(n2392) );
  NAND_GATE U3190 ( .I1(n2395), .I2(n2392), .O(n1923) );
  NAND_GATE U3191 ( .I1(n2391), .I2(n1923), .O(n1924) );
  NAND_GATE U3192 ( .I1(n2385), .I2(n1924), .O(n1957) );
  INV_GATE U3193 ( .I1(n1956), .O(n1958) );
  NAND_GATE U3194 ( .I1(n1961), .I2(n1958), .O(n1925) );
  NAND_GATE U3195 ( .I1(n1957), .I2(n1925), .O(n1926) );
  NAND_GATE U3196 ( .I1(n1951), .I2(n1926), .O(n2410) );
  INV_GATE U3197 ( .I1(n2409), .O(n2411) );
  NAND_GATE U3198 ( .I1(n2414), .I2(n2411), .O(n1927) );
  NAND_GATE U3199 ( .I1(n2410), .I2(n1927), .O(n1928) );
  NAND_GATE U3200 ( .I1(n2404), .I2(n1928), .O(n2428) );
  NAND_GATE U3201 ( .I1(n2424), .I2(n2428), .O(n2421) );
  INV_GATE U3202 ( .I1(n1940), .O(n1937) );
  NAND_GATE U3203 ( .I1(n1426), .I2(B[30]), .O(n1929) );
  NAND_GATE U3204 ( .I1(n1930), .I2(n1929), .O(n1931) );
  NAND_GATE U3205 ( .I1(A[29]), .I2(n1931), .O(n1936) );
  NAND_GATE U3206 ( .I1(n1933), .I2(n1932), .O(n1934) );
  NAND_GATE U3207 ( .I1(A[28]), .I2(n1934), .O(n1935) );
  NAND_GATE U3208 ( .I1(n1936), .I2(n1935), .O(n1938) );
  NAND_GATE U3209 ( .I1(n1937), .I2(n1938), .O(n1942) );
  INV_GATE U3210 ( .I1(n1938), .O(n1939) );
  NAND_GATE U3211 ( .I1(n1940), .I2(n1939), .O(n1941) );
  NAND_GATE U3212 ( .I1(n1942), .I2(n1941), .O(n2425) );
  INV_GATE U3213 ( .I1(n2428), .O(n2426) );
  NAND_GATE U3214 ( .I1(n2431), .I2(n2426), .O(n1943) );
  NAND_GATE U3215 ( .I1(n2425), .I2(n1943), .O(n1944) );
  NAND_GATE U3216 ( .I1(n2421), .I2(n1944), .O(n2444) );
  INV_GATE U3217 ( .I1(n2443), .O(n2445) );
  NAND_GATE U3218 ( .I1(n2448), .I2(n2445), .O(n1945) );
  NAND_GATE U3219 ( .I1(n2444), .I2(n1945), .O(n1946) );
  NAND_GATE U3220 ( .I1(n2438), .I2(n1946), .O(n15306) );
  NAND_GATE U3221 ( .I1(n1947), .I2(n15306), .O(n1950) );
  INV_GATE U3222 ( .I1(n15306), .O(n1948) );
  NAND_GATE U3223 ( .I1(n15307), .I2(n1948), .O(n1949) );
  NAND_GATE U3224 ( .I1(n1950), .I2(n1949), .O(\A1[59] ) );
  NAND_GATE U3225 ( .I1(B[28]), .I2(A[31]), .O(n2463) );
  INV_GATE U3226 ( .I1(n2463), .O(n2436) );
  NAND_GATE U3227 ( .I1(B[28]), .I2(A[30]), .O(n2474) );
  INV_GATE U3228 ( .I1(n2474), .O(n2419) );
  NAND_GATE U3229 ( .I1(B[28]), .I2(A[29]), .O(n2485) );
  INV_GATE U3230 ( .I1(n2485), .O(n2402) );
  INV_GATE U3231 ( .I1(n1951), .O(n1952) );
  NAND_GATE U3232 ( .I1(n1952), .I2(n1957), .O(n1965) );
  INV_GATE U3233 ( .I1(n1957), .O(n1955) );
  NAND_GATE U3234 ( .I1(n1958), .I2(n1955), .O(n1953) );
  NAND_GATE U3235 ( .I1(n1954), .I2(n1953), .O(n1963) );
  NAND_GATE U3236 ( .I1(n1956), .I2(n1955), .O(n1960) );
  NAND_GATE U3237 ( .I1(n1958), .I2(n1957), .O(n1959) );
  NAND3_GATE U3238 ( .I1(n1961), .I2(n1960), .I3(n1959), .O(n1962) );
  NAND_GATE U3239 ( .I1(n1963), .I2(n1962), .O(n1964) );
  NAND_GATE U3240 ( .I1(n1965), .I2(n1964), .O(n2483) );
  NAND_GATE U3241 ( .I1(n2402), .I2(n2483), .O(n2480) );
  NAND_GATE U3242 ( .I1(B[28]), .I2(A[28]), .O(n2496) );
  INV_GATE U3243 ( .I1(n2496), .O(n2400) );
  NAND_GATE U3244 ( .I1(B[28]), .I2(A[27]), .O(n2858) );
  INV_GATE U3245 ( .I1(n2858), .O(n2383) );
  NAND_GATE U3246 ( .I1(B[28]), .I2(A[26]), .O(n2507) );
  INV_GATE U3247 ( .I1(n2507), .O(n2366) );
  NAND_GATE U3248 ( .I1(B[28]), .I2(A[25]), .O(n2518) );
  INV_GATE U3249 ( .I1(n2518), .O(n2349) );
  NAND_GATE U3250 ( .I1(B[28]), .I2(A[24]), .O(n2529) );
  INV_GATE U3251 ( .I1(n2529), .O(n2332) );
  NAND_GATE U3252 ( .I1(B[28]), .I2(A[23]), .O(n2540) );
  INV_GATE U3253 ( .I1(n2540), .O(n2315) );
  NAND_GATE U3254 ( .I1(B[28]), .I2(A[22]), .O(n2551) );
  INV_GATE U3255 ( .I1(n2551), .O(n2298) );
  NAND_GATE U3256 ( .I1(B[28]), .I2(A[21]), .O(n2565) );
  INV_GATE U3257 ( .I1(n2565), .O(n2281) );
  NAND_GATE U3258 ( .I1(B[28]), .I2(A[20]), .O(n2579) );
  INV_GATE U3259 ( .I1(n2579), .O(n2265) );
  NAND_GATE U3260 ( .I1(B[28]), .I2(A[19]), .O(n2593) );
  INV_GATE U3261 ( .I1(n2593), .O(n2249) );
  NAND_GATE U3262 ( .I1(B[28]), .I2(A[18]), .O(n2604) );
  INV_GATE U3263 ( .I1(n2604), .O(n2233) );
  NAND_GATE U3264 ( .I1(B[28]), .I2(A[17]), .O(n2615) );
  INV_GATE U3265 ( .I1(n2615), .O(n2216) );
  NAND_GATE U3266 ( .I1(B[28]), .I2(A[16]), .O(n2626) );
  INV_GATE U3267 ( .I1(n2626), .O(n2199) );
  NAND_GATE U3268 ( .I1(B[28]), .I2(A[15]), .O(n2637) );
  INV_GATE U3269 ( .I1(n2637), .O(n2182) );
  NAND_GATE U3270 ( .I1(B[28]), .I2(A[14]), .O(n2648) );
  INV_GATE U3271 ( .I1(n2648), .O(n2165) );
  NAND_GATE U3272 ( .I1(B[28]), .I2(A[13]), .O(n2659) );
  INV_GATE U3273 ( .I1(n2659), .O(n2148) );
  NAND_GATE U3274 ( .I1(B[28]), .I2(A[12]), .O(n2670) );
  INV_GATE U3275 ( .I1(n2670), .O(n2131) );
  NAND_GATE U3276 ( .I1(B[28]), .I2(A[9]), .O(n2700) );
  INV_GATE U3277 ( .I1(n2700), .O(n2705) );
  NAND_GATE U3278 ( .I1(B[28]), .I2(A[8]), .O(n2711) );
  INV_GATE U3279 ( .I1(n2711), .O(n2715) );
  INV_GATE U3280 ( .I1(n1966), .O(n1967) );
  NAND_GATE U3281 ( .I1(n1967), .I2(n1972), .O(n1980) );
  OR_GATE U3282 ( .I1(n1972), .I2(n1971), .O(n1968) );
  NAND_GATE U3283 ( .I1(n1969), .I2(n1968), .O(n1978) );
  NAND3_GATE U3284 ( .I1(n1971), .I2(n1981), .I3(n1970), .O(n1975) );
  NAND_GATE U3285 ( .I1(n1973), .I2(n1972), .O(n1974) );
  NAND3_GATE U3286 ( .I1(n1976), .I2(n1975), .I3(n1974), .O(n1977) );
  NAND_GATE U3287 ( .I1(n1978), .I2(n1977), .O(n1979) );
  NAND_GATE U3288 ( .I1(B[28]), .I2(A[6]), .O(n2738) );
  INV_GATE U3289 ( .I1(n2738), .O(n2731) );
  NAND_GATE U3290 ( .I1(n1987), .I2(n663), .O(n1984) );
  NAND_GATE U3291 ( .I1(n797), .I2(n1986), .O(n1983) );
  NAND3_GATE U3292 ( .I1(n1984), .I2(n1983), .I3(n1982), .O(n1992) );
  NAND_GATE U3293 ( .I1(n1985), .I2(n663), .O(n1990) );
  NAND_GATE U3294 ( .I1(n1987), .I2(n1986), .O(n1989) );
  NAND3_GATE U3295 ( .I1(n1990), .I2(n1989), .I3(n1988), .O(n1991) );
  NAND_GATE U3296 ( .I1(n1992), .I2(n1991), .O(n2735) );
  INV_GATE U3297 ( .I1(n1997), .O(n1999) );
  NAND_GATE U3298 ( .I1(n1999), .I2(n2000), .O(n1995) );
  INV_GATE U3299 ( .I1(n2000), .O(n1996) );
  NAND_GATE U3300 ( .I1(n1997), .I2(n1996), .O(n1994) );
  NAND3_GATE U3301 ( .I1(n1997), .I2(n1996), .I3(n1998), .O(n2002) );
  NAND3_GATE U3302 ( .I1(n2000), .I2(n1999), .I3(n1998), .O(n2001) );
  NAND_GATE U3303 ( .I1(n2002), .I2(n2001), .O(n2003) );
  NAND_GATE U3304 ( .I1(B[28]), .I2(A[4]), .O(n2795) );
  INV_GATE U3305 ( .I1(n2795), .O(n2799) );
  NAND_GATE U3306 ( .I1(n2795), .I2(n2003), .O(n2744) );
  NAND_GATE U3307 ( .I1(n2795), .I2(n1307), .O(n2743) );
  NAND3_GATE U3308 ( .I1(B[28]), .I2(B[29]), .I3(n1196), .O(n2764) );
  INV_GATE U3309 ( .I1(n2764), .O(n2767) );
  NAND_GATE U3310 ( .I1(n1398), .I2(A[1]), .O(n14784) );
  NAND_GATE U3311 ( .I1(n1396), .I2(A[1]), .O(n2004) );
  NAND_GATE U3312 ( .I1(n14784), .I2(n2004), .O(n2005) );
  NAND_GATE U3313 ( .I1(B[29]), .I2(n2005), .O(n2758) );
  NAND_GATE U3314 ( .I1(A[0]), .I2(n1399), .O(n14781) );
  NAND_GATE U3315 ( .I1(n1395), .I2(A[0]), .O(n2006) );
  NAND_GATE U3316 ( .I1(n14781), .I2(n2006), .O(n2007) );
  NAND_GATE U3317 ( .I1(B[30]), .I2(n2007), .O(n2759) );
  NAND_GATE U3318 ( .I1(n2758), .I2(n2759), .O(n2765) );
  NAND_GATE U3319 ( .I1(B[28]), .I2(A[2]), .O(n2766) );
  NAND_GATE U3320 ( .I1(n2763), .I2(n2766), .O(n2008) );
  NAND_GATE U3321 ( .I1(n2767), .I2(n2008), .O(n2010) );
  INV_GATE U3322 ( .I1(n2766), .O(n2761) );
  NAND_GATE U3323 ( .I1(n2765), .I2(n2761), .O(n2009) );
  NAND_GATE U3324 ( .I1(n2010), .I2(n2009), .O(n2785) );
  NAND3_GATE U3325 ( .I1(n2013), .I2(n2018), .I3(n2012), .O(n2016) );
  NAND3_GATE U3326 ( .I1(n2014), .I2(n2011), .I3(n217), .O(n2020) );
  NAND_GATE U3327 ( .I1(n2013), .I2(n2012), .O(n2019) );
  NAND_GATE U3328 ( .I1(n2014), .I2(n217), .O(n2017) );
  NAND_GATE U3329 ( .I1(n2016), .I2(n2015), .O(n2786) );
  NAND_GATE U3330 ( .I1(n2785), .I2(n2786), .O(n2022) );
  NAND_GATE U3331 ( .I1(B[28]), .I2(A[3]), .O(n2787) );
  INV_GATE U3332 ( .I1(n2787), .O(n2781) );
  NAND_GATE U3333 ( .I1(n2018), .I2(n2017), .O(n2782) );
  NAND3_GATE U3334 ( .I1(n2781), .I2(n2782), .I3(n1194), .O(n2021) );
  NAND_GATE U3335 ( .I1(n2781), .I2(n2785), .O(n2780) );
  NAND3_GATE U3336 ( .I1(n2022), .I2(n2021), .I3(n2780), .O(n2794) );
  NAND3_GATE U3337 ( .I1(n2744), .I2(n2743), .I3(n2794), .O(n2023) );
  NAND_GATE U3338 ( .I1(n2742), .I2(n2023), .O(n2751) );
  NAND_GATE U3339 ( .I1(n225), .I2(n2028), .O(n2032) );
  NAND4_GATE U3340 ( .I1(n2027), .I2(n1297), .I3(n2026), .I4(n2025), .O(n2033)
         );
  NAND3_GATE U3341 ( .I1(n2032), .I2(n2033), .I3(n2034), .O(n2031) );
  NAND_GATE U3342 ( .I1(n1297), .I2(n2028), .O(n2036) );
  NAND3_GATE U3343 ( .I1(n2036), .I2(n2037), .I3(n2035), .O(n2030) );
  NAND_GATE U3344 ( .I1(n2031), .I2(n2030), .O(n2750) );
  INV_GATE U3345 ( .I1(n2750), .O(n2749) );
  NAND_GATE U3346 ( .I1(n2751), .I2(n2749), .O(n2041) );
  NAND_GATE U3347 ( .I1(B[28]), .I2(A[5]), .O(n2754) );
  INV_GATE U3348 ( .I1(n2754), .O(n2745) );
  NAND_GATE U3349 ( .I1(n2745), .I2(n2751), .O(n2040) );
  NAND3_GATE U3350 ( .I1(n2034), .I2(n2033), .I3(n2032), .O(n2039) );
  NAND3_GATE U3351 ( .I1(n2037), .I2(n2036), .I3(n2035), .O(n2038) );
  NAND3_GATE U3352 ( .I1(n2745), .I2(n2039), .I3(n2038), .O(n2741) );
  NAND3_GATE U3353 ( .I1(n2041), .I2(n2040), .I3(n2741), .O(n2734) );
  NAND_GATE U3354 ( .I1(n2738), .I2(n2735), .O(n2042) );
  NAND_GATE U3355 ( .I1(n2734), .I2(n2042), .O(n2043) );
  NAND_GATE U3356 ( .I1(n2730), .I2(n2043), .O(n2726) );
  NAND_GATE U3357 ( .I1(n2720), .I2(n2726), .O(n2045) );
  NAND_GATE U3358 ( .I1(B[28]), .I2(A[7]), .O(n2723) );
  INV_GATE U3359 ( .I1(n2723), .O(n2725) );
  NAND_GATE U3360 ( .I1(n2725), .I2(n2726), .O(n2044) );
  NAND_GATE U3361 ( .I1(n2725), .I2(n2720), .O(n2724) );
  NAND3_GATE U3362 ( .I1(n2045), .I2(n2044), .I3(n2724), .O(n2716) );
  NAND_GATE U3363 ( .I1(n2715), .I2(n2716), .O(n2062) );
  INV_GATE U3364 ( .I1(n2046), .O(n2047) );
  NAND_GATE U3365 ( .I1(n2047), .I2(n2052), .O(n2060) );
  INV_GATE U3366 ( .I1(n2052), .O(n2050) );
  NAND_GATE U3367 ( .I1(n2053), .I2(n2050), .O(n2048) );
  NAND_GATE U3368 ( .I1(n2049), .I2(n2048), .O(n2058) );
  NAND_GATE U3369 ( .I1(n2051), .I2(n2050), .O(n2055) );
  NAND_GATE U3370 ( .I1(n2053), .I2(n2052), .O(n2054) );
  NAND3_GATE U3371 ( .I1(n2056), .I2(n2055), .I3(n2054), .O(n2057) );
  NAND_GATE U3372 ( .I1(n2058), .I2(n2057), .O(n2059) );
  NAND_GATE U3373 ( .I1(n2060), .I2(n2059), .O(n2710) );
  NAND_GATE U3374 ( .I1(n2710), .I2(n2716), .O(n2061) );
  NAND_GATE U3375 ( .I1(n2715), .I2(n2710), .O(n2714) );
  NAND3_GATE U3376 ( .I1(n2062), .I2(n2061), .I3(n2714), .O(n2706) );
  NAND_GATE U3377 ( .I1(n2705), .I2(n2706), .O(n2078) );
  INV_GATE U3378 ( .I1(n2063), .O(n2064) );
  NAND_GATE U3379 ( .I1(n2064), .I2(n2068), .O(n2076) );
  NAND_GATE U3380 ( .I1(n2069), .I2(n6), .O(n2065) );
  NAND_GATE U3381 ( .I1(n2066), .I2(n2065), .O(n2074) );
  NAND_GATE U3382 ( .I1(n2067), .I2(n6), .O(n2071) );
  NAND_GATE U3383 ( .I1(n2069), .I2(n2068), .O(n2070) );
  NAND3_GATE U3384 ( .I1(n2072), .I2(n2071), .I3(n2070), .O(n2073) );
  NAND_GATE U3385 ( .I1(n2074), .I2(n2073), .O(n2075) );
  NAND_GATE U3386 ( .I1(n2076), .I2(n2075), .O(n2699) );
  NAND_GATE U3387 ( .I1(n2699), .I2(n2706), .O(n2077) );
  NAND_GATE U3388 ( .I1(n2705), .I2(n2699), .O(n2703) );
  NAND3_GATE U3389 ( .I1(n2078), .I2(n2077), .I3(n2703), .O(n2689) );
  NAND_GATE U3390 ( .I1(B[28]), .I2(A[11]), .O(n2678) );
  INV_GATE U3391 ( .I1(n2678), .O(n2681) );
  INV_GATE U3392 ( .I1(n2079), .O(n2080) );
  NAND_GATE U3393 ( .I1(n2080), .I2(n2085), .O(n2093) );
  INV_GATE U3394 ( .I1(n2085), .O(n2083) );
  NAND_GATE U3395 ( .I1(n2086), .I2(n2083), .O(n2081) );
  NAND_GATE U3396 ( .I1(n2082), .I2(n2081), .O(n2091) );
  NAND_GATE U3397 ( .I1(n2084), .I2(n2083), .O(n2088) );
  NAND_GATE U3398 ( .I1(n2086), .I2(n2085), .O(n2087) );
  NAND3_GATE U3399 ( .I1(n2089), .I2(n2088), .I3(n2087), .O(n2090) );
  NAND_GATE U3400 ( .I1(n2091), .I2(n2090), .O(n2092) );
  NAND_GATE U3401 ( .I1(n2093), .I2(n2092), .O(n2692) );
  NAND3_GATE U3402 ( .I1(n2689), .I2(n2681), .I3(n2692), .O(n2115) );
  NAND_GATE U3403 ( .I1(B[28]), .I2(A[10]), .O(n2695) );
  INV_GATE U3404 ( .I1(n2695), .O(n2687) );
  NAND3_GATE U3405 ( .I1(n2687), .I2(n2681), .I3(n2689), .O(n2114) );
  INV_GATE U3406 ( .I1(n2094), .O(n2095) );
  NAND_GATE U3407 ( .I1(n2095), .I2(n2100), .O(n2108) );
  INV_GATE U3408 ( .I1(n2100), .O(n2098) );
  NAND_GATE U3409 ( .I1(n2101), .I2(n2098), .O(n2096) );
  NAND_GATE U3410 ( .I1(n2097), .I2(n2096), .O(n2106) );
  NAND_GATE U3411 ( .I1(n2099), .I2(n2098), .O(n2103) );
  NAND_GATE U3412 ( .I1(n2101), .I2(n2100), .O(n2102) );
  NAND3_GATE U3413 ( .I1(n2104), .I2(n2103), .I3(n2102), .O(n2105) );
  NAND_GATE U3414 ( .I1(n2106), .I2(n2105), .O(n2107) );
  NAND_GATE U3415 ( .I1(n2108), .I2(n2107), .O(n2675) );
  NAND_GATE U3416 ( .I1(n2687), .I2(n2689), .O(n2110) );
  NAND_GATE U3417 ( .I1(n2692), .I2(n2689), .O(n2109) );
  NAND_GATE U3418 ( .I1(n2687), .I2(n2692), .O(n2111) );
  NAND3_GATE U3419 ( .I1(n2110), .I2(n2109), .I3(n2111), .O(n2680) );
  NAND_GATE U3420 ( .I1(n2675), .I2(n2680), .O(n2113) );
  NAND_GATE U3421 ( .I1(n2681), .I2(n2675), .O(n2684) );
  INV_GATE U3422 ( .I1(n2111), .O(n2688) );
  NAND_GATE U3423 ( .I1(n2681), .I2(n2688), .O(n2112) );
  NAND5_GATE U3424 ( .I1(n2115), .I2(n2114), .I3(n2113), .I4(n2684), .I5(n2112), .O(n2669) );
  NAND_GATE U3425 ( .I1(n2131), .I2(n2669), .O(n2665) );
  INV_GATE U3426 ( .I1(n2116), .O(n2117) );
  NAND_GATE U3427 ( .I1(n2117), .I2(n2122), .O(n2130) );
  INV_GATE U3428 ( .I1(n2122), .O(n2120) );
  NAND_GATE U3429 ( .I1(n2123), .I2(n2120), .O(n2118) );
  NAND_GATE U3430 ( .I1(n2119), .I2(n2118), .O(n2128) );
  NAND_GATE U3431 ( .I1(n2121), .I2(n2120), .O(n2125) );
  NAND_GATE U3432 ( .I1(n2123), .I2(n2122), .O(n2124) );
  NAND3_GATE U3433 ( .I1(n2126), .I2(n2125), .I3(n2124), .O(n2127) );
  NAND_GATE U3434 ( .I1(n2128), .I2(n2127), .O(n2129) );
  NAND_GATE U3435 ( .I1(n2130), .I2(n2129), .O(n2668) );
  NAND_GATE U3436 ( .I1(n2131), .I2(n2668), .O(n2664) );
  NAND_GATE U3437 ( .I1(n2669), .I2(n2668), .O(n2132) );
  NAND3_GATE U3438 ( .I1(n2665), .I2(n2664), .I3(n2132), .O(n2658) );
  NAND_GATE U3439 ( .I1(n2148), .I2(n2658), .O(n2654) );
  INV_GATE U3440 ( .I1(n2133), .O(n2134) );
  NAND_GATE U3441 ( .I1(n2134), .I2(n2139), .O(n2147) );
  INV_GATE U3442 ( .I1(n2139), .O(n2137) );
  NAND_GATE U3443 ( .I1(n2140), .I2(n2137), .O(n2135) );
  NAND_GATE U3444 ( .I1(n2136), .I2(n2135), .O(n2145) );
  NAND_GATE U3445 ( .I1(n2138), .I2(n2137), .O(n2142) );
  NAND_GATE U3446 ( .I1(n2140), .I2(n2139), .O(n2141) );
  NAND3_GATE U3447 ( .I1(n2143), .I2(n2142), .I3(n2141), .O(n2144) );
  NAND_GATE U3448 ( .I1(n2145), .I2(n2144), .O(n2146) );
  NAND_GATE U3449 ( .I1(n2147), .I2(n2146), .O(n2657) );
  NAND_GATE U3450 ( .I1(n2148), .I2(n2657), .O(n2653) );
  NAND_GATE U3451 ( .I1(n2658), .I2(n2657), .O(n2149) );
  NAND3_GATE U3452 ( .I1(n2654), .I2(n2653), .I3(n2149), .O(n2647) );
  NAND_GATE U3453 ( .I1(n2165), .I2(n2647), .O(n2643) );
  INV_GATE U3454 ( .I1(n2150), .O(n2151) );
  NAND_GATE U3455 ( .I1(n2151), .I2(n2156), .O(n2164) );
  INV_GATE U3456 ( .I1(n2156), .O(n2154) );
  NAND_GATE U3457 ( .I1(n2157), .I2(n2154), .O(n2152) );
  NAND_GATE U3458 ( .I1(n2153), .I2(n2152), .O(n2162) );
  NAND_GATE U3459 ( .I1(n2155), .I2(n2154), .O(n2159) );
  NAND_GATE U3460 ( .I1(n2157), .I2(n2156), .O(n2158) );
  NAND3_GATE U3461 ( .I1(n2160), .I2(n2159), .I3(n2158), .O(n2161) );
  NAND_GATE U3462 ( .I1(n2162), .I2(n2161), .O(n2163) );
  NAND_GATE U3463 ( .I1(n2164), .I2(n2163), .O(n2646) );
  NAND_GATE U3464 ( .I1(n2165), .I2(n2646), .O(n2642) );
  NAND_GATE U3465 ( .I1(n2647), .I2(n2646), .O(n2166) );
  NAND3_GATE U3466 ( .I1(n2643), .I2(n2642), .I3(n2166), .O(n2636) );
  NAND_GATE U3467 ( .I1(n2182), .I2(n2636), .O(n2632) );
  INV_GATE U3468 ( .I1(n2167), .O(n2168) );
  NAND_GATE U3469 ( .I1(n2168), .I2(n2173), .O(n2181) );
  INV_GATE U3470 ( .I1(n2173), .O(n2171) );
  NAND_GATE U3471 ( .I1(n2174), .I2(n2171), .O(n2169) );
  NAND_GATE U3472 ( .I1(n2170), .I2(n2169), .O(n2179) );
  NAND_GATE U3473 ( .I1(n2172), .I2(n2171), .O(n2176) );
  NAND_GATE U3474 ( .I1(n2174), .I2(n2173), .O(n2175) );
  NAND3_GATE U3475 ( .I1(n2177), .I2(n2176), .I3(n2175), .O(n2178) );
  NAND_GATE U3476 ( .I1(n2179), .I2(n2178), .O(n2180) );
  NAND_GATE U3477 ( .I1(n2181), .I2(n2180), .O(n2635) );
  NAND_GATE U3478 ( .I1(n2182), .I2(n2635), .O(n2631) );
  NAND_GATE U3479 ( .I1(n2636), .I2(n2635), .O(n2183) );
  NAND3_GATE U3480 ( .I1(n2632), .I2(n2631), .I3(n2183), .O(n2625) );
  NAND_GATE U3481 ( .I1(n2199), .I2(n2625), .O(n2621) );
  INV_GATE U3482 ( .I1(n2184), .O(n2185) );
  NAND_GATE U3483 ( .I1(n2185), .I2(n2190), .O(n2198) );
  INV_GATE U3484 ( .I1(n2190), .O(n2188) );
  NAND_GATE U3485 ( .I1(n2191), .I2(n2188), .O(n2186) );
  NAND_GATE U3486 ( .I1(n2187), .I2(n2186), .O(n2196) );
  NAND_GATE U3487 ( .I1(n2189), .I2(n2188), .O(n2193) );
  NAND_GATE U3488 ( .I1(n2191), .I2(n2190), .O(n2192) );
  NAND3_GATE U3489 ( .I1(n2194), .I2(n2193), .I3(n2192), .O(n2195) );
  NAND_GATE U3490 ( .I1(n2196), .I2(n2195), .O(n2197) );
  NAND_GATE U3491 ( .I1(n2198), .I2(n2197), .O(n2624) );
  NAND_GATE U3492 ( .I1(n2199), .I2(n2624), .O(n2620) );
  NAND_GATE U3493 ( .I1(n2625), .I2(n2624), .O(n2200) );
  NAND3_GATE U3494 ( .I1(n2621), .I2(n2620), .I3(n2200), .O(n2614) );
  NAND_GATE U3495 ( .I1(n2216), .I2(n2614), .O(n2610) );
  INV_GATE U3496 ( .I1(n2201), .O(n2202) );
  NAND_GATE U3497 ( .I1(n2202), .I2(n2207), .O(n2215) );
  INV_GATE U3498 ( .I1(n2207), .O(n2205) );
  NAND_GATE U3499 ( .I1(n2208), .I2(n2205), .O(n2203) );
  NAND_GATE U3500 ( .I1(n2204), .I2(n2203), .O(n2213) );
  NAND_GATE U3501 ( .I1(n2206), .I2(n2205), .O(n2210) );
  NAND_GATE U3502 ( .I1(n2208), .I2(n2207), .O(n2209) );
  NAND3_GATE U3503 ( .I1(n2211), .I2(n2210), .I3(n2209), .O(n2212) );
  NAND_GATE U3504 ( .I1(n2213), .I2(n2212), .O(n2214) );
  NAND_GATE U3505 ( .I1(n2215), .I2(n2214), .O(n2613) );
  NAND_GATE U3506 ( .I1(n2216), .I2(n2613), .O(n2609) );
  NAND_GATE U3507 ( .I1(n2614), .I2(n2613), .O(n2217) );
  NAND3_GATE U3508 ( .I1(n2610), .I2(n2609), .I3(n2217), .O(n2603) );
  NAND_GATE U3509 ( .I1(n2233), .I2(n2603), .O(n2599) );
  INV_GATE U3510 ( .I1(n2218), .O(n2219) );
  NAND_GATE U3511 ( .I1(n2219), .I2(n2224), .O(n2232) );
  INV_GATE U3512 ( .I1(n2224), .O(n2222) );
  NAND_GATE U3513 ( .I1(n2225), .I2(n2222), .O(n2220) );
  NAND_GATE U3514 ( .I1(n2221), .I2(n2220), .O(n2230) );
  NAND_GATE U3515 ( .I1(n2223), .I2(n2222), .O(n2227) );
  NAND_GATE U3516 ( .I1(n2225), .I2(n2224), .O(n2226) );
  NAND3_GATE U3517 ( .I1(n2228), .I2(n2227), .I3(n2226), .O(n2229) );
  NAND_GATE U3518 ( .I1(n2230), .I2(n2229), .O(n2231) );
  NAND_GATE U3519 ( .I1(n2232), .I2(n2231), .O(n2602) );
  NAND_GATE U3520 ( .I1(n2233), .I2(n2602), .O(n2598) );
  NAND_GATE U3521 ( .I1(n2599), .I2(n2598), .O(n2589) );
  NAND_GATE U3522 ( .I1(n2603), .I2(n2602), .O(n2588) );
  NAND_GATE U3523 ( .I1(n2249), .I2(n2590), .O(n2585) );
  INV_GATE U3524 ( .I1(n2234), .O(n2235) );
  NAND_GATE U3525 ( .I1(n2235), .I2(n2240), .O(n2248) );
  INV_GATE U3526 ( .I1(n2240), .O(n2238) );
  NAND_GATE U3527 ( .I1(n2241), .I2(n2238), .O(n2236) );
  NAND_GATE U3528 ( .I1(n2237), .I2(n2236), .O(n2246) );
  NAND_GATE U3529 ( .I1(n2239), .I2(n2238), .O(n2243) );
  NAND_GATE U3530 ( .I1(n2241), .I2(n2240), .O(n2242) );
  NAND3_GATE U3531 ( .I1(n2244), .I2(n2243), .I3(n2242), .O(n2245) );
  NAND_GATE U3532 ( .I1(n2246), .I2(n2245), .O(n2247) );
  NAND_GATE U3533 ( .I1(n2248), .I2(n2247), .O(n2591) );
  NAND_GATE U3534 ( .I1(n2249), .I2(n2591), .O(n2584) );
  NAND_GATE U3535 ( .I1(n2585), .I2(n2584), .O(n2575) );
  NAND_GATE U3536 ( .I1(n2590), .I2(n2591), .O(n2574) );
  NAND_GATE U3537 ( .I1(n2265), .I2(n2576), .O(n2571) );
  INV_GATE U3538 ( .I1(n2250), .O(n2251) );
  NAND_GATE U3539 ( .I1(n2251), .I2(n2256), .O(n2264) );
  INV_GATE U3540 ( .I1(n2256), .O(n2254) );
  NAND_GATE U3541 ( .I1(n2257), .I2(n2254), .O(n2252) );
  NAND_GATE U3542 ( .I1(n2253), .I2(n2252), .O(n2262) );
  NAND_GATE U3543 ( .I1(n2255), .I2(n2254), .O(n2259) );
  NAND_GATE U3544 ( .I1(n2257), .I2(n2256), .O(n2258) );
  NAND3_GATE U3545 ( .I1(n2260), .I2(n2259), .I3(n2258), .O(n2261) );
  NAND_GATE U3546 ( .I1(n2262), .I2(n2261), .O(n2263) );
  NAND_GATE U3547 ( .I1(n2264), .I2(n2263), .O(n2577) );
  NAND_GATE U3548 ( .I1(n2265), .I2(n2577), .O(n2570) );
  NAND_GATE U3549 ( .I1(n2571), .I2(n2570), .O(n2561) );
  NAND_GATE U3550 ( .I1(n2576), .I2(n2577), .O(n2560) );
  NAND_GATE U3551 ( .I1(n2281), .I2(n2562), .O(n2557) );
  INV_GATE U3552 ( .I1(n2266), .O(n2267) );
  NAND_GATE U3553 ( .I1(n2267), .I2(n2272), .O(n2280) );
  INV_GATE U3554 ( .I1(n2272), .O(n2270) );
  NAND_GATE U3555 ( .I1(n2273), .I2(n2270), .O(n2268) );
  NAND_GATE U3556 ( .I1(n2269), .I2(n2268), .O(n2278) );
  NAND_GATE U3557 ( .I1(n2271), .I2(n2270), .O(n2275) );
  NAND_GATE U3558 ( .I1(n2273), .I2(n2272), .O(n2274) );
  NAND3_GATE U3559 ( .I1(n2276), .I2(n2275), .I3(n2274), .O(n2277) );
  NAND_GATE U3560 ( .I1(n2278), .I2(n2277), .O(n2279) );
  NAND_GATE U3561 ( .I1(n2280), .I2(n2279), .O(n2563) );
  NAND_GATE U3562 ( .I1(n2281), .I2(n2563), .O(n2556) );
  NAND_GATE U3563 ( .I1(n2562), .I2(n2563), .O(n2282) );
  NAND3_GATE U3564 ( .I1(n2557), .I2(n2556), .I3(n2282), .O(n2550) );
  NAND_GATE U3565 ( .I1(n2298), .I2(n2550), .O(n2546) );
  INV_GATE U3566 ( .I1(n2283), .O(n2284) );
  NAND_GATE U3567 ( .I1(n2284), .I2(n2289), .O(n2297) );
  INV_GATE U3568 ( .I1(n2289), .O(n2287) );
  NAND_GATE U3569 ( .I1(n2290), .I2(n2287), .O(n2285) );
  NAND_GATE U3570 ( .I1(n2286), .I2(n2285), .O(n2295) );
  NAND_GATE U3571 ( .I1(n2288), .I2(n2287), .O(n2292) );
  NAND_GATE U3572 ( .I1(n2290), .I2(n2289), .O(n2291) );
  NAND3_GATE U3573 ( .I1(n2293), .I2(n2292), .I3(n2291), .O(n2294) );
  NAND_GATE U3574 ( .I1(n2295), .I2(n2294), .O(n2296) );
  NAND_GATE U3575 ( .I1(n2297), .I2(n2296), .O(n2549) );
  NAND_GATE U3576 ( .I1(n2298), .I2(n2549), .O(n2545) );
  NAND_GATE U3577 ( .I1(n2550), .I2(n2549), .O(n2299) );
  NAND3_GATE U3578 ( .I1(n2546), .I2(n2545), .I3(n2299), .O(n2539) );
  NAND_GATE U3579 ( .I1(n2315), .I2(n2539), .O(n2535) );
  INV_GATE U3580 ( .I1(n2300), .O(n2301) );
  NAND_GATE U3581 ( .I1(n2301), .I2(n2306), .O(n2314) );
  INV_GATE U3582 ( .I1(n2306), .O(n2304) );
  NAND_GATE U3583 ( .I1(n2307), .I2(n2304), .O(n2302) );
  NAND_GATE U3584 ( .I1(n2303), .I2(n2302), .O(n2312) );
  NAND_GATE U3585 ( .I1(n2305), .I2(n2304), .O(n2309) );
  NAND_GATE U3586 ( .I1(n2307), .I2(n2306), .O(n2308) );
  NAND3_GATE U3587 ( .I1(n2310), .I2(n2309), .I3(n2308), .O(n2311) );
  NAND_GATE U3588 ( .I1(n2312), .I2(n2311), .O(n2313) );
  NAND_GATE U3589 ( .I1(n2314), .I2(n2313), .O(n2538) );
  NAND_GATE U3590 ( .I1(n2315), .I2(n2538), .O(n2534) );
  NAND_GATE U3591 ( .I1(n2539), .I2(n2538), .O(n2316) );
  NAND3_GATE U3592 ( .I1(n2535), .I2(n2534), .I3(n2316), .O(n2528) );
  NAND_GATE U3593 ( .I1(n2332), .I2(n2528), .O(n2524) );
  INV_GATE U3594 ( .I1(n2317), .O(n2318) );
  NAND_GATE U3595 ( .I1(n2318), .I2(n2323), .O(n2331) );
  INV_GATE U3596 ( .I1(n2323), .O(n2321) );
  NAND_GATE U3597 ( .I1(n2324), .I2(n2321), .O(n2319) );
  NAND_GATE U3598 ( .I1(n2320), .I2(n2319), .O(n2329) );
  NAND_GATE U3599 ( .I1(n2322), .I2(n2321), .O(n2326) );
  NAND_GATE U3600 ( .I1(n2324), .I2(n2323), .O(n2325) );
  NAND3_GATE U3601 ( .I1(n2327), .I2(n2326), .I3(n2325), .O(n2328) );
  NAND_GATE U3602 ( .I1(n2329), .I2(n2328), .O(n2330) );
  NAND_GATE U3603 ( .I1(n2331), .I2(n2330), .O(n2527) );
  NAND_GATE U3604 ( .I1(n2332), .I2(n2527), .O(n2523) );
  NAND_GATE U3605 ( .I1(n2528), .I2(n2527), .O(n2333) );
  NAND3_GATE U3606 ( .I1(n2524), .I2(n2523), .I3(n2333), .O(n2517) );
  NAND_GATE U3607 ( .I1(n2349), .I2(n2517), .O(n2513) );
  INV_GATE U3608 ( .I1(n2334), .O(n2335) );
  NAND_GATE U3609 ( .I1(n2335), .I2(n2340), .O(n2348) );
  INV_GATE U3610 ( .I1(n2340), .O(n2338) );
  NAND_GATE U3611 ( .I1(n2341), .I2(n2338), .O(n2336) );
  NAND_GATE U3612 ( .I1(n2337), .I2(n2336), .O(n2346) );
  NAND_GATE U3613 ( .I1(n2339), .I2(n2338), .O(n2343) );
  NAND_GATE U3614 ( .I1(n2341), .I2(n2340), .O(n2342) );
  NAND3_GATE U3615 ( .I1(n2344), .I2(n2343), .I3(n2342), .O(n2345) );
  NAND_GATE U3616 ( .I1(n2346), .I2(n2345), .O(n2347) );
  NAND_GATE U3617 ( .I1(n2348), .I2(n2347), .O(n2516) );
  NAND_GATE U3618 ( .I1(n2349), .I2(n2516), .O(n2512) );
  NAND_GATE U3619 ( .I1(n2517), .I2(n2516), .O(n2350) );
  NAND3_GATE U3620 ( .I1(n2513), .I2(n2512), .I3(n2350), .O(n2506) );
  NAND_GATE U3621 ( .I1(n2366), .I2(n2506), .O(n2502) );
  INV_GATE U3622 ( .I1(n2351), .O(n2352) );
  NAND_GATE U3623 ( .I1(n2352), .I2(n2357), .O(n2365) );
  INV_GATE U3624 ( .I1(n2357), .O(n2355) );
  NAND_GATE U3625 ( .I1(n2358), .I2(n2355), .O(n2353) );
  NAND_GATE U3626 ( .I1(n2354), .I2(n2353), .O(n2363) );
  NAND_GATE U3627 ( .I1(n2356), .I2(n2355), .O(n2360) );
  NAND_GATE U3628 ( .I1(n2358), .I2(n2357), .O(n2359) );
  NAND3_GATE U3629 ( .I1(n2361), .I2(n2360), .I3(n2359), .O(n2362) );
  NAND_GATE U3630 ( .I1(n2363), .I2(n2362), .O(n2364) );
  NAND_GATE U3631 ( .I1(n2365), .I2(n2364), .O(n2505) );
  NAND_GATE U3632 ( .I1(n2366), .I2(n2505), .O(n2501) );
  NAND_GATE U3633 ( .I1(n2506), .I2(n2505), .O(n2367) );
  NAND3_GATE U3634 ( .I1(n2502), .I2(n2501), .I3(n2367), .O(n2857) );
  NAND_GATE U3635 ( .I1(n2383), .I2(n2857), .O(n2853) );
  INV_GATE U3636 ( .I1(n2368), .O(n2369) );
  NAND_GATE U3637 ( .I1(n2369), .I2(n2374), .O(n2382) );
  INV_GATE U3638 ( .I1(n2374), .O(n2372) );
  NAND_GATE U3639 ( .I1(n2375), .I2(n2372), .O(n2370) );
  NAND_GATE U3640 ( .I1(n2371), .I2(n2370), .O(n2380) );
  NAND_GATE U3641 ( .I1(n2373), .I2(n2372), .O(n2377) );
  NAND_GATE U3642 ( .I1(n2375), .I2(n2374), .O(n2376) );
  NAND3_GATE U3643 ( .I1(n2378), .I2(n2377), .I3(n2376), .O(n2379) );
  NAND_GATE U3644 ( .I1(n2380), .I2(n2379), .O(n2381) );
  NAND_GATE U3645 ( .I1(n2382), .I2(n2381), .O(n2856) );
  NAND_GATE U3646 ( .I1(n2383), .I2(n2856), .O(n2852) );
  NAND_GATE U3647 ( .I1(n2857), .I2(n2856), .O(n2384) );
  NAND3_GATE U3648 ( .I1(n2853), .I2(n2852), .I3(n2384), .O(n2495) );
  NAND_GATE U3649 ( .I1(n2400), .I2(n2495), .O(n2491) );
  INV_GATE U3650 ( .I1(n2385), .O(n2386) );
  NAND_GATE U3651 ( .I1(n2386), .I2(n2391), .O(n2399) );
  INV_GATE U3652 ( .I1(n2391), .O(n2389) );
  NAND_GATE U3653 ( .I1(n2392), .I2(n2389), .O(n2387) );
  NAND_GATE U3654 ( .I1(n2388), .I2(n2387), .O(n2397) );
  NAND_GATE U3655 ( .I1(n2390), .I2(n2389), .O(n2394) );
  NAND_GATE U3656 ( .I1(n2392), .I2(n2391), .O(n2393) );
  NAND3_GATE U3657 ( .I1(n2395), .I2(n2394), .I3(n2393), .O(n2396) );
  NAND_GATE U3658 ( .I1(n2397), .I2(n2396), .O(n2398) );
  NAND_GATE U3659 ( .I1(n2399), .I2(n2398), .O(n2494) );
  NAND_GATE U3660 ( .I1(n2400), .I2(n2494), .O(n2490) );
  NAND_GATE U3661 ( .I1(n2495), .I2(n2494), .O(n2401) );
  NAND3_GATE U3662 ( .I1(n2491), .I2(n2490), .I3(n2401), .O(n2484) );
  NAND_GATE U3663 ( .I1(n2402), .I2(n2484), .O(n2479) );
  NAND_GATE U3664 ( .I1(n2483), .I2(n2484), .O(n2403) );
  NAND3_GATE U3665 ( .I1(n2480), .I2(n2479), .I3(n2403), .O(n2473) );
  NAND_GATE U3666 ( .I1(n2419), .I2(n2473), .O(n2469) );
  INV_GATE U3667 ( .I1(n2404), .O(n2405) );
  NAND_GATE U3668 ( .I1(n2405), .I2(n2410), .O(n2418) );
  INV_GATE U3669 ( .I1(n2410), .O(n2408) );
  NAND_GATE U3670 ( .I1(n2411), .I2(n2408), .O(n2406) );
  NAND_GATE U3671 ( .I1(n2407), .I2(n2406), .O(n2416) );
  NAND_GATE U3672 ( .I1(n2409), .I2(n2408), .O(n2413) );
  NAND_GATE U3673 ( .I1(n2411), .I2(n2410), .O(n2412) );
  NAND3_GATE U3674 ( .I1(n2414), .I2(n2413), .I3(n2412), .O(n2415) );
  NAND_GATE U3675 ( .I1(n2416), .I2(n2415), .O(n2417) );
  NAND_GATE U3676 ( .I1(n2418), .I2(n2417), .O(n2472) );
  NAND_GATE U3677 ( .I1(n2419), .I2(n2472), .O(n2468) );
  NAND_GATE U3678 ( .I1(n2473), .I2(n2472), .O(n2420) );
  NAND3_GATE U3679 ( .I1(n2469), .I2(n2468), .I3(n2420), .O(n2462) );
  NAND_GATE U3680 ( .I1(n2436), .I2(n2462), .O(n2458) );
  INV_GATE U3681 ( .I1(n2421), .O(n2422) );
  NAND_GATE U3682 ( .I1(n2422), .I2(n2425), .O(n2435) );
  INV_GATE U3683 ( .I1(n2425), .O(n2427) );
  NAND_GATE U3684 ( .I1(n2426), .I2(n2427), .O(n2423) );
  NAND_GATE U3685 ( .I1(n2424), .I2(n2423), .O(n2433) );
  NAND_GATE U3686 ( .I1(n2426), .I2(n2425), .O(n2430) );
  NAND_GATE U3687 ( .I1(n2428), .I2(n2427), .O(n2429) );
  NAND3_GATE U3688 ( .I1(n2431), .I2(n2430), .I3(n2429), .O(n2432) );
  NAND_GATE U3689 ( .I1(n2433), .I2(n2432), .O(n2434) );
  NAND_GATE U3690 ( .I1(n2435), .I2(n2434), .O(n2461) );
  NAND_GATE U3691 ( .I1(n2436), .I2(n2461), .O(n2457) );
  NAND_GATE U3692 ( .I1(n2462), .I2(n2461), .O(n2437) );
  NAND3_GATE U3693 ( .I1(n2458), .I2(n2457), .I3(n2437), .O(n15309) );
  INV_GATE U3694 ( .I1(n15309), .O(n2453) );
  INV_GATE U3695 ( .I1(n2438), .O(n2439) );
  NAND_GATE U3696 ( .I1(n2439), .I2(n2444), .O(n2452) );
  INV_GATE U3697 ( .I1(n2444), .O(n2442) );
  NAND_GATE U3698 ( .I1(n2445), .I2(n2442), .O(n2440) );
  NAND_GATE U3699 ( .I1(n2441), .I2(n2440), .O(n2450) );
  NAND_GATE U3700 ( .I1(n2443), .I2(n2442), .O(n2447) );
  NAND_GATE U3701 ( .I1(n2445), .I2(n2444), .O(n2446) );
  NAND3_GATE U3702 ( .I1(n2448), .I2(n2447), .I3(n2446), .O(n2449) );
  NAND_GATE U3703 ( .I1(n2450), .I2(n2449), .O(n2451) );
  NAND_GATE U3704 ( .I1(n2452), .I2(n2451), .O(n15308) );
  NAND_GATE U3705 ( .I1(n2453), .I2(n15308), .O(n2456) );
  INV_GATE U3706 ( .I1(n15308), .O(n2454) );
  NAND_GATE U3707 ( .I1(n15309), .I2(n2454), .O(n2455) );
  NAND_GATE U3708 ( .I1(n2456), .I2(n2455), .O(\A1[58] ) );
  OR_GATE U3709 ( .I1(n2457), .I2(n2462), .O(n2460) );
  OR_GATE U3710 ( .I1(n2461), .I2(n2458), .O(n2459) );
  AND_GATE U3711 ( .I1(n2460), .I2(n2459), .O(n2467) );
  NAND_GATE U3712 ( .I1(n2462), .I2(n1138), .O(n2464) );
  NAND3_GATE U3713 ( .I1(n2465), .I2(n2464), .I3(n2463), .O(n2466) );
  OR_GATE U3714 ( .I1(n2468), .I2(n2473), .O(n2471) );
  OR_GATE U3715 ( .I1(n2472), .I2(n2469), .O(n2470) );
  AND_GATE U3716 ( .I1(n2471), .I2(n2470), .O(n2478) );
  NAND_GATE U3717 ( .I1(n2473), .I2(n1137), .O(n2475) );
  NAND3_GATE U3718 ( .I1(n2476), .I2(n2475), .I3(n2474), .O(n2477) );
  NAND_GATE U3719 ( .I1(n2478), .I2(n2477), .O(n3340) );
  INV_GATE U3720 ( .I1(n3340), .O(n3343) );
  NAND_GATE U3721 ( .I1(B[27]), .I2(A[31]), .O(n3347) );
  INV_GATE U3722 ( .I1(n3347), .O(n3341) );
  NAND_GATE U3723 ( .I1(n3343), .I2(n3341), .O(n3338) );
  OR_GATE U3724 ( .I1(n2479), .I2(n2483), .O(n2482) );
  OR_GATE U3725 ( .I1(n2484), .I2(n2480), .O(n2481) );
  AND_GATE U3726 ( .I1(n2482), .I2(n2481), .O(n2489) );
  NAND_GATE U3727 ( .I1(n1136), .I2(n2484), .O(n2486) );
  NAND3_GATE U3728 ( .I1(n2487), .I2(n2486), .I3(n2485), .O(n2488) );
  NAND_GATE U3729 ( .I1(n2489), .I2(n2488), .O(n3324) );
  INV_GATE U3730 ( .I1(n3324), .O(n3327) );
  NAND_GATE U3731 ( .I1(B[27]), .I2(A[30]), .O(n3331) );
  INV_GATE U3732 ( .I1(n3331), .O(n3325) );
  NAND_GATE U3733 ( .I1(n3327), .I2(n3325), .O(n3322) );
  OR_GATE U3734 ( .I1(n2490), .I2(n2495), .O(n2493) );
  OR_GATE U3735 ( .I1(n2494), .I2(n2491), .O(n2492) );
  AND_GATE U3736 ( .I1(n2493), .I2(n2492), .O(n2500) );
  NAND_GATE U3737 ( .I1(n2495), .I2(n1134), .O(n2497) );
  NAND3_GATE U3738 ( .I1(n2498), .I2(n2497), .I3(n2496), .O(n2499) );
  NAND_GATE U3739 ( .I1(n2500), .I2(n2499), .O(n3308) );
  INV_GATE U3740 ( .I1(n3308), .O(n3311) );
  NAND_GATE U3741 ( .I1(B[27]), .I2(A[29]), .O(n3315) );
  INV_GATE U3742 ( .I1(n3315), .O(n3309) );
  NAND_GATE U3743 ( .I1(n3311), .I2(n3309), .O(n3306) );
  NAND_GATE U3744 ( .I1(B[27]), .I2(A[28]), .O(n3299) );
  INV_GATE U3745 ( .I1(n3299), .O(n3293) );
  OR_GATE U3746 ( .I1(n2501), .I2(n2506), .O(n2504) );
  OR_GATE U3747 ( .I1(n2505), .I2(n2502), .O(n2503) );
  AND_GATE U3748 ( .I1(n2504), .I2(n2503), .O(n2511) );
  NAND_GATE U3749 ( .I1(n2506), .I2(n1129), .O(n2508) );
  NAND3_GATE U3750 ( .I1(n2509), .I2(n2508), .I3(n2507), .O(n2510) );
  NAND_GATE U3751 ( .I1(n2511), .I2(n2510), .O(n3276) );
  INV_GATE U3752 ( .I1(n3276), .O(n3279) );
  NAND_GATE U3753 ( .I1(B[27]), .I2(A[27]), .O(n3283) );
  INV_GATE U3754 ( .I1(n3283), .O(n3277) );
  NAND_GATE U3755 ( .I1(n3279), .I2(n3277), .O(n3274) );
  OR_GATE U3756 ( .I1(n2512), .I2(n2517), .O(n2515) );
  OR_GATE U3757 ( .I1(n2516), .I2(n2513), .O(n2514) );
  AND_GATE U3758 ( .I1(n2515), .I2(n2514), .O(n2522) );
  NAND_GATE U3759 ( .I1(n2517), .I2(n1126), .O(n2519) );
  NAND3_GATE U3760 ( .I1(n2520), .I2(n2519), .I3(n2518), .O(n2521) );
  NAND_GATE U3761 ( .I1(n2522), .I2(n2521), .O(n2875) );
  INV_GATE U3762 ( .I1(n2875), .O(n2878) );
  NAND_GATE U3763 ( .I1(B[27]), .I2(A[26]), .O(n2882) );
  INV_GATE U3764 ( .I1(n2882), .O(n2876) );
  NAND_GATE U3765 ( .I1(n2878), .I2(n2876), .O(n2873) );
  OR_GATE U3766 ( .I1(n2523), .I2(n2528), .O(n2526) );
  OR_GATE U3767 ( .I1(n2527), .I2(n2524), .O(n2525) );
  AND_GATE U3768 ( .I1(n2526), .I2(n2525), .O(n2533) );
  NAND_GATE U3769 ( .I1(n2528), .I2(n1119), .O(n2530) );
  NAND3_GATE U3770 ( .I1(n2531), .I2(n2530), .I3(n2529), .O(n2532) );
  NAND_GATE U3771 ( .I1(n2533), .I2(n2532), .O(n3258) );
  INV_GATE U3772 ( .I1(n3258), .O(n3261) );
  NAND_GATE U3773 ( .I1(B[27]), .I2(A[25]), .O(n3265) );
  INV_GATE U3774 ( .I1(n3265), .O(n3259) );
  NAND_GATE U3775 ( .I1(n3261), .I2(n3259), .O(n3256) );
  OR_GATE U3776 ( .I1(n2534), .I2(n2539), .O(n2537) );
  OR_GATE U3777 ( .I1(n2538), .I2(n2535), .O(n2536) );
  AND_GATE U3778 ( .I1(n2537), .I2(n2536), .O(n2544) );
  NAND_GATE U3779 ( .I1(n2539), .I2(n1112), .O(n2541) );
  NAND3_GATE U3780 ( .I1(n2542), .I2(n2541), .I3(n2540), .O(n2543) );
  NAND_GATE U3781 ( .I1(n2544), .I2(n2543), .O(n3242) );
  INV_GATE U3782 ( .I1(n3242), .O(n3245) );
  NAND_GATE U3783 ( .I1(B[27]), .I2(A[24]), .O(n3249) );
  INV_GATE U3784 ( .I1(n3249), .O(n3243) );
  NAND_GATE U3785 ( .I1(n3245), .I2(n3243), .O(n3240) );
  OR_GATE U3786 ( .I1(n2545), .I2(n2550), .O(n2548) );
  OR_GATE U3787 ( .I1(n2549), .I2(n2546), .O(n2547) );
  AND_GATE U3788 ( .I1(n2548), .I2(n2547), .O(n2555) );
  NAND_GATE U3789 ( .I1(n2550), .I2(n1104), .O(n2552) );
  NAND3_GATE U3790 ( .I1(n2553), .I2(n2552), .I3(n2551), .O(n2554) );
  NAND_GATE U3791 ( .I1(n2555), .I2(n2554), .O(n3226) );
  INV_GATE U3792 ( .I1(n3226), .O(n3229) );
  NAND_GATE U3793 ( .I1(B[27]), .I2(A[23]), .O(n3233) );
  INV_GATE U3794 ( .I1(n3233), .O(n3227) );
  NAND_GATE U3795 ( .I1(n3229), .I2(n3227), .O(n3224) );
  OR_GATE U3796 ( .I1(n2556), .I2(n2562), .O(n2559) );
  OR_GATE U3797 ( .I1(n2563), .I2(n2557), .O(n2558) );
  AND_GATE U3798 ( .I1(n2559), .I2(n2558), .O(n2569) );
  OR_GATE U3799 ( .I1(n2563), .I2(n2560), .O(n2567) );
  NAND_GATE U3800 ( .I1(n2561), .I2(n1097), .O(n2566) );
  NAND4_GATE U3801 ( .I1(n2567), .I2(n2566), .I3(n2565), .I4(n2564), .O(n2568)
         );
  NAND_GATE U3802 ( .I1(n2569), .I2(n2568), .O(n3210) );
  INV_GATE U3803 ( .I1(n3210), .O(n3213) );
  NAND_GATE U3804 ( .I1(B[27]), .I2(A[22]), .O(n3217) );
  INV_GATE U3805 ( .I1(n3217), .O(n3211) );
  NAND_GATE U3806 ( .I1(n3213), .I2(n3211), .O(n3207) );
  OR_GATE U3807 ( .I1(n2570), .I2(n2576), .O(n2573) );
  OR_GATE U3808 ( .I1(n2577), .I2(n2571), .O(n2572) );
  AND_GATE U3809 ( .I1(n2573), .I2(n2572), .O(n2583) );
  OR_GATE U3810 ( .I1(n2577), .I2(n2574), .O(n2581) );
  NAND_GATE U3811 ( .I1(n2575), .I2(n1088), .O(n2580) );
  NAND4_GATE U3812 ( .I1(n2581), .I2(n2580), .I3(n2579), .I4(n2578), .O(n2582)
         );
  NAND_GATE U3813 ( .I1(n2583), .I2(n2582), .O(n3193) );
  INV_GATE U3814 ( .I1(n3193), .O(n3196) );
  NAND_GATE U3815 ( .I1(B[27]), .I2(A[21]), .O(n3200) );
  INV_GATE U3816 ( .I1(n3200), .O(n3194) );
  NAND_GATE U3817 ( .I1(n3196), .I2(n3194), .O(n3190) );
  OR_GATE U3818 ( .I1(n2584), .I2(n2590), .O(n2587) );
  OR_GATE U3819 ( .I1(n2591), .I2(n2585), .O(n2586) );
  AND_GATE U3820 ( .I1(n2587), .I2(n2586), .O(n2597) );
  OR_GATE U3821 ( .I1(n2591), .I2(n2588), .O(n2595) );
  NAND_GATE U3822 ( .I1(n2589), .I2(n1095), .O(n2594) );
  NAND4_GATE U3823 ( .I1(n2595), .I2(n2594), .I3(n2593), .I4(n2592), .O(n2596)
         );
  NAND_GATE U3824 ( .I1(n2597), .I2(n2596), .O(n3176) );
  INV_GATE U3825 ( .I1(n3176), .O(n3179) );
  NAND_GATE U3826 ( .I1(B[27]), .I2(A[20]), .O(n3183) );
  INV_GATE U3827 ( .I1(n3183), .O(n3177) );
  NAND_GATE U3828 ( .I1(n3179), .I2(n3177), .O(n3173) );
  OR_GATE U3829 ( .I1(n2598), .I2(n2603), .O(n2601) );
  OR_GATE U3830 ( .I1(n2602), .I2(n2599), .O(n2600) );
  AND_GATE U3831 ( .I1(n2601), .I2(n2600), .O(n2608) );
  NAND_GATE U3832 ( .I1(n2603), .I2(n1096), .O(n2605) );
  NAND3_GATE U3833 ( .I1(n2606), .I2(n2605), .I3(n2604), .O(n2607) );
  NAND_GATE U3834 ( .I1(n2608), .I2(n2607), .O(n3159) );
  INV_GATE U3835 ( .I1(n3159), .O(n3162) );
  NAND_GATE U3836 ( .I1(B[27]), .I2(A[19]), .O(n3166) );
  INV_GATE U3837 ( .I1(n3166), .O(n3160) );
  NAND_GATE U3838 ( .I1(n3162), .I2(n3160), .O(n3157) );
  OR_GATE U3839 ( .I1(n2609), .I2(n2614), .O(n2612) );
  OR_GATE U3840 ( .I1(n2613), .I2(n2610), .O(n2611) );
  AND_GATE U3841 ( .I1(n2612), .I2(n2611), .O(n2619) );
  NAND_GATE U3842 ( .I1(n2614), .I2(n1090), .O(n2616) );
  NAND3_GATE U3843 ( .I1(n2617), .I2(n2616), .I3(n2615), .O(n2618) );
  NAND_GATE U3844 ( .I1(n2619), .I2(n2618), .O(n3143) );
  INV_GATE U3845 ( .I1(n3143), .O(n3146) );
  NAND_GATE U3846 ( .I1(B[27]), .I2(A[18]), .O(n3150) );
  INV_GATE U3847 ( .I1(n3150), .O(n3144) );
  NAND_GATE U3848 ( .I1(n3146), .I2(n3144), .O(n3141) );
  OR_GATE U3849 ( .I1(n2620), .I2(n2625), .O(n2623) );
  OR_GATE U3850 ( .I1(n2624), .I2(n2621), .O(n2622) );
  AND_GATE U3851 ( .I1(n2623), .I2(n2622), .O(n2630) );
  NAND_GATE U3852 ( .I1(n2625), .I2(n1083), .O(n2627) );
  NAND3_GATE U3853 ( .I1(n2628), .I2(n2627), .I3(n2626), .O(n2629) );
  NAND_GATE U3854 ( .I1(n2630), .I2(n2629), .O(n3127) );
  INV_GATE U3855 ( .I1(n3127), .O(n3130) );
  NAND_GATE U3856 ( .I1(B[27]), .I2(A[17]), .O(n3134) );
  INV_GATE U3857 ( .I1(n3134), .O(n3128) );
  NAND_GATE U3858 ( .I1(n3130), .I2(n3128), .O(n3125) );
  OR_GATE U3859 ( .I1(n2631), .I2(n2636), .O(n2634) );
  OR_GATE U3860 ( .I1(n2635), .I2(n2632), .O(n2633) );
  AND_GATE U3861 ( .I1(n2634), .I2(n2633), .O(n2641) );
  NAND_GATE U3862 ( .I1(n2636), .I2(n1082), .O(n2638) );
  NAND3_GATE U3863 ( .I1(n2639), .I2(n2638), .I3(n2637), .O(n2640) );
  NAND_GATE U3864 ( .I1(n2641), .I2(n2640), .O(n3111) );
  INV_GATE U3865 ( .I1(n3111), .O(n3114) );
  NAND_GATE U3866 ( .I1(B[27]), .I2(A[16]), .O(n3118) );
  INV_GATE U3867 ( .I1(n3118), .O(n3112) );
  NAND_GATE U3868 ( .I1(n3114), .I2(n3112), .O(n3109) );
  OR_GATE U3869 ( .I1(n2642), .I2(n2647), .O(n2645) );
  OR_GATE U3870 ( .I1(n2646), .I2(n2643), .O(n2644) );
  AND_GATE U3871 ( .I1(n2645), .I2(n2644), .O(n2652) );
  NAND_GATE U3872 ( .I1(n2647), .I2(n1081), .O(n2649) );
  NAND3_GATE U3873 ( .I1(n2650), .I2(n2649), .I3(n2648), .O(n2651) );
  NAND_GATE U3874 ( .I1(n2652), .I2(n2651), .O(n3095) );
  INV_GATE U3875 ( .I1(n3095), .O(n3098) );
  NAND_GATE U3876 ( .I1(B[27]), .I2(A[15]), .O(n3102) );
  INV_GATE U3877 ( .I1(n3102), .O(n3096) );
  NAND_GATE U3878 ( .I1(n3098), .I2(n3096), .O(n3093) );
  OR_GATE U3879 ( .I1(n2653), .I2(n2658), .O(n2656) );
  OR_GATE U3880 ( .I1(n2657), .I2(n2654), .O(n2655) );
  AND_GATE U3881 ( .I1(n2656), .I2(n2655), .O(n2663) );
  NAND_GATE U3882 ( .I1(n2658), .I2(n1080), .O(n2660) );
  NAND3_GATE U3883 ( .I1(n2661), .I2(n2660), .I3(n2659), .O(n2662) );
  NAND_GATE U3884 ( .I1(n2663), .I2(n2662), .O(n3083) );
  INV_GATE U3885 ( .I1(n3083), .O(n3081) );
  NAND_GATE U3886 ( .I1(B[27]), .I2(A[14]), .O(n3086) );
  INV_GATE U3887 ( .I1(n3086), .O(n3079) );
  NAND_GATE U3888 ( .I1(n3081), .I2(n3079), .O(n3076) );
  OR_GATE U3889 ( .I1(n2664), .I2(n2669), .O(n2667) );
  OR_GATE U3890 ( .I1(n2668), .I2(n2665), .O(n2666) );
  AND_GATE U3891 ( .I1(n2667), .I2(n2666), .O(n2674) );
  NAND_GATE U3892 ( .I1(n2669), .I2(n1078), .O(n2671) );
  NAND3_GATE U3893 ( .I1(n2672), .I2(n2671), .I3(n2670), .O(n2673) );
  NAND_GATE U3894 ( .I1(n2674), .I2(n2673), .O(n3066) );
  INV_GATE U3895 ( .I1(n3066), .O(n3065) );
  NAND_GATE U3896 ( .I1(B[27]), .I2(A[13]), .O(n3069) );
  INV_GATE U3897 ( .I1(n3069), .O(n3063) );
  NAND_GATE U3898 ( .I1(n3065), .I2(n3063), .O(n3060) );
  INV_GATE U3899 ( .I1(n2675), .O(n2679) );
  NAND_GATE U3900 ( .I1(n2679), .I2(n2680), .O(n2677) );
  NAND_GATE U3901 ( .I1(n2675), .I2(n800), .O(n2676) );
  NAND3_GATE U3902 ( .I1(n2678), .I2(n2677), .I3(n2676), .O(n2683) );
  NAND3_GATE U3903 ( .I1(n2681), .I2(n2680), .I3(n2679), .O(n2682) );
  NAND_GATE U3904 ( .I1(n2683), .I2(n2682), .O(n2686) );
  INV_GATE U3905 ( .I1(n2684), .O(n2685) );
  NAND_GATE U3906 ( .I1(B[27]), .I2(A[12]), .O(n3053) );
  INV_GATE U3907 ( .I1(n3053), .O(n3047) );
  NAND_GATE U3908 ( .I1(n1309), .I2(n3047), .O(n3048) );
  NAND_GATE U3909 ( .I1(n2686), .I2(n3053), .O(n2820) );
  NAND_GATE U3910 ( .I1(n280), .I2(n3053), .O(n2819) );
  INV_GATE U3911 ( .I1(n2692), .O(n2690) );
  NAND3_GATE U3912 ( .I1(n2687), .I2(n2690), .I3(n2689), .O(n2698) );
  INV_GATE U3913 ( .I1(n2689), .O(n2691) );
  NAND_GATE U3914 ( .I1(n2688), .I2(n2691), .O(n2697) );
  NAND_GATE U3915 ( .I1(n2690), .I2(n2689), .O(n2694) );
  NAND_GATE U3916 ( .I1(n2692), .I2(n2691), .O(n2693) );
  NAND3_GATE U3917 ( .I1(n2695), .I2(n2694), .I3(n2693), .O(n2696) );
  NAND3_GATE U3918 ( .I1(n2698), .I2(n2697), .I3(n2696), .O(n2894) );
  NAND_GATE U3919 ( .I1(B[27]), .I2(A[11]), .O(n2892) );
  INV_GATE U3920 ( .I1(n2892), .O(n2890) );
  NAND_GATE U3921 ( .I1(n224), .I2(n2890), .O(n2887) );
  INV_GATE U3922 ( .I1(n2699), .O(n2704) );
  NAND_GATE U3923 ( .I1(n2704), .I2(n2706), .O(n2701) );
  NAND3_GATE U3924 ( .I1(n2702), .I2(n2701), .I3(n2700), .O(n2709) );
  OR_GATE U3925 ( .I1(n2706), .I2(n2703), .O(n2708) );
  NAND3_GATE U3926 ( .I1(n2706), .I2(n2705), .I3(n2704), .O(n2707) );
  NAND3_GATE U3927 ( .I1(n2709), .I2(n2708), .I3(n2707), .O(n3030) );
  INV_GATE U3928 ( .I1(n3030), .O(n3028) );
  NAND_GATE U3929 ( .I1(B[27]), .I2(A[10]), .O(n3031) );
  INV_GATE U3930 ( .I1(n3031), .O(n3026) );
  NAND_GATE U3931 ( .I1(n3028), .I2(n3026), .O(n3027) );
  NAND_GATE U3932 ( .I1(n274), .I2(n2716), .O(n2712) );
  NAND3_GATE U3933 ( .I1(n2713), .I2(n2712), .I3(n2711), .O(n2719) );
  OR_GATE U3934 ( .I1(n2716), .I2(n2714), .O(n2718) );
  NAND3_GATE U3935 ( .I1(n2716), .I2(n2715), .I3(n274), .O(n2717) );
  NAND3_GATE U3936 ( .I1(n2719), .I2(n2718), .I3(n2717), .O(n3013) );
  NAND_GATE U3937 ( .I1(B[27]), .I2(A[9]), .O(n3012) );
  INV_GATE U3938 ( .I1(n3012), .O(n3020) );
  NAND_GATE U3939 ( .I1(n273), .I2(n3020), .O(n3011) );
  NAND_GATE U3940 ( .I1(n804), .I2(n2726), .O(n2722) );
  NAND3_GATE U3941 ( .I1(n2723), .I2(n2722), .I3(n2721), .O(n2729) );
  OR_GATE U3942 ( .I1(n2726), .I2(n2724), .O(n2728) );
  NAND3_GATE U3943 ( .I1(n804), .I2(n2726), .I3(n2725), .O(n2727) );
  NAND3_GATE U3944 ( .I1(n2729), .I2(n2728), .I3(n2727), .O(n2999) );
  NAND_GATE U3945 ( .I1(B[27]), .I2(A[8]), .O(n2998) );
  INV_GATE U3946 ( .I1(n2998), .O(n3006) );
  NAND_GATE U3947 ( .I1(n871), .I2(n3006), .O(n2996) );
  NAND_GATE U3948 ( .I1(B[27]), .I2(A[7]), .O(n2987) );
  INV_GATE U3949 ( .I1(n2987), .O(n3685) );
  OR_GATE U3950 ( .I1(n2734), .I2(n2730), .O(n2733) );
  NAND3_GATE U3951 ( .I1(n2731), .I2(n2735), .I3(n2734), .O(n2732) );
  AND_GATE U3952 ( .I1(n2733), .I2(n2732), .O(n2740) );
  NAND_GATE U3953 ( .I1(n2735), .I2(n2734), .O(n2736) );
  NAND3_GATE U3954 ( .I1(n2738), .I2(n2737), .I3(n2736), .O(n2739) );
  NAND_GATE U3955 ( .I1(n2740), .I2(n2739), .O(n2986) );
  INV_GATE U3956 ( .I1(n2986), .O(n2988) );
  NAND_GATE U3957 ( .I1(n3685), .I2(n2988), .O(n2990) );
  OR_GATE U3958 ( .I1(n2751), .I2(n2741), .O(n2757) );
  INV_GATE U3959 ( .I1(n2742), .O(n2793) );
  NAND_GATE U3960 ( .I1(n2745), .I2(n2793), .O(n2747) );
  NAND4_GATE U3961 ( .I1(n2745), .I2(n2744), .I3(n2743), .I4(n2794), .O(n2746)
         );
  NAND_GATE U3962 ( .I1(n2747), .I2(n2746), .O(n2748) );
  NAND_GATE U3963 ( .I1(n2750), .I2(n2748), .O(n2756) );
  NAND_GATE U3964 ( .I1(n2751), .I2(n2750), .O(n2752) );
  NAND3_GATE U3965 ( .I1(n2754), .I2(n2753), .I3(n2752), .O(n2755) );
  NAND3_GATE U3966 ( .I1(n2757), .I2(n2756), .I3(n2755), .O(n2976) );
  NAND_GATE U3967 ( .I1(B[27]), .I2(A[6]), .O(n2971) );
  INV_GATE U3968 ( .I1(n2971), .O(n2979) );
  NAND_GATE U3969 ( .I1(B[27]), .I2(A[5]), .O(n2909) );
  INV_GATE U3970 ( .I1(n2909), .O(n2901) );
  NAND3_GATE U3971 ( .I1(n2759), .I2(n2758), .I3(n2764), .O(n2760) );
  NAND_GATE U3972 ( .I1(n2761), .I2(n2760), .O(n2933) );
  INV_GATE U3973 ( .I1(n2933), .O(n2762) );
  NAND3_GATE U3974 ( .I1(n2767), .I2(n2761), .I3(n2765), .O(n2936) );
  NAND_GATE U3975 ( .I1(n2762), .I2(n2936), .O(n2777) );
  NAND3_GATE U3976 ( .I1(n2764), .I2(n2766), .I3(n2763), .O(n2769) );
  NAND3_GATE U3977 ( .I1(n2767), .I2(n2766), .I3(n2765), .O(n2768) );
  AND_GATE U3978 ( .I1(n2769), .I2(n2768), .O(n2934) );
  NAND3_GATE U3979 ( .I1(B[27]), .I2(B[28]), .I3(n1196), .O(n2916) );
  INV_GATE U3980 ( .I1(n2916), .O(n2919) );
  NAND_GATE U3981 ( .I1(n1395), .I2(A[1]), .O(n2770) );
  NAND_GATE U3982 ( .I1(n14784), .I2(n2770), .O(n2771) );
  NAND_GATE U3983 ( .I1(B[28]), .I2(n2771), .O(n2910) );
  NAND_GATE U3984 ( .I1(n1394), .I2(A[0]), .O(n2772) );
  NAND_GATE U3985 ( .I1(n14781), .I2(n2772), .O(n2773) );
  NAND_GATE U3986 ( .I1(B[29]), .I2(n2773), .O(n2911) );
  NAND_GATE U3987 ( .I1(n2910), .I2(n2911), .O(n2917) );
  NAND_GATE U3988 ( .I1(B[27]), .I2(A[2]), .O(n2918) );
  NAND_GATE U3989 ( .I1(n2915), .I2(n2918), .O(n2774) );
  NAND_GATE U3990 ( .I1(n2919), .I2(n2774), .O(n2776) );
  INV_GATE U3991 ( .I1(n2918), .O(n2913) );
  NAND_GATE U3992 ( .I1(n2917), .I2(n2913), .O(n2775) );
  NAND_GATE U3993 ( .I1(n2776), .I2(n2775), .O(n2940) );
  NAND3_GATE U3994 ( .I1(n2777), .I2(n2934), .I3(n2940), .O(n2779) );
  NAND_GATE U3995 ( .I1(B[27]), .I2(A[3]), .O(n2943) );
  INV_GATE U3996 ( .I1(n2943), .O(n2932) );
  NAND3_GATE U3997 ( .I1(n2932), .I2(n2933), .I3(n2934), .O(n2778) );
  NAND_GATE U3998 ( .I1(n2932), .I2(n2940), .O(n2937) );
  NAND3_GATE U3999 ( .I1(n2779), .I2(n2778), .I3(n2937), .O(n2954) );
  NAND_GATE U4000 ( .I1(B[27]), .I2(A[4]), .O(n2953) );
  OR_GATE U4001 ( .I1(n2786), .I2(n2780), .O(n2784) );
  NAND4_GATE U4002 ( .I1(n2782), .I2(n1194), .I3(n2781), .I4(n1193), .O(n2783)
         );
  AND_GATE U4003 ( .I1(n2784), .I2(n2783), .O(n2950) );
  NAND_GATE U4004 ( .I1(n1193), .I2(n2786), .O(n2788) );
  NAND3_GATE U4005 ( .I1(n2789), .I2(n2788), .I3(n2787), .O(n2951) );
  NAND_GATE U4006 ( .I1(n2953), .I2(n2960), .O(n2790) );
  NAND_GATE U4007 ( .I1(n2954), .I2(n2790), .O(n2792) );
  INV_GATE U4008 ( .I1(n2953), .O(n2963) );
  INV_GATE U4009 ( .I1(n2960), .O(n2952) );
  NAND_GATE U4010 ( .I1(n2963), .I2(n2952), .O(n2791) );
  NAND_GATE U4011 ( .I1(n2792), .I2(n2791), .O(n2906) );
  NAND_GATE U4012 ( .I1(n2901), .I2(n2906), .O(n2900) );
  INV_GATE U4013 ( .I1(n2794), .O(n2796) );
  NAND_GATE U4014 ( .I1(n2793), .I2(n2794), .O(n2804) );
  NAND3_GATE U4015 ( .I1(n2798), .I2(n2804), .I3(n2799), .O(n2902) );
  NAND3_GATE U4016 ( .I1(n2794), .I2(n185), .I3(n2795), .O(n2800) );
  NAND3_GATE U4017 ( .I1(n2797), .I2(n2796), .I3(n2795), .O(n2801) );
  NAND3_GATE U4018 ( .I1(n2901), .I2(n2902), .I3(n1143), .O(n2806) );
  NAND_GATE U4019 ( .I1(n2799), .I2(n2798), .O(n2802) );
  NAND3_GATE U4020 ( .I1(n2802), .I2(n2801), .I3(n2800), .O(n2803) );
  NAND_GATE U4021 ( .I1(n2804), .I2(n2803), .O(n2905) );
  NAND_GATE U4022 ( .I1(n2906), .I2(n2905), .O(n2805) );
  NAND3_GATE U4023 ( .I1(n2900), .I2(n2806), .I3(n2805), .O(n2970) );
  NAND_GATE U4024 ( .I1(n2976), .I2(n2971), .O(n2807) );
  NAND_GATE U4025 ( .I1(n2970), .I2(n2807), .O(n2808) );
  NAND_GATE U4026 ( .I1(n2987), .I2(n2986), .O(n2809) );
  NAND_GATE U4027 ( .I1(n2991), .I2(n2809), .O(n2810) );
  NAND_GATE U4028 ( .I1(n2990), .I2(n2810), .O(n2997) );
  NAND_GATE U4029 ( .I1(n2999), .I2(n2998), .O(n2811) );
  NAND_GATE U4030 ( .I1(n2997), .I2(n2811), .O(n2812) );
  NAND_GATE U4031 ( .I1(n3013), .I2(n3012), .O(n2813) );
  NAND_GATE U4032 ( .I1(n781), .I2(n2813), .O(n2814) );
  NAND_GATE U4033 ( .I1(n3011), .I2(n2814), .O(n3029) );
  NAND_GATE U4034 ( .I1(n3030), .I2(n3031), .O(n2815) );
  NAND_GATE U4035 ( .I1(n3029), .I2(n2815), .O(n2816) );
  NAND_GATE U4036 ( .I1(n3027), .I2(n2816), .O(n2891) );
  NAND_GATE U4037 ( .I1(n2894), .I2(n2892), .O(n2817) );
  NAND_GATE U4038 ( .I1(n2891), .I2(n2817), .O(n2818) );
  NAND_GATE U4039 ( .I1(n2887), .I2(n2818), .O(n3049) );
  NAND3_GATE U4040 ( .I1(n2820), .I2(n2819), .I3(n3049), .O(n2821) );
  NAND_GATE U4041 ( .I1(n3048), .I2(n2821), .O(n3064) );
  NAND_GATE U4042 ( .I1(n3066), .I2(n3069), .O(n2822) );
  NAND_GATE U4043 ( .I1(n3064), .I2(n2822), .O(n2823) );
  NAND_GATE U4044 ( .I1(n3060), .I2(n2823), .O(n3080) );
  NAND_GATE U4045 ( .I1(n3083), .I2(n3086), .O(n2824) );
  NAND_GATE U4046 ( .I1(n3080), .I2(n2824), .O(n2825) );
  NAND_GATE U4047 ( .I1(n3076), .I2(n2825), .O(n3097) );
  NAND_GATE U4048 ( .I1(n3095), .I2(n3102), .O(n2826) );
  NAND_GATE U4049 ( .I1(n3097), .I2(n2826), .O(n2827) );
  NAND_GATE U4050 ( .I1(n3093), .I2(n2827), .O(n3113) );
  NAND_GATE U4051 ( .I1(n3111), .I2(n3118), .O(n2828) );
  NAND_GATE U4052 ( .I1(n3113), .I2(n2828), .O(n2829) );
  NAND_GATE U4053 ( .I1(n3109), .I2(n2829), .O(n3129) );
  NAND_GATE U4054 ( .I1(n3127), .I2(n3134), .O(n2830) );
  NAND_GATE U4055 ( .I1(n3129), .I2(n2830), .O(n2831) );
  NAND_GATE U4056 ( .I1(n3125), .I2(n2831), .O(n3145) );
  NAND_GATE U4057 ( .I1(n3143), .I2(n3150), .O(n2832) );
  NAND_GATE U4058 ( .I1(n3145), .I2(n2832), .O(n2833) );
  NAND_GATE U4059 ( .I1(n3141), .I2(n2833), .O(n3161) );
  NAND_GATE U4060 ( .I1(n3159), .I2(n3166), .O(n2834) );
  NAND_GATE U4061 ( .I1(n3161), .I2(n2834), .O(n2835) );
  NAND_GATE U4062 ( .I1(n3157), .I2(n2835), .O(n3178) );
  NAND_GATE U4063 ( .I1(n3176), .I2(n3183), .O(n2836) );
  NAND_GATE U4064 ( .I1(n3178), .I2(n2836), .O(n2837) );
  NAND_GATE U4065 ( .I1(n3173), .I2(n2837), .O(n3195) );
  NAND_GATE U4066 ( .I1(n3193), .I2(n3200), .O(n2838) );
  NAND_GATE U4067 ( .I1(n3195), .I2(n2838), .O(n2839) );
  NAND_GATE U4068 ( .I1(n3190), .I2(n2839), .O(n3212) );
  NAND_GATE U4069 ( .I1(n3210), .I2(n3217), .O(n2840) );
  NAND_GATE U4070 ( .I1(n3212), .I2(n2840), .O(n2841) );
  NAND_GATE U4071 ( .I1(n3207), .I2(n2841), .O(n3228) );
  NAND_GATE U4072 ( .I1(n3226), .I2(n3233), .O(n2842) );
  NAND_GATE U4073 ( .I1(n3228), .I2(n2842), .O(n2843) );
  NAND_GATE U4074 ( .I1(n3224), .I2(n2843), .O(n3244) );
  NAND_GATE U4075 ( .I1(n3242), .I2(n3249), .O(n2844) );
  NAND_GATE U4076 ( .I1(n3244), .I2(n2844), .O(n2845) );
  NAND_GATE U4077 ( .I1(n3240), .I2(n2845), .O(n3260) );
  NAND_GATE U4078 ( .I1(n3258), .I2(n3265), .O(n2846) );
  NAND_GATE U4079 ( .I1(n3260), .I2(n2846), .O(n2847) );
  NAND_GATE U4080 ( .I1(n3256), .I2(n2847), .O(n2877) );
  NAND_GATE U4081 ( .I1(n2875), .I2(n2882), .O(n2848) );
  NAND_GATE U4082 ( .I1(n2877), .I2(n2848), .O(n2849) );
  NAND_GATE U4083 ( .I1(n2873), .I2(n2849), .O(n3278) );
  NAND_GATE U4084 ( .I1(n3276), .I2(n3283), .O(n2850) );
  NAND_GATE U4085 ( .I1(n3278), .I2(n2850), .O(n2851) );
  NAND_GATE U4086 ( .I1(n3274), .I2(n2851), .O(n3295) );
  NAND_GATE U4087 ( .I1(n3293), .I2(n3295), .O(n3290) );
  OR_GATE U4088 ( .I1(n2852), .I2(n2857), .O(n2855) );
  OR_GATE U4089 ( .I1(n2856), .I2(n2853), .O(n2854) );
  AND_GATE U4090 ( .I1(n2855), .I2(n2854), .O(n2862) );
  NAND_GATE U4091 ( .I1(n2857), .I2(n1132), .O(n2859) );
  NAND3_GATE U4092 ( .I1(n2860), .I2(n2859), .I3(n2858), .O(n2861) );
  NAND_GATE U4093 ( .I1(n2862), .I2(n2861), .O(n3291) );
  INV_GATE U4094 ( .I1(n3291), .O(n3294) );
  INV_GATE U4095 ( .I1(n3295), .O(n3292) );
  NAND_GATE U4096 ( .I1(n3299), .I2(n3292), .O(n2863) );
  NAND_GATE U4097 ( .I1(n3294), .I2(n2863), .O(n2864) );
  NAND_GATE U4098 ( .I1(n3290), .I2(n2864), .O(n3310) );
  NAND_GATE U4099 ( .I1(n3308), .I2(n3315), .O(n2865) );
  NAND_GATE U4100 ( .I1(n3310), .I2(n2865), .O(n2866) );
  NAND_GATE U4101 ( .I1(n3306), .I2(n2866), .O(n3326) );
  NAND_GATE U4102 ( .I1(n3324), .I2(n3331), .O(n2867) );
  NAND_GATE U4103 ( .I1(n3326), .I2(n2867), .O(n2868) );
  NAND_GATE U4104 ( .I1(n3322), .I2(n2868), .O(n3342) );
  NAND_GATE U4105 ( .I1(n3340), .I2(n3347), .O(n2869) );
  NAND_GATE U4106 ( .I1(n3342), .I2(n2869), .O(n2870) );
  NAND_GATE U4107 ( .I1(n3338), .I2(n2870), .O(n2871) );
  NAND_GATE U4108 ( .I1(n288), .I2(n2871), .O(n15310) );
  AND_GATE U4109 ( .I1(n15310), .I2(n2872), .O(\A1[57] ) );
  NAND_GATE U4110 ( .I1(B[26]), .I2(A[31]), .O(n3362) );
  INV_GATE U4111 ( .I1(n3362), .O(n3336) );
  NAND_GATE U4112 ( .I1(B[26]), .I2(A[30]), .O(n3373) );
  INV_GATE U4113 ( .I1(n3373), .O(n3320) );
  NAND_GATE U4114 ( .I1(B[26]), .I2(A[29]), .O(n3384) );
  INV_GATE U4115 ( .I1(n3384), .O(n3304) );
  NAND_GATE U4116 ( .I1(B[26]), .I2(A[28]), .O(n3395) );
  INV_GATE U4117 ( .I1(n3395), .O(n3288) );
  NAND_GATE U4118 ( .I1(B[26]), .I2(A[27]), .O(n3406) );
  INV_GATE U4119 ( .I1(n3406), .O(n3272) );
  INV_GATE U4120 ( .I1(n2873), .O(n2874) );
  NAND_GATE U4121 ( .I1(n2874), .I2(n2877), .O(n2886) );
  NAND_GATE U4122 ( .I1(n2876), .I2(n2880), .O(n2884) );
  NAND_GATE U4123 ( .I1(n2878), .I2(n2877), .O(n2879) );
  NAND_GATE U4124 ( .I1(n2880), .I2(n2879), .O(n2881) );
  NAND_GATE U4125 ( .I1(n2882), .I2(n2881), .O(n2883) );
  NAND_GATE U4126 ( .I1(n2884), .I2(n2883), .O(n2885) );
  NAND_GATE U4127 ( .I1(n2886), .I2(n2885), .O(n3404) );
  NAND_GATE U4128 ( .I1(n3272), .I2(n3404), .O(n3401) );
  NAND_GATE U4129 ( .I1(B[26]), .I2(A[26]), .O(n3417) );
  INV_GATE U4130 ( .I1(n3417), .O(n3270) );
  NAND_GATE U4131 ( .I1(B[26]), .I2(A[25]), .O(n3753) );
  INV_GATE U4132 ( .I1(n3753), .O(n3254) );
  NAND_GATE U4133 ( .I1(B[26]), .I2(A[24]), .O(n3428) );
  INV_GATE U4134 ( .I1(n3428), .O(n3238) );
  NAND_GATE U4135 ( .I1(B[26]), .I2(A[23]), .O(n3439) );
  INV_GATE U4136 ( .I1(n3439), .O(n3222) );
  NAND_GATE U4137 ( .I1(B[26]), .I2(A[22]), .O(n3450) );
  INV_GATE U4138 ( .I1(n3450), .O(n3205) );
  NAND_GATE U4139 ( .I1(B[26]), .I2(A[21]), .O(n3461) );
  INV_GATE U4140 ( .I1(n3461), .O(n3188) );
  NAND_GATE U4141 ( .I1(B[26]), .I2(A[20]), .O(n3472) );
  INV_GATE U4142 ( .I1(n3472), .O(n3171) );
  NAND_GATE U4143 ( .I1(B[26]), .I2(A[19]), .O(n3483) );
  INV_GATE U4144 ( .I1(n3483), .O(n3155) );
  NAND_GATE U4145 ( .I1(B[26]), .I2(A[18]), .O(n3494) );
  INV_GATE U4146 ( .I1(n3494), .O(n3139) );
  NAND_GATE U4147 ( .I1(B[26]), .I2(A[17]), .O(n3505) );
  INV_GATE U4148 ( .I1(n3505), .O(n3123) );
  NAND_GATE U4149 ( .I1(B[26]), .I2(A[16]), .O(n3516) );
  INV_GATE U4150 ( .I1(n3516), .O(n3107) );
  NAND_GATE U4151 ( .I1(B[26]), .I2(A[15]), .O(n3527) );
  INV_GATE U4152 ( .I1(n3527), .O(n3091) );
  NAND_GATE U4153 ( .I1(B[26]), .I2(A[14]), .O(n3538) );
  INV_GATE U4154 ( .I1(n3538), .O(n3074) );
  INV_GATE U4155 ( .I1(n2887), .O(n2888) );
  NAND_GATE U4156 ( .I1(n2888), .I2(n2891), .O(n2899) );
  INV_GATE U4157 ( .I1(n2891), .O(n2893) );
  NAND_GATE U4158 ( .I1(n2894), .I2(n2893), .O(n2889) );
  NAND_GATE U4159 ( .I1(n2890), .I2(n2889), .O(n2897) );
  NAND_GATE U4160 ( .I1(n224), .I2(n2891), .O(n2896) );
  NAND3_GATE U4161 ( .I1(n2894), .I2(n2893), .I3(n2892), .O(n2895) );
  NAND3_GATE U4162 ( .I1(n2897), .I2(n2896), .I3(n2895), .O(n2898) );
  NAND_GATE U4163 ( .I1(n2899), .I2(n2898), .O(n3557) );
  NAND_GATE U4164 ( .I1(B[26]), .I2(A[11]), .O(n3564) );
  INV_GATE U4165 ( .I1(n3564), .O(n3034) );
  NAND_GATE U4166 ( .I1(B[26]), .I2(A[6]), .O(n3591) );
  INV_GATE U4167 ( .I1(n3591), .O(n3811) );
  OR_GATE U4168 ( .I1(n2905), .I2(n2900), .O(n2904) );
  NAND4_GATE U4169 ( .I1(n2902), .I2(n1143), .I3(n2901), .I4(n215), .O(n2903)
         );
  NAND_GATE U4170 ( .I1(n215), .I2(n2905), .O(n2908) );
  NAND3_GATE U4171 ( .I1(n2908), .I2(n2907), .I3(n2909), .O(n3661) );
  NAND_GATE U4172 ( .I1(n861), .I2(n3661), .O(n3657) );
  NAND4_GATE U4173 ( .I1(n2909), .I2(n3591), .I3(n2908), .I4(n2907), .O(n2967)
         );
  NAND_GATE U4174 ( .I1(n3591), .I2(n749), .O(n2966) );
  NAND3_GATE U4175 ( .I1(n2911), .I2(n2910), .I3(n2916), .O(n2912) );
  NAND_GATE U4176 ( .I1(n2913), .I2(n2912), .O(n3614) );
  INV_GATE U4177 ( .I1(n3614), .O(n2914) );
  NAND3_GATE U4178 ( .I1(n2917), .I2(n2913), .I3(n2919), .O(n3617) );
  NAND_GATE U4179 ( .I1(n2914), .I2(n3617), .O(n2929) );
  NAND3_GATE U4180 ( .I1(n2916), .I2(n2918), .I3(n2915), .O(n2921) );
  NAND3_GATE U4181 ( .I1(n2919), .I2(n2918), .I3(n2917), .O(n2920) );
  AND_GATE U4182 ( .I1(n2921), .I2(n2920), .O(n3615) );
  NAND3_GATE U4183 ( .I1(B[26]), .I2(B[27]), .I3(n1196), .O(n3600) );
  INV_GATE U4184 ( .I1(n3600), .O(n3598) );
  NAND_GATE U4185 ( .I1(n1393), .I2(A[0]), .O(n2922) );
  NAND_GATE U4186 ( .I1(n14781), .I2(n2922), .O(n2923) );
  NAND_GATE U4187 ( .I1(B[28]), .I2(n2923), .O(n3592) );
  NAND_GATE U4188 ( .I1(n1394), .I2(A[1]), .O(n2924) );
  NAND_GATE U4189 ( .I1(n14784), .I2(n2924), .O(n2925) );
  NAND_GATE U4190 ( .I1(B[27]), .I2(n2925), .O(n3593) );
  NAND_GATE U4191 ( .I1(n3592), .I2(n3593), .O(n3597) );
  NAND_GATE U4192 ( .I1(B[26]), .I2(A[2]), .O(n3599) );
  NAND_GATE U4193 ( .I1(n744), .I2(n3599), .O(n2926) );
  NAND_GATE U4194 ( .I1(n3598), .I2(n2926), .O(n2928) );
  INV_GATE U4195 ( .I1(n3599), .O(n3595) );
  NAND_GATE U4196 ( .I1(n3597), .I2(n3595), .O(n2927) );
  NAND_GATE U4197 ( .I1(n2928), .I2(n2927), .O(n3621) );
  NAND3_GATE U4198 ( .I1(n2929), .I2(n3615), .I3(n3621), .O(n2931) );
  NAND_GATE U4199 ( .I1(B[26]), .I2(A[3]), .O(n3624) );
  INV_GATE U4200 ( .I1(n3624), .O(n3613) );
  NAND3_GATE U4201 ( .I1(n3613), .I2(n3614), .I3(n3615), .O(n2930) );
  NAND_GATE U4202 ( .I1(n3613), .I2(n3621), .O(n3618) );
  NAND3_GATE U4203 ( .I1(n2931), .I2(n2930), .I3(n3618), .O(n3632) );
  NAND_GATE U4204 ( .I1(B[26]), .I2(A[4]), .O(n3871) );
  INV_GATE U4205 ( .I1(n2940), .O(n2938) );
  NAND4_GATE U4206 ( .I1(n2933), .I2(n2934), .I3(n2932), .I4(n2938), .O(n2946)
         );
  NAND_GATE U4207 ( .I1(n2934), .I2(n2933), .O(n2935) );
  NAND_GATE U4208 ( .I1(n2936), .I2(n2935), .O(n2939) );
  OR_GATE U4209 ( .I1(n2939), .I2(n2937), .O(n2945) );
  NAND_GATE U4210 ( .I1(n2938), .I2(n2939), .O(n2942) );
  NAND3_GATE U4211 ( .I1(n2943), .I2(n2942), .I3(n2941), .O(n2944) );
  NAND3_GATE U4212 ( .I1(n2946), .I2(n2945), .I3(n2944), .O(n3637) );
  NAND_GATE U4213 ( .I1(n3871), .I2(n3637), .O(n2947) );
  NAND_GATE U4214 ( .I1(n3632), .I2(n2947), .O(n2949) );
  INV_GATE U4215 ( .I1(n3871), .O(n3869) );
  NAND_GATE U4216 ( .I1(n3869), .I2(n573), .O(n2948) );
  NAND_GATE U4217 ( .I1(n2949), .I2(n2948), .O(n3641) );
  NAND4_GATE U4218 ( .I1(n2954), .I2(n2951), .I3(n2963), .I4(n2950), .O(n2962)
         );
  NAND3_GATE U4219 ( .I1(n2963), .I2(n2951), .I3(n2950), .O(n2956) );
  NAND_GATE U4220 ( .I1(n2954), .I2(n2963), .O(n2955) );
  NAND3_GATE U4221 ( .I1(n751), .I2(n2953), .I3(n2960), .O(n2959) );
  NAND4_GATE U4222 ( .I1(n2956), .I2(n2955), .I3(n2959), .I4(n2958), .O(n2957)
         );
  NAND_GATE U4223 ( .I1(n2962), .I2(n2957), .O(n3649) );
  NAND_GATE U4224 ( .I1(n3641), .I2(n3649), .O(n2965) );
  NAND_GATE U4225 ( .I1(n751), .I2(n2960), .O(n2961) );
  NAND3_GATE U4226 ( .I1(n2963), .I2(n2962), .I3(n2961), .O(n3646) );
  NAND_GATE U4227 ( .I1(B[26]), .I2(A[5]), .O(n3644) );
  INV_GATE U4228 ( .I1(n3644), .O(n3647) );
  NAND3_GATE U4229 ( .I1(n1153), .I2(n3646), .I3(n3647), .O(n2964) );
  NAND_GATE U4230 ( .I1(n3647), .I2(n3641), .O(n3648) );
  NAND3_GATE U4231 ( .I1(n2965), .I2(n2964), .I3(n3648), .O(n3660) );
  NAND3_GATE U4232 ( .I1(n2967), .I2(n2966), .I3(n3660), .O(n2968) );
  NAND_GATE U4233 ( .I1(n2969), .I2(n2968), .O(n3672) );
  NAND_GATE U4234 ( .I1(n1262), .I2(n2970), .O(n2977) );
  INV_GATE U4235 ( .I1(n2970), .O(n2975) );
  NAND_GATE U4236 ( .I1(n2979), .I2(n2970), .O(n2973) );
  NAND3_GATE U4237 ( .I1(n750), .I2(n2971), .I3(n2970), .O(n2980) );
  NAND4_GATE U4238 ( .I1(n2981), .I2(n2973), .I3(n2972), .I4(n2980), .O(n2974)
         );
  NAND_GATE U4239 ( .I1(n2977), .I2(n2974), .O(n3667) );
  NAND_GATE U4240 ( .I1(n3672), .I2(n3667), .O(n2985) );
  NAND_GATE U4241 ( .I1(B[26]), .I2(A[7]), .O(n3678) );
  INV_GATE U4242 ( .I1(n3678), .O(n3670) );
  NAND_GATE U4243 ( .I1(n2976), .I2(n2975), .O(n2978) );
  NAND3_GATE U4244 ( .I1(n2979), .I2(n2978), .I3(n2977), .O(n3669) );
  NAND_GATE U4245 ( .I1(n2981), .I2(n2980), .O(n2982) );
  INV_GATE U4246 ( .I1(n2982), .O(n3668) );
  NAND3_GATE U4247 ( .I1(n3670), .I2(n3669), .I3(n3668), .O(n2984) );
  NAND_GATE U4248 ( .I1(n3670), .I2(n3672), .O(n2983) );
  NAND3_GATE U4249 ( .I1(n2985), .I2(n2984), .I3(n2983), .O(n3692) );
  NAND_GATE U4250 ( .I1(n2986), .I2(n839), .O(n3686) );
  NAND_GATE U4251 ( .I1(n3685), .I2(n3686), .O(n2989) );
  NAND3_GATE U4252 ( .I1(n2986), .I2(n839), .I3(n2987), .O(n3687) );
  NAND3_GATE U4253 ( .I1(n2991), .I2(n2988), .I3(n2987), .O(n3688) );
  NAND3_GATE U4254 ( .I1(n2989), .I2(n3687), .I3(n3688), .O(n2992) );
  NAND_GATE U4255 ( .I1(n2992), .I2(n3684), .O(n3683) );
  NAND_GATE U4256 ( .I1(n3692), .I2(n3683), .O(n2995) );
  NAND_GATE U4257 ( .I1(B[26]), .I2(A[8]), .O(n3700) );
  INV_GATE U4258 ( .I1(n3700), .O(n3693) );
  NAND_GATE U4259 ( .I1(n3693), .I2(n3683), .O(n2994) );
  NAND_GATE U4260 ( .I1(n3693), .I2(n3692), .O(n2993) );
  NAND3_GATE U4261 ( .I1(n2995), .I2(n2994), .I3(n2993), .O(n3587) );
  NAND3_GATE U4262 ( .I1(n871), .I2(n2998), .I3(n2997), .O(n3002) );
  NAND_GATE U4263 ( .I1(n3006), .I2(n3005), .O(n3000) );
  NAND_GATE U4264 ( .I1(n3004), .I2(n3001), .O(n3585) );
  NAND_GATE U4265 ( .I1(n3587), .I2(n3585), .O(n3010) );
  NAND_GATE U4266 ( .I1(B[26]), .I2(A[9]), .O(n3709) );
  INV_GATE U4267 ( .I1(n3709), .O(n3588) );
  NAND_GATE U4268 ( .I1(n3588), .I2(n3587), .O(n3009) );
  AND3_GATE U4269 ( .I1(n3003), .I2(n3002), .I3(n3588), .O(n3008) );
  NAND3_GATE U4270 ( .I1(n3006), .I2(n3005), .I3(n3004), .O(n3007) );
  NAND_GATE U4271 ( .I1(n3008), .I2(n3007), .O(n3586) );
  NAND3_GATE U4272 ( .I1(n3010), .I2(n3009), .I3(n3586), .O(n3578) );
  NAND3_GATE U4273 ( .I1(n3013), .I2(n3012), .I3(n873), .O(n3017) );
  NAND3_GATE U4274 ( .I1(n781), .I2(n3012), .I3(n273), .O(n3016) );
  NAND_GATE U4275 ( .I1(n3013), .I2(n873), .O(n3019) );
  NAND_GATE U4276 ( .I1(n3020), .I2(n3019), .O(n3014) );
  NAND3_GATE U4277 ( .I1(n3017), .I2(n3016), .I3(n3014), .O(n3015) );
  NAND_GATE U4278 ( .I1(n3578), .I2(n3579), .O(n3024) );
  NAND_GATE U4279 ( .I1(B[26]), .I2(A[10]), .O(n3582) );
  INV_GATE U4280 ( .I1(n3582), .O(n3575) );
  NAND_GATE U4281 ( .I1(n3575), .I2(n3578), .O(n3023) );
  AND3_GATE U4282 ( .I1(n3017), .I2(n3016), .I3(n3575), .O(n3022) );
  NAND3_GATE U4283 ( .I1(n3020), .I2(n3019), .I3(n3018), .O(n3021) );
  NAND_GATE U4284 ( .I1(n3022), .I2(n3021), .O(n3574) );
  NAND3_GATE U4285 ( .I1(n3024), .I2(n3023), .I3(n3574), .O(n3567) );
  NAND_GATE U4286 ( .I1(n3034), .I2(n3567), .O(n3569) );
  NAND_GATE U4287 ( .I1(n3030), .I2(n1150), .O(n3025) );
  NAND_GATE U4288 ( .I1(n3026), .I2(n3025), .O(n3036) );
  NAND3_GATE U4289 ( .I1(n3029), .I2(n3031), .I3(n3028), .O(n3033) );
  NAND3_GATE U4290 ( .I1(n1150), .I2(n3031), .I3(n3030), .O(n3032) );
  AND_GATE U4291 ( .I1(n3033), .I2(n3032), .O(n3037) );
  NAND3_GATE U4292 ( .I1(n3035), .I2(n3037), .I3(n3034), .O(n3568) );
  NAND_GATE U4293 ( .I1(n3037), .I2(n3036), .O(n3038) );
  NAND_GATE U4294 ( .I1(n3039), .I2(n3038), .O(n3570) );
  NAND_GATE U4295 ( .I1(n3567), .I2(n3570), .O(n3040) );
  NAND3_GATE U4296 ( .I1(n3569), .I2(n3568), .I3(n3040), .O(n3558) );
  NAND_GATE U4297 ( .I1(n3557), .I2(n3558), .O(n3059) );
  NAND_GATE U4298 ( .I1(B[26]), .I2(A[13]), .O(n3546) );
  INV_GATE U4299 ( .I1(n3546), .O(n3548) );
  NAND_GATE U4300 ( .I1(B[26]), .I2(A[12]), .O(n3559) );
  INV_GATE U4301 ( .I1(n3559), .O(n3041) );
  NAND_GATE U4302 ( .I1(n3558), .I2(n3041), .O(n3553) );
  NAND_GATE U4303 ( .I1(n3557), .I2(n3041), .O(n3552) );
  NAND_GATE U4304 ( .I1(n3553), .I2(n3552), .O(n3058) );
  NAND_GATE U4305 ( .I1(n1309), .I2(n3049), .O(n3043) );
  INV_GATE U4306 ( .I1(n3049), .O(n3044) );
  NAND_GATE U4307 ( .I1(n3043), .I2(n3042), .O(n3052) );
  NAND_GATE U4308 ( .I1(n3045), .I2(n3044), .O(n3046) );
  NAND_GATE U4309 ( .I1(n3047), .I2(n3046), .O(n3055) );
  INV_GATE U4310 ( .I1(n3055), .O(n3050) );
  NAND_GATE U4311 ( .I1(n3050), .I2(n3057), .O(n3051) );
  NAND_GATE U4312 ( .I1(n3053), .I2(n3052), .O(n3054) );
  NAND_GATE U4313 ( .I1(n3055), .I2(n3054), .O(n3056) );
  NAND_GATE U4314 ( .I1(n3057), .I2(n3056), .O(n3543) );
  NAND_GATE U4315 ( .I1(n3074), .I2(n3537), .O(n3533) );
  INV_GATE U4316 ( .I1(n3060), .O(n3061) );
  NAND_GATE U4317 ( .I1(n3061), .I2(n3064), .O(n3073) );
  NAND_GATE U4318 ( .I1(n3066), .I2(n222), .O(n3062) );
  NAND_GATE U4319 ( .I1(n3063), .I2(n3062), .O(n3071) );
  NAND_GATE U4320 ( .I1(n3065), .I2(n3064), .O(n3067) );
  NAND_GATE U4321 ( .I1(n3067), .I2(n3062), .O(n3068) );
  NAND_GATE U4322 ( .I1(n3069), .I2(n3068), .O(n3070) );
  NAND_GATE U4323 ( .I1(n3071), .I2(n3070), .O(n3072) );
  NAND_GATE U4324 ( .I1(n3073), .I2(n3072), .O(n3536) );
  NAND_GATE U4325 ( .I1(n3074), .I2(n3536), .O(n3532) );
  NAND_GATE U4326 ( .I1(n3537), .I2(n3536), .O(n3075) );
  NAND3_GATE U4327 ( .I1(n3533), .I2(n3532), .I3(n3075), .O(n3526) );
  NAND_GATE U4328 ( .I1(n3091), .I2(n3526), .O(n3522) );
  INV_GATE U4329 ( .I1(n3076), .O(n3077) );
  NAND_GATE U4330 ( .I1(n3077), .I2(n3080), .O(n3090) );
  INV_GATE U4331 ( .I1(n3080), .O(n3082) );
  NAND_GATE U4332 ( .I1(n3083), .I2(n3082), .O(n3078) );
  NAND_GATE U4333 ( .I1(n3079), .I2(n3078), .O(n3088) );
  NAND_GATE U4334 ( .I1(n3081), .I2(n3080), .O(n3084) );
  NAND_GATE U4335 ( .I1(n3084), .I2(n3078), .O(n3085) );
  NAND_GATE U4336 ( .I1(n3086), .I2(n3085), .O(n3087) );
  NAND_GATE U4337 ( .I1(n3088), .I2(n3087), .O(n3089) );
  NAND_GATE U4338 ( .I1(n3090), .I2(n3089), .O(n3525) );
  NAND_GATE U4339 ( .I1(n3091), .I2(n3525), .O(n3521) );
  NAND_GATE U4340 ( .I1(n3526), .I2(n3525), .O(n3092) );
  NAND3_GATE U4341 ( .I1(n3522), .I2(n3521), .I3(n3092), .O(n3515) );
  NAND_GATE U4342 ( .I1(n3107), .I2(n3515), .O(n3511) );
  INV_GATE U4343 ( .I1(n3093), .O(n3094) );
  NAND_GATE U4344 ( .I1(n3094), .I2(n3097), .O(n3106) );
  NAND_GATE U4345 ( .I1(n3096), .I2(n3100), .O(n3104) );
  NAND_GATE U4346 ( .I1(n3098), .I2(n3097), .O(n3099) );
  NAND_GATE U4347 ( .I1(n3100), .I2(n3099), .O(n3101) );
  NAND_GATE U4348 ( .I1(n3102), .I2(n3101), .O(n3103) );
  NAND_GATE U4349 ( .I1(n3104), .I2(n3103), .O(n3105) );
  NAND_GATE U4350 ( .I1(n3106), .I2(n3105), .O(n3514) );
  NAND_GATE U4351 ( .I1(n3107), .I2(n3514), .O(n3510) );
  NAND_GATE U4352 ( .I1(n3515), .I2(n3514), .O(n3108) );
  NAND3_GATE U4353 ( .I1(n3511), .I2(n3510), .I3(n3108), .O(n3504) );
  NAND_GATE U4354 ( .I1(n3123), .I2(n3504), .O(n3500) );
  INV_GATE U4355 ( .I1(n3109), .O(n3110) );
  NAND_GATE U4356 ( .I1(n3110), .I2(n3113), .O(n3122) );
  NAND_GATE U4357 ( .I1(n3112), .I2(n3116), .O(n3120) );
  NAND_GATE U4358 ( .I1(n3114), .I2(n3113), .O(n3115) );
  NAND_GATE U4359 ( .I1(n3116), .I2(n3115), .O(n3117) );
  NAND_GATE U4360 ( .I1(n3118), .I2(n3117), .O(n3119) );
  NAND_GATE U4361 ( .I1(n3120), .I2(n3119), .O(n3121) );
  NAND_GATE U4362 ( .I1(n3122), .I2(n3121), .O(n3503) );
  NAND_GATE U4363 ( .I1(n3123), .I2(n3503), .O(n3499) );
  NAND_GATE U4364 ( .I1(n3504), .I2(n3503), .O(n3124) );
  NAND3_GATE U4365 ( .I1(n3500), .I2(n3499), .I3(n3124), .O(n3493) );
  NAND_GATE U4366 ( .I1(n3139), .I2(n3493), .O(n3489) );
  INV_GATE U4367 ( .I1(n3125), .O(n3126) );
  NAND_GATE U4368 ( .I1(n3126), .I2(n3129), .O(n3138) );
  NAND_GATE U4369 ( .I1(n3128), .I2(n3132), .O(n3136) );
  NAND_GATE U4370 ( .I1(n3130), .I2(n3129), .O(n3131) );
  NAND_GATE U4371 ( .I1(n3132), .I2(n3131), .O(n3133) );
  NAND_GATE U4372 ( .I1(n3134), .I2(n3133), .O(n3135) );
  NAND_GATE U4373 ( .I1(n3136), .I2(n3135), .O(n3137) );
  NAND_GATE U4374 ( .I1(n3138), .I2(n3137), .O(n3492) );
  NAND_GATE U4375 ( .I1(n3139), .I2(n3492), .O(n3488) );
  NAND_GATE U4376 ( .I1(n3493), .I2(n3492), .O(n3140) );
  NAND3_GATE U4377 ( .I1(n3489), .I2(n3488), .I3(n3140), .O(n3482) );
  NAND_GATE U4378 ( .I1(n3155), .I2(n3482), .O(n3478) );
  INV_GATE U4379 ( .I1(n3141), .O(n3142) );
  NAND_GATE U4380 ( .I1(n3142), .I2(n3145), .O(n3154) );
  NAND_GATE U4381 ( .I1(n3144), .I2(n3148), .O(n3152) );
  NAND_GATE U4382 ( .I1(n3146), .I2(n3145), .O(n3147) );
  NAND_GATE U4383 ( .I1(n3148), .I2(n3147), .O(n3149) );
  NAND_GATE U4384 ( .I1(n3150), .I2(n3149), .O(n3151) );
  NAND_GATE U4385 ( .I1(n3152), .I2(n3151), .O(n3153) );
  NAND_GATE U4386 ( .I1(n3154), .I2(n3153), .O(n3481) );
  NAND_GATE U4387 ( .I1(n3155), .I2(n3481), .O(n3477) );
  NAND_GATE U4388 ( .I1(n3482), .I2(n3481), .O(n3156) );
  NAND3_GATE U4389 ( .I1(n3478), .I2(n3477), .I3(n3156), .O(n3471) );
  NAND_GATE U4390 ( .I1(n3171), .I2(n3471), .O(n3467) );
  INV_GATE U4391 ( .I1(n3157), .O(n3158) );
  NAND_GATE U4392 ( .I1(n3158), .I2(n3161), .O(n3170) );
  NAND_GATE U4393 ( .I1(n3160), .I2(n3164), .O(n3168) );
  NAND_GATE U4394 ( .I1(n3162), .I2(n3161), .O(n3163) );
  NAND_GATE U4395 ( .I1(n3164), .I2(n3163), .O(n3165) );
  NAND_GATE U4396 ( .I1(n3166), .I2(n3165), .O(n3167) );
  NAND_GATE U4397 ( .I1(n3168), .I2(n3167), .O(n3169) );
  NAND_GATE U4398 ( .I1(n3170), .I2(n3169), .O(n3470) );
  NAND_GATE U4399 ( .I1(n3171), .I2(n3470), .O(n3466) );
  NAND_GATE U4400 ( .I1(n3471), .I2(n3470), .O(n3172) );
  NAND3_GATE U4401 ( .I1(n3467), .I2(n3466), .I3(n3172), .O(n3460) );
  NAND_GATE U4402 ( .I1(n3188), .I2(n3460), .O(n3456) );
  INV_GATE U4403 ( .I1(n3173), .O(n3174) );
  NAND_GATE U4404 ( .I1(n3174), .I2(n3178), .O(n3187) );
  INV_GATE U4405 ( .I1(n3178), .O(n3175) );
  NAND_GATE U4406 ( .I1(n3176), .I2(n3175), .O(n3181) );
  NAND_GATE U4407 ( .I1(n3177), .I2(n3181), .O(n3185) );
  NAND_GATE U4408 ( .I1(n3179), .I2(n3178), .O(n3180) );
  NAND_GATE U4409 ( .I1(n3181), .I2(n3180), .O(n3182) );
  NAND_GATE U4410 ( .I1(n3183), .I2(n3182), .O(n3184) );
  NAND_GATE U4411 ( .I1(n3185), .I2(n3184), .O(n3186) );
  NAND_GATE U4412 ( .I1(n3187), .I2(n3186), .O(n3459) );
  NAND_GATE U4413 ( .I1(n3188), .I2(n3459), .O(n3455) );
  NAND_GATE U4414 ( .I1(n3460), .I2(n3459), .O(n3189) );
  NAND3_GATE U4415 ( .I1(n3456), .I2(n3455), .I3(n3189), .O(n3449) );
  NAND_GATE U4416 ( .I1(n3205), .I2(n3449), .O(n3445) );
  INV_GATE U4417 ( .I1(n3190), .O(n3191) );
  NAND_GATE U4418 ( .I1(n3191), .I2(n3195), .O(n3204) );
  INV_GATE U4419 ( .I1(n3195), .O(n3192) );
  NAND_GATE U4420 ( .I1(n3193), .I2(n3192), .O(n3198) );
  NAND_GATE U4421 ( .I1(n3194), .I2(n3198), .O(n3202) );
  NAND_GATE U4422 ( .I1(n3196), .I2(n3195), .O(n3197) );
  NAND_GATE U4423 ( .I1(n3198), .I2(n3197), .O(n3199) );
  NAND_GATE U4424 ( .I1(n3200), .I2(n3199), .O(n3201) );
  NAND_GATE U4425 ( .I1(n3202), .I2(n3201), .O(n3203) );
  NAND_GATE U4426 ( .I1(n3204), .I2(n3203), .O(n3448) );
  NAND_GATE U4427 ( .I1(n3205), .I2(n3448), .O(n3444) );
  NAND_GATE U4428 ( .I1(n3449), .I2(n3448), .O(n3206) );
  NAND3_GATE U4429 ( .I1(n3445), .I2(n3444), .I3(n3206), .O(n3438) );
  NAND_GATE U4430 ( .I1(n3222), .I2(n3438), .O(n3434) );
  INV_GATE U4431 ( .I1(n3207), .O(n3208) );
  NAND_GATE U4432 ( .I1(n3208), .I2(n3212), .O(n3221) );
  INV_GATE U4433 ( .I1(n3212), .O(n3209) );
  NAND_GATE U4434 ( .I1(n3210), .I2(n3209), .O(n3215) );
  NAND_GATE U4435 ( .I1(n3211), .I2(n3215), .O(n3219) );
  NAND_GATE U4436 ( .I1(n3213), .I2(n3212), .O(n3214) );
  NAND_GATE U4437 ( .I1(n3215), .I2(n3214), .O(n3216) );
  NAND_GATE U4438 ( .I1(n3217), .I2(n3216), .O(n3218) );
  NAND_GATE U4439 ( .I1(n3219), .I2(n3218), .O(n3220) );
  NAND_GATE U4440 ( .I1(n3221), .I2(n3220), .O(n3437) );
  NAND_GATE U4441 ( .I1(n3222), .I2(n3437), .O(n3433) );
  NAND_GATE U4442 ( .I1(n3438), .I2(n3437), .O(n3223) );
  NAND3_GATE U4443 ( .I1(n3434), .I2(n3433), .I3(n3223), .O(n3427) );
  NAND_GATE U4444 ( .I1(n3238), .I2(n3427), .O(n3423) );
  INV_GATE U4445 ( .I1(n3224), .O(n3225) );
  NAND_GATE U4446 ( .I1(n3225), .I2(n3228), .O(n3237) );
  NAND_GATE U4447 ( .I1(n3227), .I2(n3231), .O(n3235) );
  NAND_GATE U4448 ( .I1(n3229), .I2(n3228), .O(n3230) );
  NAND_GATE U4449 ( .I1(n3231), .I2(n3230), .O(n3232) );
  NAND_GATE U4450 ( .I1(n3233), .I2(n3232), .O(n3234) );
  NAND_GATE U4451 ( .I1(n3235), .I2(n3234), .O(n3236) );
  NAND_GATE U4452 ( .I1(n3237), .I2(n3236), .O(n3426) );
  NAND_GATE U4453 ( .I1(n3238), .I2(n3426), .O(n3422) );
  NAND_GATE U4454 ( .I1(n3427), .I2(n3426), .O(n3239) );
  NAND3_GATE U4455 ( .I1(n3423), .I2(n3422), .I3(n3239), .O(n3752) );
  NAND_GATE U4456 ( .I1(n3254), .I2(n3752), .O(n3748) );
  INV_GATE U4457 ( .I1(n3240), .O(n3241) );
  NAND_GATE U4458 ( .I1(n3241), .I2(n3244), .O(n3253) );
  NAND_GATE U4459 ( .I1(n3243), .I2(n3247), .O(n3251) );
  NAND_GATE U4460 ( .I1(n3245), .I2(n3244), .O(n3246) );
  NAND_GATE U4461 ( .I1(n3247), .I2(n3246), .O(n3248) );
  NAND_GATE U4462 ( .I1(n3249), .I2(n3248), .O(n3250) );
  NAND_GATE U4463 ( .I1(n3251), .I2(n3250), .O(n3252) );
  NAND_GATE U4464 ( .I1(n3253), .I2(n3252), .O(n3751) );
  NAND_GATE U4465 ( .I1(n3254), .I2(n3751), .O(n3747) );
  NAND_GATE U4466 ( .I1(n3752), .I2(n3751), .O(n3255) );
  NAND3_GATE U4467 ( .I1(n3748), .I2(n3747), .I3(n3255), .O(n3416) );
  NAND_GATE U4468 ( .I1(n3270), .I2(n3416), .O(n3412) );
  INV_GATE U4469 ( .I1(n3256), .O(n3257) );
  NAND_GATE U4470 ( .I1(n3257), .I2(n3260), .O(n3269) );
  NAND_GATE U4471 ( .I1(n3259), .I2(n3263), .O(n3267) );
  NAND_GATE U4472 ( .I1(n3261), .I2(n3260), .O(n3262) );
  NAND_GATE U4473 ( .I1(n3263), .I2(n3262), .O(n3264) );
  NAND_GATE U4474 ( .I1(n3265), .I2(n3264), .O(n3266) );
  NAND_GATE U4475 ( .I1(n3267), .I2(n3266), .O(n3268) );
  NAND_GATE U4476 ( .I1(n3269), .I2(n3268), .O(n3415) );
  NAND_GATE U4477 ( .I1(n3270), .I2(n3415), .O(n3411) );
  NAND_GATE U4478 ( .I1(n3416), .I2(n3415), .O(n3271) );
  NAND3_GATE U4479 ( .I1(n3412), .I2(n3411), .I3(n3271), .O(n3405) );
  NAND_GATE U4480 ( .I1(n3272), .I2(n3405), .O(n3400) );
  NAND_GATE U4481 ( .I1(n3404), .I2(n3405), .O(n3273) );
  NAND3_GATE U4482 ( .I1(n3401), .I2(n3400), .I3(n3273), .O(n3394) );
  NAND_GATE U4483 ( .I1(n3288), .I2(n3394), .O(n3390) );
  INV_GATE U4484 ( .I1(n3274), .O(n3275) );
  NAND_GATE U4485 ( .I1(n3275), .I2(n3278), .O(n3287) );
  NAND_GATE U4486 ( .I1(n3277), .I2(n3281), .O(n3285) );
  NAND_GATE U4487 ( .I1(n3279), .I2(n3278), .O(n3280) );
  NAND_GATE U4488 ( .I1(n3281), .I2(n3280), .O(n3282) );
  NAND_GATE U4489 ( .I1(n3283), .I2(n3282), .O(n3284) );
  NAND_GATE U4490 ( .I1(n3285), .I2(n3284), .O(n3286) );
  NAND_GATE U4491 ( .I1(n3287), .I2(n3286), .O(n3393) );
  NAND_GATE U4492 ( .I1(n3288), .I2(n3393), .O(n3389) );
  NAND_GATE U4493 ( .I1(n3394), .I2(n3393), .O(n3289) );
  NAND3_GATE U4494 ( .I1(n3390), .I2(n3389), .I3(n3289), .O(n3383) );
  NAND_GATE U4495 ( .I1(n3304), .I2(n3383), .O(n3379) );
  OR_GATE U4496 ( .I1(n3291), .I2(n3290), .O(n3303) );
  NAND_GATE U4497 ( .I1(n3292), .I2(n3291), .O(n3297) );
  NAND_GATE U4498 ( .I1(n3293), .I2(n3297), .O(n3301) );
  NAND_GATE U4499 ( .I1(n3295), .I2(n3294), .O(n3296) );
  NAND_GATE U4500 ( .I1(n3297), .I2(n3296), .O(n3298) );
  NAND_GATE U4501 ( .I1(n3299), .I2(n3298), .O(n3300) );
  NAND_GATE U4502 ( .I1(n3301), .I2(n3300), .O(n3302) );
  NAND_GATE U4503 ( .I1(n3303), .I2(n3302), .O(n3382) );
  NAND_GATE U4504 ( .I1(n3304), .I2(n3382), .O(n3378) );
  NAND_GATE U4505 ( .I1(n3383), .I2(n3382), .O(n3305) );
  NAND3_GATE U4506 ( .I1(n3379), .I2(n3378), .I3(n3305), .O(n3372) );
  NAND_GATE U4507 ( .I1(n3320), .I2(n3372), .O(n3368) );
  INV_GATE U4508 ( .I1(n3306), .O(n3307) );
  NAND_GATE U4509 ( .I1(n3307), .I2(n3310), .O(n3319) );
  NAND_GATE U4510 ( .I1(n3309), .I2(n3313), .O(n3317) );
  NAND_GATE U4511 ( .I1(n3311), .I2(n3310), .O(n3312) );
  NAND_GATE U4512 ( .I1(n3313), .I2(n3312), .O(n3314) );
  NAND_GATE U4513 ( .I1(n3315), .I2(n3314), .O(n3316) );
  NAND_GATE U4514 ( .I1(n3317), .I2(n3316), .O(n3318) );
  NAND_GATE U4515 ( .I1(n3319), .I2(n3318), .O(n3371) );
  NAND_GATE U4516 ( .I1(n3320), .I2(n3371), .O(n3367) );
  NAND_GATE U4517 ( .I1(n3372), .I2(n3371), .O(n3321) );
  NAND3_GATE U4518 ( .I1(n3368), .I2(n3367), .I3(n3321), .O(n3361) );
  NAND_GATE U4519 ( .I1(n3336), .I2(n3361), .O(n3357) );
  INV_GATE U4520 ( .I1(n3322), .O(n3323) );
  NAND_GATE U4521 ( .I1(n3323), .I2(n3326), .O(n3335) );
  NAND_GATE U4522 ( .I1(n3325), .I2(n3329), .O(n3333) );
  NAND_GATE U4523 ( .I1(n3327), .I2(n3326), .O(n3328) );
  NAND_GATE U4524 ( .I1(n3329), .I2(n3328), .O(n3330) );
  NAND_GATE U4525 ( .I1(n3331), .I2(n3330), .O(n3332) );
  NAND_GATE U4526 ( .I1(n3333), .I2(n3332), .O(n3334) );
  NAND_GATE U4527 ( .I1(n3335), .I2(n3334), .O(n3360) );
  NAND_GATE U4528 ( .I1(n3336), .I2(n3360), .O(n3356) );
  NAND_GATE U4529 ( .I1(n3361), .I2(n3360), .O(n3337) );
  NAND3_GATE U4530 ( .I1(n3357), .I2(n3356), .I3(n3337), .O(n15312) );
  INV_GATE U4531 ( .I1(n15312), .O(n3352) );
  INV_GATE U4532 ( .I1(n3338), .O(n3339) );
  NAND_GATE U4533 ( .I1(n3339), .I2(n3342), .O(n3351) );
  NAND_GATE U4534 ( .I1(n3341), .I2(n3345), .O(n3349) );
  NAND_GATE U4535 ( .I1(n3343), .I2(n3342), .O(n3344) );
  NAND_GATE U4536 ( .I1(n3345), .I2(n3344), .O(n3346) );
  NAND_GATE U4537 ( .I1(n3347), .I2(n3346), .O(n3348) );
  NAND_GATE U4538 ( .I1(n3349), .I2(n3348), .O(n3350) );
  NAND_GATE U4539 ( .I1(n3351), .I2(n3350), .O(n15311) );
  NAND_GATE U4540 ( .I1(n3352), .I2(n15311), .O(n3355) );
  INV_GATE U4541 ( .I1(n15311), .O(n3353) );
  NAND_GATE U4542 ( .I1(n15312), .I2(n3353), .O(n3354) );
  NAND_GATE U4543 ( .I1(n3355), .I2(n3354), .O(\A1[56] ) );
  OR_GATE U4544 ( .I1(n3356), .I2(n3361), .O(n3359) );
  OR_GATE U4545 ( .I1(n3360), .I2(n3357), .O(n3358) );
  AND_GATE U4546 ( .I1(n3359), .I2(n3358), .O(n3366) );
  NAND_GATE U4547 ( .I1(n3361), .I2(n1135), .O(n3363) );
  NAND3_GATE U4548 ( .I1(n3364), .I2(n3363), .I3(n3362), .O(n3365) );
  OR_GATE U4549 ( .I1(n3367), .I2(n3372), .O(n3370) );
  OR_GATE U4550 ( .I1(n3371), .I2(n3368), .O(n3369) );
  AND_GATE U4551 ( .I1(n3370), .I2(n3369), .O(n3377) );
  NAND_GATE U4552 ( .I1(n1133), .I2(n3371), .O(n3375) );
  NAND3_GATE U4553 ( .I1(n3375), .I2(n3374), .I3(n3373), .O(n3376) );
  NAND_GATE U4554 ( .I1(n3377), .I2(n3376), .O(n4221) );
  INV_GATE U4555 ( .I1(n4221), .O(n4224) );
  NAND_GATE U4556 ( .I1(B[25]), .I2(A[31]), .O(n4228) );
  INV_GATE U4557 ( .I1(n4228), .O(n4222) );
  NAND_GATE U4558 ( .I1(n4224), .I2(n4222), .O(n4219) );
  OR_GATE U4559 ( .I1(n3378), .I2(n3383), .O(n3381) );
  OR_GATE U4560 ( .I1(n3382), .I2(n3379), .O(n3380) );
  AND_GATE U4561 ( .I1(n3381), .I2(n3380), .O(n3388) );
  NAND_GATE U4562 ( .I1(n3383), .I2(n1131), .O(n3385) );
  NAND3_GATE U4563 ( .I1(n3386), .I2(n3385), .I3(n3384), .O(n3387) );
  NAND_GATE U4564 ( .I1(n3388), .I2(n3387), .O(n4205) );
  INV_GATE U4565 ( .I1(n4205), .O(n4208) );
  NAND_GATE U4566 ( .I1(B[25]), .I2(A[30]), .O(n4212) );
  INV_GATE U4567 ( .I1(n4212), .O(n4206) );
  NAND_GATE U4568 ( .I1(n4208), .I2(n4206), .O(n4203) );
  OR_GATE U4569 ( .I1(n3389), .I2(n3394), .O(n3392) );
  OR_GATE U4570 ( .I1(n3393), .I2(n3390), .O(n3391) );
  AND_GATE U4571 ( .I1(n3392), .I2(n3391), .O(n3399) );
  NAND_GATE U4572 ( .I1(n3394), .I2(n1128), .O(n3396) );
  NAND3_GATE U4573 ( .I1(n3397), .I2(n3396), .I3(n3395), .O(n3398) );
  NAND_GATE U4574 ( .I1(n3399), .I2(n3398), .O(n4189) );
  INV_GATE U4575 ( .I1(n4189), .O(n4192) );
  NAND_GATE U4576 ( .I1(B[25]), .I2(A[29]), .O(n4196) );
  INV_GATE U4577 ( .I1(n4196), .O(n4190) );
  NAND_GATE U4578 ( .I1(n4192), .I2(n4190), .O(n4187) );
  OR_GATE U4579 ( .I1(n3400), .I2(n3404), .O(n3403) );
  OR_GATE U4580 ( .I1(n3405), .I2(n3401), .O(n3402) );
  AND_GATE U4581 ( .I1(n3403), .I2(n3402), .O(n3410) );
  NAND_GATE U4582 ( .I1(n1125), .I2(n3405), .O(n3407) );
  NAND3_GATE U4583 ( .I1(n3408), .I2(n3407), .I3(n3406), .O(n3409) );
  NAND_GATE U4584 ( .I1(n3410), .I2(n3409), .O(n4173) );
  INV_GATE U4585 ( .I1(n4173), .O(n4176) );
  NAND_GATE U4586 ( .I1(B[25]), .I2(A[28]), .O(n4180) );
  INV_GATE U4587 ( .I1(n4180), .O(n4174) );
  NAND_GATE U4588 ( .I1(n4176), .I2(n4174), .O(n4171) );
  OR_GATE U4589 ( .I1(n3411), .I2(n3416), .O(n3414) );
  OR_GATE U4590 ( .I1(n3415), .I2(n3412), .O(n3413) );
  AND_GATE U4591 ( .I1(n3414), .I2(n3413), .O(n3421) );
  NAND_GATE U4592 ( .I1(n3416), .I2(n1117), .O(n3418) );
  NAND3_GATE U4593 ( .I1(n3419), .I2(n3418), .I3(n3417), .O(n3420) );
  NAND_GATE U4594 ( .I1(n3421), .I2(n3420), .O(n4157) );
  INV_GATE U4595 ( .I1(n4157), .O(n4160) );
  NAND_GATE U4596 ( .I1(B[25]), .I2(A[27]), .O(n4164) );
  INV_GATE U4597 ( .I1(n4164), .O(n4158) );
  NAND_GATE U4598 ( .I1(n4160), .I2(n4158), .O(n4155) );
  NAND_GATE U4599 ( .I1(B[25]), .I2(A[26]), .O(n4148) );
  INV_GATE U4600 ( .I1(n4148), .O(n4142) );
  OR_GATE U4601 ( .I1(n3422), .I2(n3427), .O(n3425) );
  OR_GATE U4602 ( .I1(n3426), .I2(n3423), .O(n3424) );
  AND_GATE U4603 ( .I1(n3425), .I2(n3424), .O(n3432) );
  NAND_GATE U4604 ( .I1(n1099), .I2(n3426), .O(n3430) );
  NAND3_GATE U4605 ( .I1(n3430), .I2(n3429), .I3(n3428), .O(n3431) );
  NAND_GATE U4606 ( .I1(n3432), .I2(n3431), .O(n4125) );
  INV_GATE U4607 ( .I1(n4125), .O(n4128) );
  NAND_GATE U4608 ( .I1(B[25]), .I2(A[25]), .O(n4132) );
  INV_GATE U4609 ( .I1(n4132), .O(n4126) );
  NAND_GATE U4610 ( .I1(n4128), .I2(n4126), .O(n4122) );
  OR_GATE U4611 ( .I1(n3433), .I2(n3438), .O(n3436) );
  OR_GATE U4612 ( .I1(n3437), .I2(n3434), .O(n3435) );
  AND_GATE U4613 ( .I1(n3436), .I2(n3435), .O(n3443) );
  NAND_GATE U4614 ( .I1(n1093), .I2(n3437), .O(n3441) );
  NAND3_GATE U4615 ( .I1(n3441), .I2(n3440), .I3(n3439), .O(n3442) );
  NAND_GATE U4616 ( .I1(n3443), .I2(n3442), .O(n3775) );
  INV_GATE U4617 ( .I1(n3775), .O(n3778) );
  NAND_GATE U4618 ( .I1(B[25]), .I2(A[24]), .O(n3782) );
  INV_GATE U4619 ( .I1(n3782), .O(n3776) );
  NAND_GATE U4620 ( .I1(n3778), .I2(n3776), .O(n3772) );
  OR_GATE U4621 ( .I1(n3444), .I2(n3449), .O(n3447) );
  OR_GATE U4622 ( .I1(n3448), .I2(n3445), .O(n3446) );
  AND_GATE U4623 ( .I1(n3447), .I2(n3446), .O(n3454) );
  NAND_GATE U4624 ( .I1(n1087), .I2(n3448), .O(n3452) );
  NAND3_GATE U4625 ( .I1(n3452), .I2(n3451), .I3(n3450), .O(n3453) );
  NAND_GATE U4626 ( .I1(n3454), .I2(n3453), .O(n4106) );
  INV_GATE U4627 ( .I1(n4106), .O(n4109) );
  NAND_GATE U4628 ( .I1(B[25]), .I2(A[23]), .O(n4113) );
  INV_GATE U4629 ( .I1(n4113), .O(n4107) );
  NAND_GATE U4630 ( .I1(n4109), .I2(n4107), .O(n4103) );
  OR_GATE U4631 ( .I1(n3455), .I2(n3460), .O(n3458) );
  OR_GATE U4632 ( .I1(n3459), .I2(n3456), .O(n3457) );
  AND_GATE U4633 ( .I1(n3458), .I2(n3457), .O(n3465) );
  NAND_GATE U4634 ( .I1(n1094), .I2(n3459), .O(n3463) );
  NAND3_GATE U4635 ( .I1(n3463), .I2(n3462), .I3(n3461), .O(n3464) );
  NAND_GATE U4636 ( .I1(n3465), .I2(n3464), .O(n4089) );
  INV_GATE U4637 ( .I1(n4089), .O(n4092) );
  NAND_GATE U4638 ( .I1(B[25]), .I2(A[22]), .O(n4096) );
  INV_GATE U4639 ( .I1(n4096), .O(n4090) );
  NAND_GATE U4640 ( .I1(n4092), .I2(n4090), .O(n4087) );
  OR_GATE U4641 ( .I1(n3466), .I2(n3471), .O(n3469) );
  OR_GATE U4642 ( .I1(n3470), .I2(n3467), .O(n3468) );
  AND_GATE U4643 ( .I1(n3469), .I2(n3468), .O(n3476) );
  NAND_GATE U4644 ( .I1(n3471), .I2(n1079), .O(n3473) );
  NAND3_GATE U4645 ( .I1(n3474), .I2(n3473), .I3(n3472), .O(n3475) );
  NAND_GATE U4646 ( .I1(n3476), .I2(n3475), .O(n4073) );
  INV_GATE U4647 ( .I1(n4073), .O(n4076) );
  NAND_GATE U4648 ( .I1(B[25]), .I2(A[21]), .O(n4080) );
  INV_GATE U4649 ( .I1(n4080), .O(n4074) );
  NAND_GATE U4650 ( .I1(n4076), .I2(n4074), .O(n4071) );
  OR_GATE U4651 ( .I1(n3477), .I2(n3482), .O(n3480) );
  OR_GATE U4652 ( .I1(n3481), .I2(n3478), .O(n3479) );
  AND_GATE U4653 ( .I1(n3480), .I2(n3479), .O(n3487) );
  NAND_GATE U4654 ( .I1(n3482), .I2(n1063), .O(n3484) );
  NAND3_GATE U4655 ( .I1(n3485), .I2(n3484), .I3(n3483), .O(n3486) );
  NAND_GATE U4656 ( .I1(n3487), .I2(n3486), .O(n4057) );
  INV_GATE U4657 ( .I1(n4057), .O(n4060) );
  NAND_GATE U4658 ( .I1(B[25]), .I2(A[20]), .O(n4064) );
  INV_GATE U4659 ( .I1(n4064), .O(n4058) );
  NAND_GATE U4660 ( .I1(n4060), .I2(n4058), .O(n4055) );
  OR_GATE U4661 ( .I1(n3488), .I2(n3493), .O(n3491) );
  OR_GATE U4662 ( .I1(n3492), .I2(n3489), .O(n3490) );
  AND_GATE U4663 ( .I1(n3491), .I2(n3490), .O(n3498) );
  NAND_GATE U4664 ( .I1(n3493), .I2(n1064), .O(n3495) );
  NAND3_GATE U4665 ( .I1(n3496), .I2(n3495), .I3(n3494), .O(n3497) );
  NAND_GATE U4666 ( .I1(n3498), .I2(n3497), .O(n4041) );
  INV_GATE U4667 ( .I1(n4041), .O(n4044) );
  NAND_GATE U4668 ( .I1(B[25]), .I2(A[19]), .O(n4048) );
  INV_GATE U4669 ( .I1(n4048), .O(n4042) );
  NAND_GATE U4670 ( .I1(n4044), .I2(n4042), .O(n4039) );
  OR_GATE U4671 ( .I1(n3499), .I2(n3504), .O(n3502) );
  OR_GATE U4672 ( .I1(n3503), .I2(n3500), .O(n3501) );
  AND_GATE U4673 ( .I1(n3502), .I2(n3501), .O(n3509) );
  NAND_GATE U4674 ( .I1(n3504), .I2(n1065), .O(n3506) );
  NAND3_GATE U4675 ( .I1(n3507), .I2(n3506), .I3(n3505), .O(n3508) );
  NAND_GATE U4676 ( .I1(n3509), .I2(n3508), .O(n4025) );
  INV_GATE U4677 ( .I1(n4025), .O(n4028) );
  NAND_GATE U4678 ( .I1(B[25]), .I2(A[18]), .O(n4032) );
  INV_GATE U4679 ( .I1(n4032), .O(n4026) );
  NAND_GATE U4680 ( .I1(n4028), .I2(n4026), .O(n4023) );
  OR_GATE U4681 ( .I1(n3510), .I2(n3515), .O(n3513) );
  OR_GATE U4682 ( .I1(n3514), .I2(n3511), .O(n3512) );
  AND_GATE U4683 ( .I1(n3513), .I2(n3512), .O(n3520) );
  NAND_GATE U4684 ( .I1(n3515), .I2(n1068), .O(n3517) );
  NAND3_GATE U4685 ( .I1(n3518), .I2(n3517), .I3(n3516), .O(n3519) );
  NAND_GATE U4686 ( .I1(n3520), .I2(n3519), .O(n4009) );
  INV_GATE U4687 ( .I1(n4009), .O(n4012) );
  NAND_GATE U4688 ( .I1(B[25]), .I2(A[17]), .O(n4016) );
  INV_GATE U4689 ( .I1(n4016), .O(n4010) );
  NAND_GATE U4690 ( .I1(n4012), .I2(n4010), .O(n4007) );
  OR_GATE U4691 ( .I1(n3521), .I2(n3526), .O(n3524) );
  OR_GATE U4692 ( .I1(n3525), .I2(n3522), .O(n3523) );
  AND_GATE U4693 ( .I1(n3524), .I2(n3523), .O(n3531) );
  NAND_GATE U4694 ( .I1(n3526), .I2(n1062), .O(n3528) );
  NAND3_GATE U4695 ( .I1(n3529), .I2(n3528), .I3(n3527), .O(n3530) );
  NAND_GATE U4696 ( .I1(n3531), .I2(n3530), .O(n3997) );
  NAND_GATE U4697 ( .I1(B[25]), .I2(A[16]), .O(n4000) );
  INV_GATE U4698 ( .I1(n4000), .O(n3995) );
  NAND_GATE U4699 ( .I1(n399), .I2(n3995), .O(n3992) );
  OR_GATE U4700 ( .I1(n3532), .I2(n3537), .O(n3535) );
  OR_GATE U4701 ( .I1(n3536), .I2(n3533), .O(n3534) );
  AND_GATE U4702 ( .I1(n3535), .I2(n3534), .O(n3542) );
  NAND_GATE U4703 ( .I1(n3537), .I2(n223), .O(n3539) );
  NAND3_GATE U4704 ( .I1(n3540), .I2(n3539), .I3(n3538), .O(n3541) );
  NAND_GATE U4705 ( .I1(n3542), .I2(n3541), .O(n3982) );
  NAND_GATE U4706 ( .I1(B[25]), .I2(A[15]), .O(n3985) );
  INV_GATE U4707 ( .I1(n3985), .O(n3980) );
  NAND_GATE U4708 ( .I1(n799), .I2(n3980), .O(n3977) );
  INV_GATE U4709 ( .I1(n3543), .O(n3547) );
  NAND_GATE U4710 ( .I1(n3547), .I2(n818), .O(n3545) );
  NAND_GATE U4711 ( .I1(n3543), .I2(n1310), .O(n3544) );
  NAND3_GATE U4712 ( .I1(n3546), .I2(n3545), .I3(n3544), .O(n3550) );
  NAND3_GATE U4713 ( .I1(n3548), .I2(n818), .I3(n3547), .O(n3549) );
  NAND_GATE U4714 ( .I1(n3550), .I2(n3549), .O(n3551) );
  NAND_GATE U4715 ( .I1(B[25]), .I2(A[14]), .O(n3970) );
  INV_GATE U4716 ( .I1(n3970), .O(n3965) );
  NAND_GATE U4717 ( .I1(n1296), .I2(n3965), .O(n3966) );
  NAND_GATE U4718 ( .I1(n3551), .I2(n3970), .O(n3723) );
  NAND_GATE U4719 ( .I1(n803), .I2(n3970), .O(n3722) );
  OR_GATE U4720 ( .I1(n3552), .I2(n3558), .O(n3555) );
  OR_GATE U4721 ( .I1(n3553), .I2(n3557), .O(n3554) );
  AND_GATE U4722 ( .I1(n3555), .I2(n3554), .O(n3563) );
  INV_GATE U4723 ( .I1(n3558), .O(n3556) );
  NAND_GATE U4724 ( .I1(n3557), .I2(n3556), .O(n3561) );
  NAND_GATE U4725 ( .I1(n8), .I2(n3558), .O(n3560) );
  NAND3_GATE U4726 ( .I1(n3561), .I2(n3560), .I3(n3559), .O(n3562) );
  NAND_GATE U4727 ( .I1(n3563), .I2(n3562), .O(n3948) );
  NAND_GATE U4728 ( .I1(B[25]), .I2(A[13]), .O(n3954) );
  INV_GATE U4729 ( .I1(n3954), .O(n3949) );
  NAND_GATE U4730 ( .I1(n3944), .I2(n3949), .O(n3950) );
  NAND3_GATE U4731 ( .I1(n3566), .I2(n3565), .I3(n3564), .O(n3573) );
  OR_GATE U4732 ( .I1(n3568), .I2(n3567), .O(n3572) );
  OR_GATE U4733 ( .I1(n3570), .I2(n3569), .O(n3571) );
  NAND3_GATE U4734 ( .I1(n3573), .I2(n3572), .I3(n3571), .O(n3936) );
  NAND_GATE U4735 ( .I1(B[25]), .I2(A[12]), .O(n3934) );
  INV_GATE U4736 ( .I1(n3934), .O(n3932) );
  NAND_GATE U4737 ( .I1(n780), .I2(n3932), .O(n3929) );
  NAND_GATE U4738 ( .I1(B[25]), .I2(A[11]), .O(n4447) );
  INV_GATE U4739 ( .I1(n4447), .O(n3791) );
  OR_GATE U4740 ( .I1(n3578), .I2(n3574), .O(n3577) );
  NAND3_GATE U4741 ( .I1(n235), .I2(n3575), .I3(n3578), .O(n3576) );
  AND_GATE U4742 ( .I1(n3577), .I2(n3576), .O(n3584) );
  NAND_GATE U4743 ( .I1(n3578), .I2(n235), .O(n3581) );
  NAND3_GATE U4744 ( .I1(n3582), .I2(n3581), .I3(n3580), .O(n3583) );
  NAND_GATE U4745 ( .I1(n3584), .I2(n3583), .O(n3787) );
  NAND_GATE U4746 ( .I1(n3791), .I2(n610), .O(n3717) );
  NAND_GATE U4747 ( .I1(B[25]), .I2(A[10]), .O(n3794) );
  NAND_GATE U4748 ( .I1(n3587), .I2(n1034), .O(n3708) );
  NAND4_GATE U4749 ( .I1(n3709), .I2(n3794), .I3(n3708), .I4(n3710), .O(n3707)
         );
  OR_GATE U4750 ( .I1(n3587), .I2(n3586), .O(n3590) );
  NAND3_GATE U4751 ( .I1(n1034), .I2(n3588), .I3(n3587), .O(n3589) );
  NAND_GATE U4752 ( .I1(n3590), .I2(n3589), .O(n3711) );
  NAND_GATE U4753 ( .I1(n3794), .I2(n3711), .O(n3706) );
  INV_GATE U4754 ( .I1(n3660), .O(n3656) );
  NAND3_GATE U4755 ( .I1(n3591), .I2(n3656), .I3(n3657), .O(n3812) );
  NAND3_GATE U4756 ( .I1(n3591), .I2(n3660), .I3(n620), .O(n3813) );
  NAND_GATE U4757 ( .I1(B[25]), .I2(A[5]), .O(n3886) );
  INV_GATE U4758 ( .I1(n3886), .O(n3876) );
  NAND3_GATE U4759 ( .I1(n3593), .I2(n3592), .I3(n3600), .O(n3594) );
  NAND_GATE U4760 ( .I1(n3595), .I2(n3594), .O(n3831) );
  INV_GATE U4761 ( .I1(n3831), .O(n3596) );
  NAND3_GATE U4762 ( .I1(n3598), .I2(n3595), .I3(n3597), .O(n3826) );
  NAND_GATE U4763 ( .I1(n3596), .I2(n3826), .O(n3610) );
  NAND3_GATE U4764 ( .I1(n3598), .I2(n3599), .I3(n3597), .O(n3602) );
  NAND3_GATE U4765 ( .I1(n3600), .I2(n3599), .I3(n744), .O(n3601) );
  AND_GATE U4766 ( .I1(n3602), .I2(n3601), .O(n3833) );
  NAND3_GATE U4767 ( .I1(B[25]), .I2(B[26]), .I3(n1196), .O(n3842) );
  INV_GATE U4768 ( .I1(n3842), .O(n3846) );
  NAND_GATE U4769 ( .I1(n1393), .I2(A[1]), .O(n3603) );
  NAND_GATE U4770 ( .I1(n14784), .I2(n3603), .O(n3604) );
  NAND_GATE U4771 ( .I1(B[26]), .I2(n3604), .O(n3837) );
  NAND_GATE U4772 ( .I1(B[25]), .I2(A[2]), .O(n3845) );
  NAND_GATE U4773 ( .I1(n3837), .I2(n3845), .O(n3605) );
  NAND_GATE U4774 ( .I1(n3846), .I2(n3605), .O(n3609) );
  INV_GATE U4775 ( .I1(n3845), .O(n3840) );
  NAND_GATE U4776 ( .I1(n1392), .I2(A[0]), .O(n3606) );
  NAND_GATE U4777 ( .I1(n14781), .I2(n3606), .O(n3607) );
  NAND_GATE U4778 ( .I1(B[27]), .I2(n3607), .O(n3838) );
  NAND_GATE U4779 ( .I1(n3837), .I2(n3838), .O(n3844) );
  NAND_GATE U4780 ( .I1(n3840), .I2(n3844), .O(n3608) );
  NAND_GATE U4781 ( .I1(n3609), .I2(n3608), .O(n3825) );
  NAND3_GATE U4782 ( .I1(n3610), .I2(n3833), .I3(n3825), .O(n3612) );
  NAND_GATE U4783 ( .I1(B[25]), .I2(A[3]), .O(n3828) );
  INV_GATE U4784 ( .I1(n3828), .O(n3832) );
  NAND3_GATE U4785 ( .I1(n3832), .I2(n3831), .I3(n3833), .O(n3611) );
  NAND_GATE U4786 ( .I1(n3832), .I2(n3825), .O(n3829) );
  NAND3_GATE U4787 ( .I1(n3612), .I2(n3611), .I3(n3829), .O(n3820) );
  NAND_GATE U4788 ( .I1(B[25]), .I2(A[4]), .O(n4493) );
  INV_GATE U4789 ( .I1(n3621), .O(n3619) );
  NAND4_GATE U4790 ( .I1(n3615), .I2(n3614), .I3(n3619), .I4(n3613), .O(n3627)
         );
  NAND_GATE U4791 ( .I1(n3615), .I2(n3614), .O(n3616) );
  NAND_GATE U4792 ( .I1(n3617), .I2(n3616), .O(n3620) );
  OR_GATE U4793 ( .I1(n3620), .I2(n3618), .O(n3626) );
  NAND_GATE U4794 ( .I1(n3619), .I2(n3620), .O(n3623) );
  NAND3_GATE U4795 ( .I1(n3624), .I2(n3623), .I3(n3622), .O(n3625) );
  NAND3_GATE U4796 ( .I1(n3627), .I2(n3626), .I3(n3625), .O(n3821) );
  NAND_GATE U4797 ( .I1(n4493), .I2(n3821), .O(n3628) );
  NAND_GATE U4798 ( .I1(n3820), .I2(n3628), .O(n3630) );
  INV_GATE U4799 ( .I1(n4493), .O(n4491) );
  NAND_GATE U4800 ( .I1(n4491), .I2(n767), .O(n3629) );
  NAND_GATE U4801 ( .I1(n3630), .I2(n3629), .O(n3880) );
  NAND_GATE U4802 ( .I1(n3876), .I2(n3880), .O(n3874) );
  NAND_GATE U4803 ( .I1(n3632), .I2(n573), .O(n3631) );
  INV_GATE U4804 ( .I1(n3632), .O(n3638) );
  NAND_GATE U4805 ( .I1(n3631), .I2(n3868), .O(n3870) );
  NAND3_GATE U4806 ( .I1(n3637), .I2(n3876), .I3(n3638), .O(n3635) );
  NAND3_GATE U4807 ( .I1(n1182), .I2(n3876), .I3(n573), .O(n3634) );
  NAND_GATE U4808 ( .I1(n3871), .I2(n3876), .O(n3633) );
  NAND3_GATE U4809 ( .I1(n3635), .I2(n3634), .I3(n3633), .O(n3636) );
  NAND_GATE U4810 ( .I1(n3872), .I2(n3636), .O(n3640) );
  NAND_GATE U4811 ( .I1(n3638), .I2(n3637), .O(n3868) );
  NAND_GATE U4812 ( .I1(n573), .I2(n1182), .O(n3875) );
  NAND3_GATE U4813 ( .I1(n3868), .I2(n3875), .I3(n3869), .O(n3882) );
  NAND3_GATE U4814 ( .I1(n3880), .I2(n3882), .I3(n3872), .O(n3639) );
  NAND3_GATE U4815 ( .I1(n3874), .I2(n3640), .I3(n3639), .O(n3892) );
  NAND_GATE U4816 ( .I1(n3645), .I2(n3649), .O(n3642) );
  NAND3_GATE U4817 ( .I1(n3644), .I2(n3643), .I3(n3642), .O(n3652) );
  NAND4_GATE U4818 ( .I1(n3647), .I2(n3646), .I3(n1153), .I4(n3645), .O(n3651)
         );
  OR_GATE U4819 ( .I1(n3649), .I2(n3648), .O(n3650) );
  NAND3_GATE U4820 ( .I1(n3652), .I2(n3651), .I3(n3650), .O(n3893) );
  NAND_GATE U4821 ( .I1(B[25]), .I2(A[6]), .O(n4567) );
  NAND_GATE U4822 ( .I1(n3893), .I2(n4567), .O(n3653) );
  NAND_GATE U4823 ( .I1(n3892), .I2(n3653), .O(n3655) );
  INV_GATE U4824 ( .I1(n4567), .O(n4561) );
  NAND_GATE U4825 ( .I1(n814), .I2(n4561), .O(n3654) );
  NAND_GATE U4826 ( .I1(n3655), .I2(n3654), .O(n3819) );
  AND3_GATE U4827 ( .I1(n3812), .I2(n3813), .I3(n3819), .O(n3659) );
  NAND_GATE U4828 ( .I1(n3657), .I2(n3656), .O(n3810) );
  NAND3_GATE U4829 ( .I1(n3811), .I2(n3660), .I3(n620), .O(n3816) );
  NAND3_GATE U4830 ( .I1(n3810), .I2(n3816), .I3(n3811), .O(n3658) );
  NAND_GATE U4831 ( .I1(n3659), .I2(n3658), .O(n3666) );
  NAND_GATE U4832 ( .I1(B[25]), .I2(A[7]), .O(n3900) );
  OR_GATE U4833 ( .I1(n3816), .I2(n3900), .O(n3663) );
  NAND_GATE U4834 ( .I1(n3811), .I2(n3660), .O(n3805) );
  INV_GATE U4835 ( .I1(n3900), .O(n3808) );
  NAND3_GATE U4836 ( .I1(n3661), .I2(n861), .I3(n3811), .O(n3804) );
  NAND3_GATE U4837 ( .I1(n3805), .I2(n3808), .I3(n3804), .O(n3662) );
  NAND_GATE U4838 ( .I1(n3663), .I2(n3662), .O(n3664) );
  NAND_GATE U4839 ( .I1(n1154), .I2(n3664), .O(n3665) );
  NAND_GATE U4840 ( .I1(n3808), .I2(n3819), .O(n3809) );
  NAND3_GATE U4841 ( .I1(n3666), .I2(n3665), .I3(n3809), .O(n3909) );
  NAND_GATE U4842 ( .I1(B[25]), .I2(A[8]), .O(n4472) );
  INV_GATE U4843 ( .I1(n3667), .O(n3671) );
  NAND_GATE U4844 ( .I1(n3672), .I2(n3671), .O(n3679) );
  NAND4_GATE U4845 ( .I1(n3678), .I2(n4472), .I3(n3680), .I4(n3679), .O(n3675)
         );
  NAND3_GATE U4846 ( .I1(n3672), .I2(n3671), .I3(n3670), .O(n3676) );
  NAND_GATE U4847 ( .I1(n3677), .I2(n3676), .O(n3673) );
  NAND_GATE U4848 ( .I1(n4472), .I2(n3673), .O(n3674) );
  NAND3_GATE U4849 ( .I1(n3909), .I2(n3675), .I3(n3674), .O(n3682) );
  INV_GATE U4850 ( .I1(n4472), .O(n4465) );
  NAND3_GATE U4851 ( .I1(n3680), .I2(n3679), .I3(n3678), .O(n3904) );
  NAND_GATE U4852 ( .I1(n1139), .I2(n3904), .O(n4463) );
  NAND_GATE U4853 ( .I1(n4465), .I2(n3908), .O(n3681) );
  NAND_GATE U4854 ( .I1(n3682), .I2(n3681), .O(n3915) );
  NAND_GATE U4855 ( .I1(B[25]), .I2(A[9]), .O(n3913) );
  INV_GATE U4856 ( .I1(n3683), .O(n3694) );
  NAND_GATE U4857 ( .I1(n3692), .I2(n3694), .O(n3699) );
  INV_GATE U4858 ( .I1(n3692), .O(n3689) );
  NAND_GATE U4859 ( .I1(n3689), .I2(n3683), .O(n3701) );
  NAND4_GATE U4860 ( .I1(n3700), .I2(n3913), .I3(n3699), .I4(n3701), .O(n3698)
         );
  NAND3_GATE U4861 ( .I1(n3686), .I2(n3685), .I3(n3684), .O(n3691) );
  AND_GATE U4862 ( .I1(n3688), .I2(n3687), .O(n3690) );
  NAND4_GATE U4863 ( .I1(n3693), .I2(n3691), .I3(n3690), .I4(n3689), .O(n3696)
         );
  NAND3_GATE U4864 ( .I1(n3694), .I2(n3693), .I3(n3692), .O(n3695) );
  NAND_GATE U4865 ( .I1(n3696), .I2(n3695), .O(n3702) );
  NAND_GATE U4866 ( .I1(n3913), .I2(n3702), .O(n3697) );
  NAND3_GATE U4867 ( .I1(n3915), .I2(n3698), .I3(n3697), .O(n3705) );
  INV_GATE U4868 ( .I1(n3913), .O(n3919) );
  AND3_GATE U4869 ( .I1(n3701), .I2(n3700), .I3(n3699), .O(n3703) );
  NAND_GATE U4870 ( .I1(n3919), .I2(n1263), .O(n3704) );
  NAND_GATE U4871 ( .I1(n3705), .I2(n3704), .O(n3793) );
  NAND3_GATE U4872 ( .I1(n3707), .I2(n3706), .I3(n3793), .O(n3714) );
  INV_GATE U4873 ( .I1(n3794), .O(n3798) );
  AND3_GATE U4874 ( .I1(n3710), .I2(n3709), .I3(n3708), .O(n3712) );
  NAND_GATE U4875 ( .I1(n3798), .I2(n1303), .O(n3713) );
  NAND_GATE U4876 ( .I1(n3714), .I2(n3713), .O(n3790) );
  NAND_GATE U4877 ( .I1(n4447), .I2(n3787), .O(n3715) );
  NAND_GATE U4878 ( .I1(n3790), .I2(n3715), .O(n3716) );
  NAND_GATE U4879 ( .I1(n3717), .I2(n3716), .O(n3933) );
  NAND_GATE U4880 ( .I1(n3936), .I2(n3934), .O(n3718) );
  NAND_GATE U4881 ( .I1(n3933), .I2(n3718), .O(n3719) );
  NAND_GATE U4882 ( .I1(n3929), .I2(n3719), .O(n3951) );
  NAND_GATE U4883 ( .I1(n3948), .I2(n3954), .O(n3720) );
  NAND_GATE U4884 ( .I1(n3951), .I2(n3720), .O(n3721) );
  NAND_GATE U4885 ( .I1(n3950), .I2(n3721), .O(n3967) );
  NAND3_GATE U4886 ( .I1(n3723), .I2(n3722), .I3(n3967), .O(n3724) );
  NAND_GATE U4887 ( .I1(n3966), .I2(n3724), .O(n3981) );
  NAND_GATE U4888 ( .I1(n3982), .I2(n3985), .O(n3725) );
  NAND_GATE U4889 ( .I1(n3981), .I2(n3725), .O(n3726) );
  NAND_GATE U4890 ( .I1(n3977), .I2(n3726), .O(n3996) );
  NAND_GATE U4891 ( .I1(n3997), .I2(n4000), .O(n3727) );
  NAND_GATE U4892 ( .I1(n3996), .I2(n3727), .O(n3728) );
  NAND_GATE U4893 ( .I1(n3992), .I2(n3728), .O(n4011) );
  NAND_GATE U4894 ( .I1(n4009), .I2(n4016), .O(n3729) );
  NAND_GATE U4895 ( .I1(n4011), .I2(n3729), .O(n3730) );
  NAND_GATE U4896 ( .I1(n4007), .I2(n3730), .O(n4027) );
  NAND_GATE U4897 ( .I1(n4025), .I2(n4032), .O(n3731) );
  NAND_GATE U4898 ( .I1(n4027), .I2(n3731), .O(n3732) );
  NAND_GATE U4899 ( .I1(n4023), .I2(n3732), .O(n4043) );
  NAND_GATE U4900 ( .I1(n4041), .I2(n4048), .O(n3733) );
  NAND_GATE U4901 ( .I1(n4043), .I2(n3733), .O(n3734) );
  NAND_GATE U4902 ( .I1(n4039), .I2(n3734), .O(n4059) );
  NAND_GATE U4903 ( .I1(n4057), .I2(n4064), .O(n3735) );
  NAND_GATE U4904 ( .I1(n4059), .I2(n3735), .O(n3736) );
  NAND_GATE U4905 ( .I1(n4055), .I2(n3736), .O(n4075) );
  NAND_GATE U4906 ( .I1(n4073), .I2(n4080), .O(n3737) );
  NAND_GATE U4907 ( .I1(n4075), .I2(n3737), .O(n3738) );
  NAND_GATE U4908 ( .I1(n4071), .I2(n3738), .O(n4091) );
  NAND_GATE U4909 ( .I1(n4089), .I2(n4096), .O(n3739) );
  NAND_GATE U4910 ( .I1(n4091), .I2(n3739), .O(n3740) );
  NAND_GATE U4911 ( .I1(n4087), .I2(n3740), .O(n4108) );
  NAND_GATE U4912 ( .I1(n4106), .I2(n4113), .O(n3741) );
  NAND_GATE U4913 ( .I1(n4108), .I2(n3741), .O(n3742) );
  NAND_GATE U4914 ( .I1(n4103), .I2(n3742), .O(n3777) );
  NAND_GATE U4915 ( .I1(n3775), .I2(n3782), .O(n3743) );
  NAND_GATE U4916 ( .I1(n3777), .I2(n3743), .O(n3744) );
  NAND_GATE U4917 ( .I1(n3772), .I2(n3744), .O(n4127) );
  NAND_GATE U4918 ( .I1(n4125), .I2(n4132), .O(n3745) );
  NAND_GATE U4919 ( .I1(n4127), .I2(n3745), .O(n3746) );
  NAND_GATE U4920 ( .I1(n4122), .I2(n3746), .O(n4144) );
  NAND_GATE U4921 ( .I1(n4142), .I2(n4144), .O(n4139) );
  OR_GATE U4922 ( .I1(n3747), .I2(n3752), .O(n3750) );
  OR_GATE U4923 ( .I1(n3751), .I2(n3748), .O(n3749) );
  AND_GATE U4924 ( .I1(n3750), .I2(n3749), .O(n3757) );
  NAND_GATE U4925 ( .I1(n3752), .I2(n1110), .O(n3754) );
  NAND3_GATE U4926 ( .I1(n3755), .I2(n3754), .I3(n3753), .O(n3756) );
  NAND_GATE U4927 ( .I1(n3757), .I2(n3756), .O(n4140) );
  INV_GATE U4928 ( .I1(n4140), .O(n4143) );
  INV_GATE U4929 ( .I1(n4144), .O(n4141) );
  NAND_GATE U4930 ( .I1(n4148), .I2(n4141), .O(n3758) );
  NAND_GATE U4931 ( .I1(n4143), .I2(n3758), .O(n3759) );
  NAND_GATE U4932 ( .I1(n4139), .I2(n3759), .O(n4159) );
  NAND_GATE U4933 ( .I1(n4157), .I2(n4164), .O(n3760) );
  NAND_GATE U4934 ( .I1(n4159), .I2(n3760), .O(n3761) );
  NAND_GATE U4935 ( .I1(n4155), .I2(n3761), .O(n4175) );
  NAND_GATE U4936 ( .I1(n4173), .I2(n4180), .O(n3762) );
  NAND_GATE U4937 ( .I1(n4175), .I2(n3762), .O(n3763) );
  NAND_GATE U4938 ( .I1(n4171), .I2(n3763), .O(n4191) );
  NAND_GATE U4939 ( .I1(n4189), .I2(n4196), .O(n3764) );
  NAND_GATE U4940 ( .I1(n4191), .I2(n3764), .O(n3765) );
  NAND_GATE U4941 ( .I1(n4187), .I2(n3765), .O(n4207) );
  NAND_GATE U4942 ( .I1(n4205), .I2(n4212), .O(n3766) );
  NAND_GATE U4943 ( .I1(n4207), .I2(n3766), .O(n3767) );
  NAND_GATE U4944 ( .I1(n4203), .I2(n3767), .O(n4223) );
  NAND_GATE U4945 ( .I1(n4221), .I2(n4228), .O(n3768) );
  NAND_GATE U4946 ( .I1(n4223), .I2(n3768), .O(n3769) );
  NAND_GATE U4947 ( .I1(n4219), .I2(n3769), .O(n3770) );
  NAND_GATE U4948 ( .I1(n287), .I2(n3770), .O(n15313) );
  AND_GATE U4949 ( .I1(n15313), .I2(n3771), .O(\A1[55] ) );
  NAND_GATE U4950 ( .I1(B[24]), .I2(A[31]), .O(n4243) );
  INV_GATE U4951 ( .I1(n4243), .O(n4217) );
  NAND_GATE U4952 ( .I1(B[24]), .I2(A[30]), .O(n4254) );
  INV_GATE U4953 ( .I1(n4254), .O(n4201) );
  NAND_GATE U4954 ( .I1(B[24]), .I2(A[29]), .O(n4265) );
  INV_GATE U4955 ( .I1(n4265), .O(n4185) );
  NAND_GATE U4956 ( .I1(B[24]), .I2(A[28]), .O(n4276) );
  INV_GATE U4957 ( .I1(n4276), .O(n4169) );
  NAND_GATE U4958 ( .I1(B[24]), .I2(A[27]), .O(n4287) );
  INV_GATE U4959 ( .I1(n4287), .O(n4153) );
  NAND_GATE U4960 ( .I1(B[24]), .I2(A[26]), .O(n4298) );
  INV_GATE U4961 ( .I1(n4298), .O(n4137) );
  NAND_GATE U4962 ( .I1(B[24]), .I2(A[25]), .O(n4309) );
  INV_GATE U4963 ( .I1(n4309), .O(n4120) );
  INV_GATE U4964 ( .I1(n3772), .O(n3773) );
  NAND_GATE U4965 ( .I1(n3773), .I2(n3777), .O(n3786) );
  INV_GATE U4966 ( .I1(n3777), .O(n3774) );
  NAND_GATE U4967 ( .I1(n3775), .I2(n3774), .O(n3780) );
  NAND_GATE U4968 ( .I1(n3776), .I2(n3780), .O(n3784) );
  NAND_GATE U4969 ( .I1(n3778), .I2(n3777), .O(n3779) );
  NAND_GATE U4970 ( .I1(n3780), .I2(n3779), .O(n3781) );
  NAND_GATE U4971 ( .I1(n3782), .I2(n3781), .O(n3783) );
  NAND_GATE U4972 ( .I1(n3784), .I2(n3783), .O(n3785) );
  NAND_GATE U4973 ( .I1(n3786), .I2(n3785), .O(n4307) );
  NAND_GATE U4974 ( .I1(n4120), .I2(n4307), .O(n4304) );
  NAND_GATE U4975 ( .I1(B[24]), .I2(A[24]), .O(n4320) );
  INV_GATE U4976 ( .I1(n4320), .O(n4118) );
  NAND_GATE U4977 ( .I1(B[24]), .I2(A[23]), .O(n4678) );
  INV_GATE U4978 ( .I1(n4678), .O(n4101) );
  NAND_GATE U4979 ( .I1(B[24]), .I2(A[22]), .O(n4331) );
  INV_GATE U4980 ( .I1(n4331), .O(n4085) );
  NAND_GATE U4981 ( .I1(B[24]), .I2(A[21]), .O(n4344) );
  INV_GATE U4982 ( .I1(n4344), .O(n4069) );
  NAND_GATE U4983 ( .I1(B[24]), .I2(A[20]), .O(n4357) );
  INV_GATE U4984 ( .I1(n4357), .O(n4053) );
  NAND_GATE U4985 ( .I1(B[24]), .I2(A[19]), .O(n4370) );
  INV_GATE U4986 ( .I1(n4370), .O(n4037) );
  NAND_GATE U4987 ( .I1(B[24]), .I2(A[18]), .O(n4382) );
  INV_GATE U4988 ( .I1(n4382), .O(n4021) );
  NAND_GATE U4989 ( .I1(B[24]), .I2(A[17]), .O(n4393) );
  INV_GATE U4990 ( .I1(n4393), .O(n4005) );
  NAND_GATE U4991 ( .I1(B[24]), .I2(A[16]), .O(n4403) );
  INV_GATE U4992 ( .I1(n4403), .O(n3990) );
  NAND_GATE U4993 ( .I1(B[24]), .I2(A[15]), .O(n4418) );
  INV_GATE U4994 ( .I1(n4418), .O(n3968) );
  NAND_GATE U4995 ( .I1(B[24]), .I2(A[14]), .O(n4429) );
  INV_GATE U4996 ( .I1(n4429), .O(n3952) );
  NAND_GATE U4997 ( .I1(B[24]), .I2(A[13]), .O(n4441) );
  INV_GATE U4998 ( .I1(n4441), .O(n3942) );
  NAND_GATE U4999 ( .I1(B[24]), .I2(A[12]), .O(n4455) );
  INV_GATE U5000 ( .I1(n4455), .O(n3927) );
  NAND_GATE U5001 ( .I1(n3791), .I2(n3789), .O(n4448) );
  NAND_GATE U5002 ( .I1(n3787), .I2(n616), .O(n3789) );
  NAND_GATE U5003 ( .I1(n610), .I2(n3790), .O(n3788) );
  NAND_GATE U5004 ( .I1(n3789), .I2(n3788), .O(n4446) );
  NAND_GATE U5005 ( .I1(n4448), .I2(n4451), .O(n3792) );
  NAND3_GATE U5006 ( .I1(n3791), .I2(n3790), .I3(n610), .O(n4449) );
  NAND_GATE U5007 ( .I1(n3792), .I2(n4449), .O(n4456) );
  NAND_GATE U5008 ( .I1(n3927), .I2(n4456), .O(n4458) );
  NAND_GATE U5009 ( .I1(B[24]), .I2(A[11]), .O(n4641) );
  INV_GATE U5010 ( .I1(n4641), .O(n4631) );
  NAND3_GATE U5011 ( .I1(n3793), .I2(n3798), .I3(n1303), .O(n3803) );
  NAND3_GATE U5012 ( .I1(n3798), .I2(n3797), .I3(n3803), .O(n3796) );
  NAND3_GATE U5013 ( .I1(n3793), .I2(n3794), .I3(n1303), .O(n3801) );
  AND_GATE U5014 ( .I1(n3801), .I2(n3800), .O(n3795) );
  NAND3_GATE U5015 ( .I1(n4631), .I2(n3796), .I3(n3795), .O(n4632) );
  NAND_GATE U5016 ( .I1(n3798), .I2(n3797), .O(n3799) );
  NAND3_GATE U5017 ( .I1(n3801), .I2(n3800), .I3(n3799), .O(n3802) );
  NAND_GATE U5018 ( .I1(n3803), .I2(n3802), .O(n4636) );
  NAND_GATE U5019 ( .I1(B[24]), .I2(A[10]), .O(n4623) );
  INV_GATE U5020 ( .I1(n4623), .O(n4615) );
  NAND_GATE U5021 ( .I1(B[24]), .I2(A[9]), .O(n4600) );
  INV_GATE U5022 ( .I1(n4600), .O(n4608) );
  NAND_GATE U5023 ( .I1(B[24]), .I2(A[8]), .O(n4585) );
  INV_GATE U5024 ( .I1(n4585), .O(n4590) );
  NAND_GATE U5025 ( .I1(n3805), .I2(n3804), .O(n3806) );
  NAND_GATE U5026 ( .I1(n3816), .I2(n3806), .O(n3807) );
  INV_GATE U5027 ( .I1(n3819), .O(n3818) );
  NAND4_GATE U5028 ( .I1(n3808), .I2(n3807), .I3(n1154), .I4(n3818), .O(n4583)
         );
  NAND_GATE U5029 ( .I1(n3811), .I2(n3810), .O(n3814) );
  NAND3_GATE U5030 ( .I1(n3814), .I2(n3813), .I3(n3812), .O(n3815) );
  NAND_GATE U5031 ( .I1(n3816), .I2(n3815), .O(n3817) );
  NAND_GATE U5032 ( .I1(n4583), .I2(n4582), .O(n3901) );
  INV_GATE U5033 ( .I1(n3901), .O(n4581) );
  NAND_GATE U5034 ( .I1(n3818), .I2(n3817), .O(n3899) );
  NAND_GATE U5035 ( .I1(n4590), .I2(n1311), .O(n4469) );
  NAND_GATE U5036 ( .I1(B[24]), .I2(A[7]), .O(n4574) );
  INV_GATE U5037 ( .I1(n4574), .O(n4560) );
  INV_GATE U5038 ( .I1(n3820), .O(n3822) );
  NAND_GATE U5039 ( .I1(n3822), .I2(n3821), .O(n4490) );
  NAND3_GATE U5040 ( .I1(n3820), .I2(n4491), .I3(n767), .O(n4488) );
  NAND3_GATE U5041 ( .I1(n4490), .I2(n4488), .I3(n4491), .O(n4498) );
  NAND_GATE U5042 ( .I1(n3820), .I2(n767), .O(n3823) );
  NAND_GATE U5043 ( .I1(n3823), .I2(n4490), .O(n4492) );
  INV_GATE U5044 ( .I1(n3825), .O(n3834) );
  NAND_GATE U5045 ( .I1(n3833), .I2(n3831), .O(n3824) );
  NAND_GATE U5046 ( .I1(n3826), .I2(n3824), .O(n3830) );
  NAND_GATE U5047 ( .I1(n3834), .I2(n3830), .O(n3860) );
  NAND3_GATE U5048 ( .I1(n3826), .I2(n3825), .I3(n3824), .O(n3827) );
  AND_GATE U5049 ( .I1(n3828), .I2(n3827), .O(n3861) );
  NAND_GATE U5050 ( .I1(B[24]), .I2(A[4]), .O(n4734) );
  NAND3_GATE U5051 ( .I1(n3860), .I2(n3861), .I3(n4734), .O(n3859) );
  OR_GATE U5052 ( .I1(n3830), .I2(n3829), .O(n3836) );
  NAND4_GATE U5053 ( .I1(n3834), .I2(n3833), .I3(n3832), .I4(n3831), .O(n3835)
         );
  NAND_GATE U5054 ( .I1(n3836), .I2(n3835), .O(n3862) );
  NAND_GATE U5055 ( .I1(n4734), .I2(n3862), .O(n3858) );
  NAND3_GATE U5056 ( .I1(n3838), .I2(n3837), .I3(n3842), .O(n3839) );
  NAND_GATE U5057 ( .I1(n3840), .I2(n3839), .O(n4534) );
  INV_GATE U5058 ( .I1(n4534), .O(n3841) );
  NAND3_GATE U5059 ( .I1(n3846), .I2(n3840), .I3(n3844), .O(n4531) );
  NAND_GATE U5060 ( .I1(n3841), .I2(n4531), .O(n3855) );
  NAND_GATE U5061 ( .I1(n3842), .I2(n3845), .O(n3843) );
  OR_GATE U5062 ( .I1(n3843), .I2(n3844), .O(n3848) );
  NAND3_GATE U5063 ( .I1(n3846), .I2(n3845), .I3(n3844), .O(n3847) );
  AND_GATE U5064 ( .I1(n3848), .I2(n3847), .O(n4533) );
  NAND_GATE U5065 ( .I1(B[24]), .I2(A[2]), .O(n4514) );
  INV_GATE U5066 ( .I1(n4514), .O(n4510) );
  NAND_GATE U5067 ( .I1(n1392), .I2(A[1]), .O(n3849) );
  NAND_GATE U5068 ( .I1(n14784), .I2(n3849), .O(n3850) );
  NAND_GATE U5069 ( .I1(B[25]), .I2(n3850), .O(n4507) );
  NAND_GATE U5070 ( .I1(n1391), .I2(A[0]), .O(n3851) );
  NAND_GATE U5071 ( .I1(n14781), .I2(n3851), .O(n3852) );
  NAND_GATE U5072 ( .I1(B[26]), .I2(n3852), .O(n4508) );
  NAND_GATE U5073 ( .I1(n4507), .I2(n4508), .O(n4512) );
  NAND_GATE U5074 ( .I1(n4510), .I2(n4512), .O(n4518) );
  NAND3_GATE U5075 ( .I1(B[24]), .I2(B[25]), .I3(n1196), .O(n4519) );
  INV_GATE U5076 ( .I1(n4519), .O(n4511) );
  INV_GATE U5077 ( .I1(n4512), .O(n4513) );
  NAND_GATE U5078 ( .I1(n4514), .I2(n4513), .O(n3853) );
  NAND_GATE U5079 ( .I1(n4511), .I2(n3853), .O(n3854) );
  NAND_GATE U5080 ( .I1(n4518), .I2(n3854), .O(n4538) );
  NAND3_GATE U5081 ( .I1(n3855), .I2(n4533), .I3(n4538), .O(n3857) );
  NAND_GATE U5082 ( .I1(B[24]), .I2(A[3]), .O(n4541) );
  INV_GATE U5083 ( .I1(n4541), .O(n4535) );
  NAND3_GATE U5084 ( .I1(n4535), .I2(n4534), .I3(n4533), .O(n3856) );
  NAND_GATE U5085 ( .I1(n4535), .I2(n4538), .O(n4532) );
  NAND3_GATE U5086 ( .I1(n3857), .I2(n3856), .I3(n4532), .O(n4505) );
  NAND3_GATE U5087 ( .I1(n3859), .I2(n3858), .I3(n4505), .O(n3865) );
  INV_GATE U5088 ( .I1(n4734), .O(n4724) );
  AND_GATE U5089 ( .I1(n3861), .I2(n3860), .O(n3863) );
  NAND_GATE U5090 ( .I1(n4724), .I2(n820), .O(n3864) );
  NAND_GATE U5091 ( .I1(n3865), .I2(n3864), .O(n4486) );
  NAND3_GATE U5092 ( .I1(n4498), .I2(n4494), .I3(n4486), .O(n3867) );
  NAND_GATE U5093 ( .I1(B[24]), .I2(A[5]), .O(n4552) );
  INV_GATE U5094 ( .I1(n4552), .O(n4499) );
  NAND3_GATE U5095 ( .I1(n4499), .I2(n4498), .I3(n4494), .O(n3866) );
  NAND_GATE U5096 ( .I1(n4499), .I2(n4486), .O(n4487) );
  NAND3_GATE U5097 ( .I1(n3867), .I2(n3866), .I3(n4487), .O(n4482) );
  NAND_GATE U5098 ( .I1(B[24]), .I2(A[6]), .O(n4801) );
  NAND_GATE U5099 ( .I1(n3869), .I2(n3868), .O(n3873) );
  NAND_GATE U5100 ( .I1(n3871), .I2(n3870), .O(n3872) );
  INV_GATE U5101 ( .I1(n3880), .O(n3881) );
  NAND4_GATE U5102 ( .I1(n3876), .I2(n3882), .I3(n3881), .I4(n3872), .O(n3877)
         );
  NAND_GATE U5103 ( .I1(n3878), .I2(n3877), .O(n3888) );
  NAND_GATE U5104 ( .I1(n4801), .I2(n3888), .O(n3884) );
  NAND_GATE U5105 ( .I1(n3872), .I2(n3882), .O(n3879) );
  NAND_GATE U5106 ( .I1(n3880), .I2(n3879), .O(n3887) );
  NAND3_GATE U5107 ( .I1(n3872), .I2(n3882), .I3(n3881), .O(n3885) );
  NAND4_GATE U5108 ( .I1(n3886), .I2(n3887), .I3(n4801), .I4(n3885), .O(n3883)
         );
  NAND3_GATE U5109 ( .I1(n4482), .I2(n3884), .I3(n3883), .O(n3891) );
  INV_GATE U5110 ( .I1(n4801), .O(n4799) );
  AND3_GATE U5111 ( .I1(n3887), .I2(n3886), .I3(n3885), .O(n3889) );
  OR_GATE U5112 ( .I1(n3889), .I2(n3888), .O(n4483) );
  NAND_GATE U5113 ( .I1(n4799), .I2(n549), .O(n3890) );
  NAND_GATE U5114 ( .I1(n3891), .I2(n3890), .O(n4571) );
  NAND_GATE U5115 ( .I1(n4560), .I2(n4571), .O(n4563) );
  INV_GATE U5116 ( .I1(n3892), .O(n3894) );
  NAND_GATE U5117 ( .I1(n3892), .I2(n814), .O(n4565) );
  NAND_GATE U5118 ( .I1(n3894), .I2(n3893), .O(n3895) );
  NAND_GATE U5119 ( .I1(n4565), .I2(n3895), .O(n4566) );
  NAND_GATE U5120 ( .I1(n4567), .I2(n4566), .O(n4559) );
  NAND3_GATE U5121 ( .I1(n4560), .I2(n4569), .I3(n4559), .O(n3897) );
  NAND3_GATE U5122 ( .I1(n4569), .I2(n4559), .I3(n4571), .O(n3896) );
  NAND3_GATE U5123 ( .I1(n4563), .I2(n3897), .I3(n3896), .O(n4584) );
  NAND4_GATE U5124 ( .I1(n3900), .I2(n4585), .I3(n3899), .I4(n3898), .O(n3903)
         );
  NAND_GATE U5125 ( .I1(n4585), .I2(n3901), .O(n3902) );
  NAND3_GATE U5126 ( .I1(n4584), .I2(n3903), .I3(n3902), .O(n4468) );
  NAND_GATE U5127 ( .I1(n4469), .I2(n4468), .O(n4606) );
  NAND3_GATE U5128 ( .I1(n3908), .I2(n4465), .I3(n3909), .O(n4476) );
  NAND_GATE U5129 ( .I1(n3909), .I2(n4465), .O(n3906) );
  NAND3_GATE U5130 ( .I1(n3904), .I2(n1139), .I3(n4465), .O(n3905) );
  NAND_GATE U5131 ( .I1(n3906), .I2(n3905), .O(n3907) );
  NAND_GATE U5132 ( .I1(n4476), .I2(n3907), .O(n4607) );
  NAND_GATE U5133 ( .I1(n3909), .I2(n3908), .O(n3910) );
  NAND_GATE U5134 ( .I1(n4464), .I2(n3910), .O(n4471) );
  NAND3_GATE U5135 ( .I1(n4608), .I2(n4607), .I3(n4473), .O(n3912) );
  NAND3_GATE U5136 ( .I1(n4606), .I2(n4607), .I3(n4473), .O(n3911) );
  NAND3_GATE U5137 ( .I1(n4470), .I2(n3912), .I3(n3911), .O(n4620) );
  NAND_GATE U5138 ( .I1(n4615), .I2(n4620), .O(n3924) );
  NAND_GATE U5139 ( .I1(n3919), .I2(n3918), .O(n3914) );
  NAND3_GATE U5140 ( .I1(n3913), .I2(n1263), .I3(n3915), .O(n3921) );
  NAND3_GATE U5141 ( .I1(n3914), .I2(n3920), .I3(n3921), .O(n3916) );
  NAND3_GATE U5142 ( .I1(n3915), .I2(n3919), .I3(n1263), .O(n3917) );
  NAND_GATE U5143 ( .I1(n3916), .I2(n3917), .O(n4617) );
  NAND_GATE U5144 ( .I1(n4620), .I2(n4617), .O(n3923) );
  NAND3_GATE U5145 ( .I1(n3919), .I2(n3918), .I3(n3917), .O(n4614) );
  NAND3_GATE U5146 ( .I1(n4615), .I2(n4614), .I3(n1152), .O(n3922) );
  NAND3_GATE U5147 ( .I1(n3924), .I2(n3923), .I3(n3922), .O(n4637) );
  NAND_GATE U5148 ( .I1(n4636), .I2(n4637), .O(n3926) );
  NAND_GATE U5149 ( .I1(n4631), .I2(n4637), .O(n3925) );
  NAND3_GATE U5150 ( .I1(n4632), .I2(n3926), .I3(n3925), .O(n4459) );
  NAND_GATE U5151 ( .I1(n4456), .I2(n4459), .O(n3928) );
  NAND_GATE U5152 ( .I1(n3927), .I2(n4459), .O(n4457) );
  NAND3_GATE U5153 ( .I1(n4458), .I2(n3928), .I3(n4457), .O(n4440) );
  NAND_GATE U5154 ( .I1(n3942), .I2(n4440), .O(n4436) );
  INV_GATE U5155 ( .I1(n3929), .O(n3930) );
  NAND_GATE U5156 ( .I1(n3930), .I2(n3933), .O(n3941) );
  INV_GATE U5157 ( .I1(n3933), .O(n3935) );
  NAND_GATE U5158 ( .I1(n3932), .I2(n3931), .O(n3939) );
  NAND_GATE U5159 ( .I1(n780), .I2(n3933), .O(n3938) );
  NAND3_GATE U5160 ( .I1(n3936), .I2(n3935), .I3(n3934), .O(n3937) );
  NAND3_GATE U5161 ( .I1(n3939), .I2(n3938), .I3(n3937), .O(n3940) );
  NAND_GATE U5162 ( .I1(n3941), .I2(n3940), .O(n4439) );
  NAND_GATE U5163 ( .I1(n3942), .I2(n4439), .O(n4435) );
  NAND_GATE U5164 ( .I1(n4440), .I2(n4439), .O(n3943) );
  NAND3_GATE U5165 ( .I1(n4436), .I2(n4435), .I3(n3943), .O(n4425) );
  NAND_GATE U5166 ( .I1(n3952), .I2(n4425), .O(n4430) );
  NAND_GATE U5167 ( .I1(n3944), .I2(n3951), .O(n3946) );
  INV_GATE U5168 ( .I1(n3951), .O(n3947) );
  NAND_GATE U5169 ( .I1(n3948), .I2(n3947), .O(n3945) );
  NAND_GATE U5170 ( .I1(n3946), .I2(n3945), .O(n3953) );
  NAND_GATE U5171 ( .I1(n3954), .I2(n3953), .O(n4422) );
  NAND_GATE U5172 ( .I1(n3949), .I2(n3945), .O(n3956) );
  NAND3_GATE U5173 ( .I1(n4422), .I2(n4423), .I3(n3952), .O(n4421) );
  AND_GATE U5174 ( .I1(n4430), .I2(n4421), .O(n3960) );
  NAND_GATE U5175 ( .I1(n3956), .I2(n3955), .O(n3957) );
  NAND_GATE U5176 ( .I1(n3958), .I2(n3957), .O(n4431) );
  NAND_GATE U5177 ( .I1(n4425), .I2(n4431), .O(n3959) );
  NAND_GATE U5178 ( .I1(n3960), .I2(n3959), .O(n4413) );
  NAND_GATE U5179 ( .I1(n1296), .I2(n3967), .O(n3962) );
  INV_GATE U5180 ( .I1(n3967), .O(n3963) );
  NAND_GATE U5181 ( .I1(n3964), .I2(n3963), .O(n3961) );
  NAND_GATE U5182 ( .I1(n3962), .I2(n3961), .O(n3969) );
  NAND_GATE U5183 ( .I1(n3965), .I2(n3961), .O(n3972) );
  NAND3_GATE U5184 ( .I1(n3971), .I2(n4411), .I3(n3968), .O(n4407) );
  AND_GATE U5185 ( .I1(n4408), .I2(n4407), .O(n3976) );
  NAND_GATE U5186 ( .I1(n3970), .I2(n3969), .O(n3971) );
  NAND_GATE U5187 ( .I1(n3972), .I2(n3971), .O(n3973) );
  NAND_GATE U5188 ( .I1(n3974), .I2(n3973), .O(n4414) );
  NAND_GATE U5189 ( .I1(n4413), .I2(n4414), .O(n3975) );
  NAND_GATE U5190 ( .I1(n3976), .I2(n3975), .O(n4402) );
  NAND_GATE U5191 ( .I1(n3990), .I2(n4402), .O(n4398) );
  INV_GATE U5192 ( .I1(n3977), .O(n3978) );
  NAND_GATE U5193 ( .I1(n3978), .I2(n3981), .O(n3989) );
  NAND_GATE U5194 ( .I1(n3980), .I2(n3979), .O(n3987) );
  NAND_GATE U5195 ( .I1(n799), .I2(n3981), .O(n3983) );
  NAND_GATE U5196 ( .I1(n3983), .I2(n3979), .O(n3984) );
  NAND_GATE U5197 ( .I1(n3985), .I2(n3984), .O(n3986) );
  NAND_GATE U5198 ( .I1(n3987), .I2(n3986), .O(n3988) );
  NAND_GATE U5199 ( .I1(n3989), .I2(n3988), .O(n4401) );
  NAND_GATE U5200 ( .I1(n3990), .I2(n4401), .O(n4397) );
  NAND_GATE U5201 ( .I1(n4402), .I2(n4401), .O(n3991) );
  NAND3_GATE U5202 ( .I1(n4398), .I2(n4397), .I3(n3991), .O(n4392) );
  NAND_GATE U5203 ( .I1(n4005), .I2(n4392), .O(n4388) );
  INV_GATE U5204 ( .I1(n3992), .O(n3993) );
  NAND_GATE U5205 ( .I1(n3993), .I2(n3996), .O(n4004) );
  NAND_GATE U5206 ( .I1(n3995), .I2(n3994), .O(n4002) );
  NAND_GATE U5207 ( .I1(n399), .I2(n3996), .O(n3998) );
  NAND_GATE U5208 ( .I1(n3998), .I2(n3994), .O(n3999) );
  NAND_GATE U5209 ( .I1(n4000), .I2(n3999), .O(n4001) );
  NAND_GATE U5210 ( .I1(n4002), .I2(n4001), .O(n4003) );
  NAND_GATE U5211 ( .I1(n4004), .I2(n4003), .O(n4391) );
  NAND_GATE U5212 ( .I1(n4392), .I2(n4391), .O(n4006) );
  NAND3_GATE U5213 ( .I1(n4388), .I2(n4387), .I3(n4006), .O(n4381) );
  NAND_GATE U5214 ( .I1(n4021), .I2(n4381), .O(n4376) );
  INV_GATE U5215 ( .I1(n4007), .O(n4008) );
  NAND_GATE U5216 ( .I1(n4008), .I2(n4011), .O(n4020) );
  NAND_GATE U5217 ( .I1(n4010), .I2(n4014), .O(n4018) );
  NAND_GATE U5218 ( .I1(n4012), .I2(n4011), .O(n4013) );
  NAND_GATE U5219 ( .I1(n4014), .I2(n4013), .O(n4015) );
  NAND_GATE U5220 ( .I1(n4016), .I2(n4015), .O(n4017) );
  NAND_GATE U5221 ( .I1(n4018), .I2(n4017), .O(n4019) );
  NAND_GATE U5222 ( .I1(n4020), .I2(n4019), .O(n4380) );
  NAND_GATE U5223 ( .I1(n4381), .I2(n4380), .O(n4022) );
  NAND3_GATE U5224 ( .I1(n4376), .I2(n4375), .I3(n4022), .O(n4369) );
  NAND_GATE U5225 ( .I1(n4037), .I2(n4369), .O(n4363) );
  INV_GATE U5226 ( .I1(n4023), .O(n4024) );
  NAND_GATE U5227 ( .I1(n4024), .I2(n4027), .O(n4036) );
  NAND_GATE U5228 ( .I1(n4026), .I2(n4030), .O(n4034) );
  NAND_GATE U5229 ( .I1(n4028), .I2(n4027), .O(n4029) );
  NAND_GATE U5230 ( .I1(n4030), .I2(n4029), .O(n4031) );
  NAND_GATE U5231 ( .I1(n4032), .I2(n4031), .O(n4033) );
  NAND_GATE U5232 ( .I1(n4034), .I2(n4033), .O(n4035) );
  NAND_GATE U5233 ( .I1(n4036), .I2(n4035), .O(n4367) );
  NAND_GATE U5234 ( .I1(n4037), .I2(n4367), .O(n4362) );
  NAND_GATE U5235 ( .I1(n4369), .I2(n4367), .O(n4038) );
  NAND3_GATE U5236 ( .I1(n4363), .I2(n4362), .I3(n4038), .O(n4356) );
  NAND_GATE U5237 ( .I1(n4053), .I2(n4356), .O(n4350) );
  INV_GATE U5238 ( .I1(n4039), .O(n4040) );
  NAND_GATE U5239 ( .I1(n4040), .I2(n4043), .O(n4052) );
  NAND_GATE U5240 ( .I1(n4042), .I2(n4046), .O(n4050) );
  NAND_GATE U5241 ( .I1(n4044), .I2(n4043), .O(n4045) );
  NAND_GATE U5242 ( .I1(n4046), .I2(n4045), .O(n4047) );
  NAND_GATE U5243 ( .I1(n4048), .I2(n4047), .O(n4049) );
  NAND_GATE U5244 ( .I1(n4050), .I2(n4049), .O(n4051) );
  NAND_GATE U5245 ( .I1(n4052), .I2(n4051), .O(n4354) );
  NAND_GATE U5246 ( .I1(n4053), .I2(n4354), .O(n4349) );
  NAND_GATE U5247 ( .I1(n4356), .I2(n4354), .O(n4054) );
  NAND3_GATE U5248 ( .I1(n4350), .I2(n4349), .I3(n4054), .O(n4343) );
  NAND_GATE U5249 ( .I1(n4069), .I2(n4343), .O(n4337) );
  INV_GATE U5250 ( .I1(n4055), .O(n4056) );
  NAND_GATE U5251 ( .I1(n4056), .I2(n4059), .O(n4068) );
  NAND_GATE U5252 ( .I1(n4058), .I2(n4062), .O(n4066) );
  NAND_GATE U5253 ( .I1(n4060), .I2(n4059), .O(n4061) );
  NAND_GATE U5254 ( .I1(n4062), .I2(n4061), .O(n4063) );
  NAND_GATE U5255 ( .I1(n4064), .I2(n4063), .O(n4065) );
  NAND_GATE U5256 ( .I1(n4066), .I2(n4065), .O(n4067) );
  NAND_GATE U5257 ( .I1(n4068), .I2(n4067), .O(n4341) );
  NAND_GATE U5258 ( .I1(n4069), .I2(n4341), .O(n4336) );
  NAND_GATE U5259 ( .I1(n4343), .I2(n4341), .O(n4070) );
  NAND3_GATE U5260 ( .I1(n4337), .I2(n4336), .I3(n4070), .O(n4330) );
  NAND_GATE U5261 ( .I1(n4085), .I2(n4330), .O(n4326) );
  INV_GATE U5262 ( .I1(n4071), .O(n4072) );
  NAND_GATE U5263 ( .I1(n4072), .I2(n4075), .O(n4084) );
  NAND_GATE U5264 ( .I1(n4074), .I2(n4078), .O(n4082) );
  NAND_GATE U5265 ( .I1(n4076), .I2(n4075), .O(n4077) );
  NAND_GATE U5266 ( .I1(n4078), .I2(n4077), .O(n4079) );
  NAND_GATE U5267 ( .I1(n4080), .I2(n4079), .O(n4081) );
  NAND_GATE U5268 ( .I1(n4082), .I2(n4081), .O(n4083) );
  NAND_GATE U5269 ( .I1(n4084), .I2(n4083), .O(n4329) );
  NAND_GATE U5270 ( .I1(n4085), .I2(n4329), .O(n4325) );
  NAND_GATE U5271 ( .I1(n4330), .I2(n4329), .O(n4086) );
  NAND3_GATE U5272 ( .I1(n4326), .I2(n4325), .I3(n4086), .O(n4677) );
  NAND_GATE U5273 ( .I1(n4101), .I2(n4677), .O(n4671) );
  INV_GATE U5274 ( .I1(n4087), .O(n4088) );
  NAND_GATE U5275 ( .I1(n4088), .I2(n4091), .O(n4100) );
  NAND_GATE U5276 ( .I1(n4090), .I2(n4094), .O(n4098) );
  NAND_GATE U5277 ( .I1(n4092), .I2(n4091), .O(n4093) );
  NAND_GATE U5278 ( .I1(n4094), .I2(n4093), .O(n4095) );
  NAND_GATE U5279 ( .I1(n4096), .I2(n4095), .O(n4097) );
  NAND_GATE U5280 ( .I1(n4098), .I2(n4097), .O(n4099) );
  NAND_GATE U5281 ( .I1(n4100), .I2(n4099), .O(n4675) );
  NAND_GATE U5282 ( .I1(n4101), .I2(n4675), .O(n4670) );
  NAND_GATE U5283 ( .I1(n4677), .I2(n4675), .O(n4102) );
  NAND3_GATE U5284 ( .I1(n4671), .I2(n4670), .I3(n4102), .O(n4319) );
  NAND_GATE U5285 ( .I1(n4118), .I2(n4319), .O(n4315) );
  INV_GATE U5286 ( .I1(n4103), .O(n4104) );
  NAND_GATE U5287 ( .I1(n4104), .I2(n4108), .O(n4117) );
  INV_GATE U5288 ( .I1(n4108), .O(n4105) );
  NAND_GATE U5289 ( .I1(n4106), .I2(n4105), .O(n4111) );
  NAND_GATE U5290 ( .I1(n4107), .I2(n4111), .O(n4115) );
  NAND_GATE U5291 ( .I1(n4109), .I2(n4108), .O(n4110) );
  NAND_GATE U5292 ( .I1(n4111), .I2(n4110), .O(n4112) );
  NAND_GATE U5293 ( .I1(n4113), .I2(n4112), .O(n4114) );
  NAND_GATE U5294 ( .I1(n4115), .I2(n4114), .O(n4116) );
  NAND_GATE U5295 ( .I1(n4117), .I2(n4116), .O(n4318) );
  NAND_GATE U5296 ( .I1(n4118), .I2(n4318), .O(n4314) );
  NAND_GATE U5297 ( .I1(n4319), .I2(n4318), .O(n4119) );
  NAND3_GATE U5298 ( .I1(n4315), .I2(n4314), .I3(n4119), .O(n4308) );
  NAND_GATE U5299 ( .I1(n4120), .I2(n4308), .O(n4303) );
  NAND_GATE U5300 ( .I1(n4307), .I2(n4308), .O(n4121) );
  NAND3_GATE U5301 ( .I1(n4304), .I2(n4303), .I3(n4121), .O(n4297) );
  NAND_GATE U5302 ( .I1(n4137), .I2(n4297), .O(n4293) );
  INV_GATE U5303 ( .I1(n4122), .O(n4123) );
  NAND_GATE U5304 ( .I1(n4123), .I2(n4127), .O(n4136) );
  INV_GATE U5305 ( .I1(n4127), .O(n4124) );
  NAND_GATE U5306 ( .I1(n4125), .I2(n4124), .O(n4130) );
  NAND_GATE U5307 ( .I1(n4126), .I2(n4130), .O(n4134) );
  NAND_GATE U5308 ( .I1(n4128), .I2(n4127), .O(n4129) );
  NAND_GATE U5309 ( .I1(n4130), .I2(n4129), .O(n4131) );
  NAND_GATE U5310 ( .I1(n4132), .I2(n4131), .O(n4133) );
  NAND_GATE U5311 ( .I1(n4134), .I2(n4133), .O(n4135) );
  NAND_GATE U5312 ( .I1(n4136), .I2(n4135), .O(n4296) );
  NAND_GATE U5313 ( .I1(n4137), .I2(n4296), .O(n4292) );
  NAND_GATE U5314 ( .I1(n4297), .I2(n4296), .O(n4138) );
  NAND3_GATE U5315 ( .I1(n4293), .I2(n4292), .I3(n4138), .O(n4286) );
  NAND_GATE U5316 ( .I1(n4153), .I2(n4286), .O(n4282) );
  OR_GATE U5317 ( .I1(n4140), .I2(n4139), .O(n4152) );
  NAND_GATE U5318 ( .I1(n4141), .I2(n4140), .O(n4146) );
  NAND_GATE U5319 ( .I1(n4142), .I2(n4146), .O(n4150) );
  NAND_GATE U5320 ( .I1(n4144), .I2(n4143), .O(n4145) );
  NAND_GATE U5321 ( .I1(n4146), .I2(n4145), .O(n4147) );
  NAND_GATE U5322 ( .I1(n4148), .I2(n4147), .O(n4149) );
  NAND_GATE U5323 ( .I1(n4150), .I2(n4149), .O(n4151) );
  NAND_GATE U5324 ( .I1(n4152), .I2(n4151), .O(n4285) );
  NAND_GATE U5325 ( .I1(n4153), .I2(n4285), .O(n4281) );
  NAND_GATE U5326 ( .I1(n4286), .I2(n4285), .O(n4154) );
  NAND3_GATE U5327 ( .I1(n4282), .I2(n4281), .I3(n4154), .O(n4275) );
  NAND_GATE U5328 ( .I1(n4169), .I2(n4275), .O(n4271) );
  INV_GATE U5329 ( .I1(n4155), .O(n4156) );
  NAND_GATE U5330 ( .I1(n4156), .I2(n4159), .O(n4168) );
  NAND_GATE U5331 ( .I1(n4158), .I2(n4162), .O(n4166) );
  NAND_GATE U5332 ( .I1(n4160), .I2(n4159), .O(n4161) );
  NAND_GATE U5333 ( .I1(n4162), .I2(n4161), .O(n4163) );
  NAND_GATE U5334 ( .I1(n4164), .I2(n4163), .O(n4165) );
  NAND_GATE U5335 ( .I1(n4166), .I2(n4165), .O(n4167) );
  NAND_GATE U5336 ( .I1(n4168), .I2(n4167), .O(n4274) );
  NAND_GATE U5337 ( .I1(n4169), .I2(n4274), .O(n4270) );
  NAND_GATE U5338 ( .I1(n4275), .I2(n4274), .O(n4170) );
  NAND3_GATE U5339 ( .I1(n4271), .I2(n4270), .I3(n4170), .O(n4264) );
  NAND_GATE U5340 ( .I1(n4185), .I2(n4264), .O(n4260) );
  INV_GATE U5341 ( .I1(n4171), .O(n4172) );
  NAND_GATE U5342 ( .I1(n4172), .I2(n4175), .O(n4184) );
  NAND_GATE U5343 ( .I1(n4174), .I2(n4178), .O(n4182) );
  NAND_GATE U5344 ( .I1(n4176), .I2(n4175), .O(n4177) );
  NAND_GATE U5345 ( .I1(n4178), .I2(n4177), .O(n4179) );
  NAND_GATE U5346 ( .I1(n4180), .I2(n4179), .O(n4181) );
  NAND_GATE U5347 ( .I1(n4182), .I2(n4181), .O(n4183) );
  NAND_GATE U5348 ( .I1(n4184), .I2(n4183), .O(n4263) );
  NAND_GATE U5349 ( .I1(n4185), .I2(n4263), .O(n4259) );
  NAND_GATE U5350 ( .I1(n4264), .I2(n4263), .O(n4186) );
  NAND3_GATE U5351 ( .I1(n4260), .I2(n4259), .I3(n4186), .O(n4253) );
  NAND_GATE U5352 ( .I1(n4201), .I2(n4253), .O(n4249) );
  INV_GATE U5353 ( .I1(n4187), .O(n4188) );
  NAND_GATE U5354 ( .I1(n4188), .I2(n4191), .O(n4200) );
  NAND_GATE U5355 ( .I1(n4190), .I2(n4194), .O(n4198) );
  NAND_GATE U5356 ( .I1(n4192), .I2(n4191), .O(n4193) );
  NAND_GATE U5357 ( .I1(n4194), .I2(n4193), .O(n4195) );
  NAND_GATE U5358 ( .I1(n4196), .I2(n4195), .O(n4197) );
  NAND_GATE U5359 ( .I1(n4198), .I2(n4197), .O(n4199) );
  NAND_GATE U5360 ( .I1(n4200), .I2(n4199), .O(n4252) );
  NAND_GATE U5361 ( .I1(n4201), .I2(n4252), .O(n4248) );
  NAND_GATE U5362 ( .I1(n4253), .I2(n4252), .O(n4202) );
  NAND3_GATE U5363 ( .I1(n4249), .I2(n4248), .I3(n4202), .O(n4242) );
  NAND_GATE U5364 ( .I1(n4217), .I2(n4242), .O(n4238) );
  INV_GATE U5365 ( .I1(n4203), .O(n4204) );
  NAND_GATE U5366 ( .I1(n4204), .I2(n4207), .O(n4216) );
  NAND_GATE U5367 ( .I1(n4206), .I2(n4210), .O(n4214) );
  NAND_GATE U5368 ( .I1(n4208), .I2(n4207), .O(n4209) );
  NAND_GATE U5369 ( .I1(n4210), .I2(n4209), .O(n4211) );
  NAND_GATE U5370 ( .I1(n4212), .I2(n4211), .O(n4213) );
  NAND_GATE U5371 ( .I1(n4214), .I2(n4213), .O(n4215) );
  NAND_GATE U5372 ( .I1(n4216), .I2(n4215), .O(n4241) );
  NAND_GATE U5373 ( .I1(n4217), .I2(n4241), .O(n4237) );
  NAND_GATE U5374 ( .I1(n4242), .I2(n4241), .O(n4218) );
  NAND3_GATE U5375 ( .I1(n4238), .I2(n4237), .I3(n4218), .O(n15315) );
  INV_GATE U5376 ( .I1(n15315), .O(n4233) );
  INV_GATE U5377 ( .I1(n4219), .O(n4220) );
  NAND_GATE U5378 ( .I1(n4220), .I2(n4223), .O(n4232) );
  NAND_GATE U5379 ( .I1(n4222), .I2(n4226), .O(n4230) );
  NAND_GATE U5380 ( .I1(n4224), .I2(n4223), .O(n4225) );
  NAND_GATE U5381 ( .I1(n4226), .I2(n4225), .O(n4227) );
  NAND_GATE U5382 ( .I1(n4228), .I2(n4227), .O(n4229) );
  NAND_GATE U5383 ( .I1(n4230), .I2(n4229), .O(n4231) );
  NAND_GATE U5384 ( .I1(n4232), .I2(n4231), .O(n15314) );
  NAND_GATE U5385 ( .I1(n4233), .I2(n15314), .O(n4236) );
  INV_GATE U5386 ( .I1(n15314), .O(n4234) );
  NAND_GATE U5387 ( .I1(n15315), .I2(n4234), .O(n4235) );
  NAND_GATE U5388 ( .I1(n4236), .I2(n4235), .O(\A1[54] ) );
  OR_GATE U5389 ( .I1(n4237), .I2(n4242), .O(n4240) );
  OR_GATE U5390 ( .I1(n4241), .I2(n4238), .O(n4239) );
  AND_GATE U5391 ( .I1(n4240), .I2(n4239), .O(n4247) );
  NAND_GATE U5392 ( .I1(n4242), .I2(n1130), .O(n4244) );
  NAND3_GATE U5393 ( .I1(n4245), .I2(n4244), .I3(n4243), .O(n4246) );
  OR_GATE U5394 ( .I1(n4248), .I2(n4253), .O(n4251) );
  OR_GATE U5395 ( .I1(n4252), .I2(n4249), .O(n4250) );
  AND_GATE U5396 ( .I1(n4251), .I2(n4250), .O(n4258) );
  NAND_GATE U5397 ( .I1(n4253), .I2(n1127), .O(n4255) );
  NAND3_GATE U5398 ( .I1(n4256), .I2(n4255), .I3(n4254), .O(n4257) );
  NAND_GATE U5399 ( .I1(n4258), .I2(n4257), .O(n5130) );
  INV_GATE U5400 ( .I1(n5130), .O(n5133) );
  NAND_GATE U5401 ( .I1(B[23]), .I2(A[31]), .O(n5137) );
  INV_GATE U5402 ( .I1(n5137), .O(n5131) );
  NAND_GATE U5403 ( .I1(n5133), .I2(n5131), .O(n5128) );
  OR_GATE U5404 ( .I1(n4259), .I2(n4264), .O(n4262) );
  OR_GATE U5405 ( .I1(n4263), .I2(n4260), .O(n4261) );
  AND_GATE U5406 ( .I1(n4262), .I2(n4261), .O(n4269) );
  NAND_GATE U5407 ( .I1(n4264), .I2(n1123), .O(n4266) );
  NAND3_GATE U5408 ( .I1(n4267), .I2(n4266), .I3(n4265), .O(n4268) );
  NAND_GATE U5409 ( .I1(n4269), .I2(n4268), .O(n5114) );
  INV_GATE U5410 ( .I1(n5114), .O(n5117) );
  NAND_GATE U5411 ( .I1(B[23]), .I2(A[30]), .O(n5121) );
  INV_GATE U5412 ( .I1(n5121), .O(n5115) );
  NAND_GATE U5413 ( .I1(n5117), .I2(n5115), .O(n5112) );
  OR_GATE U5414 ( .I1(n4270), .I2(n4275), .O(n4273) );
  OR_GATE U5415 ( .I1(n4274), .I2(n4271), .O(n4272) );
  AND_GATE U5416 ( .I1(n4273), .I2(n4272), .O(n4280) );
  NAND_GATE U5417 ( .I1(n1111), .I2(n4274), .O(n4278) );
  NAND3_GATE U5418 ( .I1(n4278), .I2(n4277), .I3(n4276), .O(n4279) );
  NAND_GATE U5419 ( .I1(n4280), .I2(n4279), .O(n5098) );
  INV_GATE U5420 ( .I1(n5098), .O(n5101) );
  NAND_GATE U5421 ( .I1(B[23]), .I2(A[29]), .O(n5105) );
  INV_GATE U5422 ( .I1(n5105), .O(n5099) );
  NAND_GATE U5423 ( .I1(n5101), .I2(n5099), .O(n5095) );
  OR_GATE U5424 ( .I1(n4281), .I2(n4286), .O(n4284) );
  OR_GATE U5425 ( .I1(n4285), .I2(n4282), .O(n4283) );
  AND_GATE U5426 ( .I1(n4284), .I2(n4283), .O(n4291) );
  NAND_GATE U5427 ( .I1(n1106), .I2(n4285), .O(n4289) );
  NAND3_GATE U5428 ( .I1(n4289), .I2(n4288), .I3(n4287), .O(n4290) );
  NAND_GATE U5429 ( .I1(n4291), .I2(n4290), .O(n5081) );
  INV_GATE U5430 ( .I1(n5081), .O(n5084) );
  NAND_GATE U5431 ( .I1(B[23]), .I2(A[28]), .O(n5088) );
  INV_GATE U5432 ( .I1(n5088), .O(n5082) );
  NAND_GATE U5433 ( .I1(n5084), .I2(n5082), .O(n5079) );
  OR_GATE U5434 ( .I1(n4292), .I2(n4297), .O(n4295) );
  OR_GATE U5435 ( .I1(n4296), .I2(n4293), .O(n4294) );
  AND_GATE U5436 ( .I1(n4295), .I2(n4294), .O(n4302) );
  NAND_GATE U5437 ( .I1(n1100), .I2(n4296), .O(n4300) );
  NAND3_GATE U5438 ( .I1(n4300), .I2(n4299), .I3(n4298), .O(n4301) );
  NAND_GATE U5439 ( .I1(n4302), .I2(n4301), .O(n5065) );
  INV_GATE U5440 ( .I1(n5065), .O(n5068) );
  NAND_GATE U5441 ( .I1(B[23]), .I2(A[27]), .O(n5072) );
  INV_GATE U5442 ( .I1(n5072), .O(n5066) );
  NAND_GATE U5443 ( .I1(n5068), .I2(n5066), .O(n5062) );
  OR_GATE U5444 ( .I1(n4303), .I2(n4307), .O(n4306) );
  OR_GATE U5445 ( .I1(n4308), .I2(n4304), .O(n4305) );
  AND_GATE U5446 ( .I1(n4306), .I2(n4305), .O(n4313) );
  NAND_GATE U5447 ( .I1(n4307), .I2(n1092), .O(n4311) );
  NAND3_GATE U5448 ( .I1(n4311), .I2(n4310), .I3(n4309), .O(n4312) );
  NAND_GATE U5449 ( .I1(n4313), .I2(n4312), .O(n5048) );
  INV_GATE U5450 ( .I1(n5048), .O(n5051) );
  NAND_GATE U5451 ( .I1(B[23]), .I2(A[26]), .O(n5055) );
  INV_GATE U5452 ( .I1(n5055), .O(n5049) );
  NAND_GATE U5453 ( .I1(n5051), .I2(n5049), .O(n5045) );
  OR_GATE U5454 ( .I1(n4314), .I2(n4319), .O(n4317) );
  OR_GATE U5455 ( .I1(n4318), .I2(n4315), .O(n4316) );
  AND_GATE U5456 ( .I1(n4317), .I2(n4316), .O(n4324) );
  NAND_GATE U5457 ( .I1(n1086), .I2(n4318), .O(n4322) );
  NAND3_GATE U5458 ( .I1(n4322), .I2(n4321), .I3(n4320), .O(n4323) );
  NAND_GATE U5459 ( .I1(n4324), .I2(n4323), .O(n5031) );
  INV_GATE U5460 ( .I1(n5031), .O(n5034) );
  NAND_GATE U5461 ( .I1(B[23]), .I2(A[25]), .O(n5038) );
  INV_GATE U5462 ( .I1(n5038), .O(n5032) );
  NAND_GATE U5463 ( .I1(n5034), .I2(n5032), .O(n5029) );
  NAND_GATE U5464 ( .I1(B[23]), .I2(A[24]), .O(n5022) );
  INV_GATE U5465 ( .I1(n5022), .O(n5016) );
  OR_GATE U5466 ( .I1(n4325), .I2(n4330), .O(n4328) );
  OR_GATE U5467 ( .I1(n4329), .I2(n4326), .O(n4327) );
  AND_GATE U5468 ( .I1(n4328), .I2(n4327), .O(n4335) );
  NAND_GATE U5469 ( .I1(n4330), .I2(n1060), .O(n4332) );
  NAND3_GATE U5470 ( .I1(n4333), .I2(n4332), .I3(n4331), .O(n4334) );
  NAND_GATE U5471 ( .I1(n4335), .I2(n4334), .O(n4999) );
  INV_GATE U5472 ( .I1(n4999), .O(n5002) );
  NAND_GATE U5473 ( .I1(B[23]), .I2(A[23]), .O(n5006) );
  INV_GATE U5474 ( .I1(n5006), .O(n5000) );
  NAND_GATE U5475 ( .I1(n5002), .I2(n5000), .O(n4997) );
  OR_GATE U5476 ( .I1(n4336), .I2(n4343), .O(n4339) );
  OR_GATE U5477 ( .I1(n4341), .I2(n4337), .O(n4338) );
  AND_GATE U5478 ( .I1(n4339), .I2(n4338), .O(n4348) );
  INV_GATE U5479 ( .I1(n4343), .O(n4340) );
  NAND_GATE U5480 ( .I1(n4340), .I2(n4341), .O(n4346) );
  INV_GATE U5481 ( .I1(n4341), .O(n4342) );
  NAND_GATE U5482 ( .I1(n4343), .I2(n4342), .O(n4345) );
  NAND3_GATE U5483 ( .I1(n4346), .I2(n4345), .I3(n4344), .O(n4347) );
  NAND_GATE U5484 ( .I1(n4348), .I2(n4347), .O(n4703) );
  INV_GATE U5485 ( .I1(n4703), .O(n4706) );
  NAND_GATE U5486 ( .I1(B[23]), .I2(A[22]), .O(n4710) );
  INV_GATE U5487 ( .I1(n4710), .O(n4704) );
  NAND_GATE U5488 ( .I1(n4706), .I2(n4704), .O(n4701) );
  OR_GATE U5489 ( .I1(n4349), .I2(n4356), .O(n4352) );
  OR_GATE U5490 ( .I1(n4354), .I2(n4350), .O(n4351) );
  AND_GATE U5491 ( .I1(n4352), .I2(n4351), .O(n4361) );
  INV_GATE U5492 ( .I1(n4356), .O(n4353) );
  NAND_GATE U5493 ( .I1(n4353), .I2(n4354), .O(n4359) );
  INV_GATE U5494 ( .I1(n4354), .O(n4355) );
  NAND_GATE U5495 ( .I1(n4356), .I2(n4355), .O(n4358) );
  NAND3_GATE U5496 ( .I1(n4359), .I2(n4358), .I3(n4357), .O(n4360) );
  NAND_GATE U5497 ( .I1(n4361), .I2(n4360), .O(n4981) );
  INV_GATE U5498 ( .I1(n4981), .O(n4984) );
  NAND_GATE U5499 ( .I1(B[23]), .I2(A[21]), .O(n4988) );
  INV_GATE U5500 ( .I1(n4988), .O(n4982) );
  NAND_GATE U5501 ( .I1(n4984), .I2(n4982), .O(n4979) );
  OR_GATE U5502 ( .I1(n4362), .I2(n4369), .O(n4365) );
  OR_GATE U5503 ( .I1(n4367), .I2(n4363), .O(n4364) );
  AND_GATE U5504 ( .I1(n4365), .I2(n4364), .O(n4374) );
  INV_GATE U5505 ( .I1(n4369), .O(n4366) );
  NAND_GATE U5506 ( .I1(n4366), .I2(n4367), .O(n4372) );
  INV_GATE U5507 ( .I1(n4367), .O(n4368) );
  NAND_GATE U5508 ( .I1(n4369), .I2(n4368), .O(n4371) );
  NAND3_GATE U5509 ( .I1(n4372), .I2(n4371), .I3(n4370), .O(n4373) );
  NAND_GATE U5510 ( .I1(n4374), .I2(n4373), .O(n4965) );
  INV_GATE U5511 ( .I1(n4965), .O(n4968) );
  NAND_GATE U5512 ( .I1(B[23]), .I2(A[20]), .O(n4972) );
  INV_GATE U5513 ( .I1(n4972), .O(n4966) );
  NAND_GATE U5514 ( .I1(n4968), .I2(n4966), .O(n4963) );
  OR_GATE U5515 ( .I1(n4375), .I2(n4381), .O(n4378) );
  OR_GATE U5516 ( .I1(n4380), .I2(n4376), .O(n4377) );
  AND_GATE U5517 ( .I1(n4378), .I2(n4377), .O(n4386) );
  INV_GATE U5518 ( .I1(n4381), .O(n4379) );
  NAND_GATE U5519 ( .I1(n4379), .I2(n4380), .O(n4384) );
  NAND_GATE U5520 ( .I1(n4381), .I2(n396), .O(n4383) );
  NAND3_GATE U5521 ( .I1(n4384), .I2(n4383), .I3(n4382), .O(n4385) );
  NAND_GATE U5522 ( .I1(n4386), .I2(n4385), .O(n4953) );
  INV_GATE U5523 ( .I1(n4953), .O(n4952) );
  NAND_GATE U5524 ( .I1(B[23]), .I2(A[19]), .O(n4956) );
  INV_GATE U5525 ( .I1(n4956), .O(n4950) );
  NAND_GATE U5526 ( .I1(n4952), .I2(n4950), .O(n4947) );
  OR_GATE U5527 ( .I1(n4387), .I2(n4392), .O(n4390) );
  OR_GATE U5528 ( .I1(n4391), .I2(n4388), .O(n4389) );
  NAND_GATE U5529 ( .I1(n397), .I2(n4391), .O(n4395) );
  NAND3_GATE U5530 ( .I1(n4395), .I2(n4394), .I3(n4393), .O(n4396) );
  NAND_GATE U5531 ( .I1(B[23]), .I2(A[18]), .O(n4941) );
  INV_GATE U5532 ( .I1(n4941), .O(n4935) );
  NAND_GATE U5533 ( .I1(n398), .I2(n4935), .O(n4932) );
  OR_GATE U5534 ( .I1(n4397), .I2(n4402), .O(n4400) );
  OR_GATE U5535 ( .I1(n4401), .I2(n4398), .O(n4399) );
  NAND_GATE U5536 ( .I1(n584), .I2(n4401), .O(n4405) );
  NAND3_GATE U5537 ( .I1(n4405), .I2(n4404), .I3(n4403), .O(n4406) );
  INV_GATE U5538 ( .I1(n4922), .O(n4921) );
  NAND_GATE U5539 ( .I1(B[23]), .I2(A[17]), .O(n4925) );
  INV_GATE U5540 ( .I1(n4925), .O(n4919) );
  NAND_GATE U5541 ( .I1(n4921), .I2(n4919), .O(n4916) );
  OR_GATE U5542 ( .I1(n4407), .I2(n4413), .O(n4410) );
  OR_GATE U5543 ( .I1(n4414), .I2(n4408), .O(n4409) );
  AND_GATE U5544 ( .I1(n4410), .I2(n4409), .O(n4420) );
  NAND_GATE U5545 ( .I1(n4411), .I2(n3971), .O(n4412) );
  NAND_GATE U5546 ( .I1(n4413), .I2(n4412), .O(n4417) );
  INV_GATE U5547 ( .I1(n4413), .O(n4415) );
  NAND_GATE U5548 ( .I1(n4415), .I2(n4414), .O(n4416) );
  NAND3_GATE U5549 ( .I1(n4418), .I2(n4417), .I3(n4416), .O(n4419) );
  NAND_GATE U5550 ( .I1(n4420), .I2(n4419), .O(n4907) );
  INV_GATE U5551 ( .I1(n4907), .O(n4905) );
  NAND_GATE U5552 ( .I1(B[23]), .I2(A[16]), .O(n4909) );
  INV_GATE U5553 ( .I1(n4909), .O(n4903) );
  NAND_GATE U5554 ( .I1(n4905), .I2(n4903), .O(n4901) );
  OR_GATE U5555 ( .I1(n4421), .I2(n4425), .O(n4434) );
  NAND_GATE U5556 ( .I1(n4423), .I2(n4422), .O(n4424) );
  NAND_GATE U5557 ( .I1(n4425), .I2(n4424), .O(n4428) );
  INV_GATE U5558 ( .I1(n4425), .O(n4426) );
  NAND_GATE U5559 ( .I1(n4426), .I2(n4431), .O(n4427) );
  NAND3_GATE U5560 ( .I1(n4429), .I2(n4428), .I3(n4427), .O(n4433) );
  OR_GATE U5561 ( .I1(n4431), .I2(n4430), .O(n4432) );
  NAND3_GATE U5562 ( .I1(n4434), .I2(n4433), .I3(n4432), .O(n4890) );
  NAND_GATE U5563 ( .I1(B[23]), .I2(A[15]), .O(n4894) );
  INV_GATE U5564 ( .I1(n4894), .O(n4887) );
  NAND_GATE U5565 ( .I1(n17), .I2(n4887), .O(n4884) );
  OR_GATE U5566 ( .I1(n4435), .I2(n4440), .O(n4438) );
  OR_GATE U5567 ( .I1(n4439), .I2(n4436), .O(n4437) );
  AND_GATE U5568 ( .I1(n4438), .I2(n4437), .O(n4445) );
  NAND_GATE U5569 ( .I1(n4440), .I2(n757), .O(n4442) );
  NAND3_GATE U5570 ( .I1(n4443), .I2(n4442), .I3(n4441), .O(n4444) );
  NAND_GATE U5571 ( .I1(n4445), .I2(n4444), .O(n4878) );
  INV_GATE U5572 ( .I1(n4878), .O(n4876) );
  NAND_GATE U5573 ( .I1(B[23]), .I2(A[14]), .O(n5316) );
  INV_GATE U5574 ( .I1(n5316), .O(n4874) );
  NAND_GATE U5575 ( .I1(n4876), .I2(n4874), .O(n4873) );
  NAND_GATE U5576 ( .I1(B[23]), .I2(A[13]), .O(n5326) );
  INV_GATE U5577 ( .I1(n5326), .O(n4720) );
  NAND_GATE U5578 ( .I1(n4447), .I2(n4446), .O(n4451) );
  NAND_GATE U5579 ( .I1(n4451), .I2(n4450), .O(n4452) );
  NAND_GATE U5580 ( .I1(n4459), .I2(n4452), .O(n4454) );
  OR_GATE U5581 ( .I1(n4452), .I2(n4459), .O(n4453) );
  NAND3_GATE U5582 ( .I1(n4455), .I2(n4454), .I3(n4453), .O(n4462) );
  OR_GATE U5583 ( .I1(n4457), .I2(n4456), .O(n4461) );
  OR_GATE U5584 ( .I1(n4459), .I2(n4458), .O(n4460) );
  NAND3_GATE U5585 ( .I1(n4462), .I2(n4461), .I3(n4460), .O(n4717) );
  INV_GATE U5586 ( .I1(n4717), .O(n4718) );
  NAND_GATE U5587 ( .I1(n4720), .I2(n4718), .O(n4649) );
  NAND_GATE U5588 ( .I1(n712), .I2(n4463), .O(n4464) );
  NAND_GATE U5589 ( .I1(n4465), .I2(n4464), .O(n4474) );
  NAND_GATE U5590 ( .I1(n4467), .I2(n4473), .O(n4466) );
  NAND_GATE U5591 ( .I1(n4606), .I2(n4466), .O(n4601) );
  NAND_GATE U5592 ( .I1(B[23]), .I2(A[10]), .O(n5375) );
  NAND4_GATE U5593 ( .I1(n4469), .I2(n4468), .I3(n4473), .I4(n4467), .O(n4599)
         );
  NAND4_GATE U5594 ( .I1(n4600), .I2(n4601), .I3(n5375), .I4(n4599), .O(n4598)
         );
  INV_GATE U5595 ( .I1(n4470), .O(n4609) );
  NAND_GATE U5596 ( .I1(n4472), .I2(n4471), .O(n4473) );
  NAND_GATE U5597 ( .I1(n4474), .I2(n4473), .O(n4475) );
  AND_GATE U5598 ( .I1(n4476), .I2(n4475), .O(n4477) );
  NAND_GATE U5599 ( .I1(n4609), .I2(n4477), .O(n4481) );
  INV_GATE U5600 ( .I1(n4606), .O(n4479) );
  AND_GATE U5601 ( .I1(n4608), .I2(n4607), .O(n4478) );
  NAND3_GATE U5602 ( .I1(n4479), .I2(n4478), .I3(n4473), .O(n4480) );
  NAND_GATE U5603 ( .I1(n4481), .I2(n4480), .O(n4602) );
  NAND_GATE U5604 ( .I1(n5375), .I2(n4602), .O(n4597) );
  NAND_GATE U5605 ( .I1(n254), .I2(n4483), .O(n4798) );
  NAND3_GATE U5606 ( .I1(n4482), .I2(n4799), .I3(n549), .O(n4805) );
  NAND3_GATE U5607 ( .I1(n4798), .I2(n4805), .I3(n4799), .O(n4812) );
  NAND_GATE U5608 ( .I1(n4484), .I2(n4798), .O(n4800) );
  NAND_GATE U5609 ( .I1(n4801), .I2(n4800), .O(n4811) );
  NAND_GATE U5610 ( .I1(B[23]), .I2(A[6]), .O(n5399) );
  INV_GATE U5611 ( .I1(n5399), .O(n4790) );
  INV_GATE U5612 ( .I1(n4486), .O(n4500) );
  NAND3_GATE U5613 ( .I1(n4494), .I2(n4498), .I3(n4500), .O(n4551) );
  NAND_GATE U5614 ( .I1(n4498), .I2(n4494), .O(n4485) );
  NAND_GATE U5615 ( .I1(n4486), .I2(n4485), .O(n4550) );
  AND3_GATE U5616 ( .I1(n4551), .I2(n4552), .I3(n4550), .O(n4503) );
  INV_GATE U5617 ( .I1(n4487), .O(n4489) );
  AND_GATE U5618 ( .I1(n4489), .I2(n4488), .O(n4497) );
  NAND_GATE U5619 ( .I1(n4491), .I2(n4490), .O(n4495) );
  NAND_GATE U5620 ( .I1(n4493), .I2(n4492), .O(n4494) );
  NAND_GATE U5621 ( .I1(n4495), .I2(n4494), .O(n4496) );
  NAND_GATE U5622 ( .I1(n4497), .I2(n4496), .O(n4502) );
  NAND4_GATE U5623 ( .I1(n4500), .I2(n4494), .I3(n4499), .I4(n4498), .O(n4501)
         );
  NAND_GATE U5624 ( .I1(n4502), .I2(n4501), .O(n4549) );
  NAND_GATE U5625 ( .I1(n4790), .I2(n854), .O(n4556) );
  NAND_GATE U5626 ( .I1(n4505), .I2(n820), .O(n4504) );
  NAND_GATE U5627 ( .I1(n4725), .I2(n4504), .O(n4733) );
  NAND_GATE U5628 ( .I1(n4724), .I2(n4725), .O(n4735) );
  INV_GATE U5629 ( .I1(n4735), .O(n4506) );
  NAND3_GATE U5630 ( .I1(n4505), .I2(n4724), .I3(n820), .O(n4737) );
  NAND_GATE U5631 ( .I1(n4506), .I2(n4737), .O(n4722) );
  NAND3_GATE U5632 ( .I1(n4508), .I2(n4507), .I3(n4519), .O(n4509) );
  NAND_GATE U5633 ( .I1(n4510), .I2(n4509), .O(n4517) );
  NAND_GATE U5634 ( .I1(n4512), .I2(n4511), .O(n4516) );
  NAND3_GATE U5635 ( .I1(n4514), .I2(n4519), .I3(n4513), .O(n4515) );
  NAND3_GATE U5636 ( .I1(n4517), .I2(n4516), .I3(n4515), .O(n4521) );
  OR_GATE U5637 ( .I1(n4519), .I2(n4518), .O(n4520) );
  NAND_GATE U5638 ( .I1(n4521), .I2(n4520), .O(n4766) );
  NAND_GATE U5639 ( .I1(B[23]), .I2(A[2]), .O(n4755) );
  INV_GATE U5640 ( .I1(n4755), .O(n4741) );
  NAND_GATE U5641 ( .I1(n1391), .I2(A[1]), .O(n4522) );
  NAND_GATE U5642 ( .I1(n14784), .I2(n4522), .O(n4523) );
  NAND_GATE U5643 ( .I1(B[24]), .I2(n4523), .O(n4738) );
  NAND_GATE U5644 ( .I1(n1390), .I2(A[0]), .O(n4524) );
  NAND_GATE U5645 ( .I1(n14781), .I2(n4524), .O(n4525) );
  NAND_GATE U5646 ( .I1(B[25]), .I2(n4525), .O(n4739) );
  NAND_GATE U5647 ( .I1(n4738), .I2(n4739), .O(n4753) );
  NAND_GATE U5648 ( .I1(n4741), .I2(n4753), .O(n4742) );
  NAND3_GATE U5649 ( .I1(B[23]), .I2(B[24]), .I3(n1196), .O(n4752) );
  INV_GATE U5650 ( .I1(n4752), .O(n4754) );
  NAND_GATE U5651 ( .I1(n4755), .I2(n199), .O(n4526) );
  NAND_GATE U5652 ( .I1(n4754), .I2(n4526), .O(n4527) );
  NAND_GATE U5653 ( .I1(n4742), .I2(n4527), .O(n4767) );
  NAND_GATE U5654 ( .I1(n4766), .I2(n4767), .O(n4529) );
  NAND_GATE U5655 ( .I1(B[23]), .I2(A[3]), .O(n4771) );
  INV_GATE U5656 ( .I1(n4771), .O(n4761) );
  NAND_GATE U5657 ( .I1(n4766), .I2(n4761), .O(n4528) );
  NAND_GATE U5658 ( .I1(n4767), .I2(n4761), .O(n4762) );
  NAND3_GATE U5659 ( .I1(n4529), .I2(n4528), .I3(n4762), .O(n4782) );
  NAND_GATE U5660 ( .I1(B[23]), .I2(A[4]), .O(n5462) );
  NAND_GATE U5661 ( .I1(n4533), .I2(n4534), .O(n4530) );
  NAND_GATE U5662 ( .I1(n4531), .I2(n4530), .O(n4539) );
  OR_GATE U5663 ( .I1(n4539), .I2(n4532), .O(n4537) );
  INV_GATE U5664 ( .I1(n4538), .O(n4540) );
  NAND4_GATE U5665 ( .I1(n4535), .I2(n4534), .I3(n4533), .I4(n4540), .O(n4536)
         );
  AND_GATE U5666 ( .I1(n4537), .I2(n4536), .O(n4777) );
  NAND_GATE U5667 ( .I1(n4540), .I2(n4539), .O(n4542) );
  NAND3_GATE U5668 ( .I1(n4543), .I2(n4542), .I3(n4541), .O(n4778) );
  NAND_GATE U5669 ( .I1(n4777), .I2(n4778), .O(n5452) );
  NAND_GATE U5670 ( .I1(n5462), .I2(n5452), .O(n4544) );
  NAND_GATE U5671 ( .I1(n4782), .I2(n4544), .O(n4546) );
  INV_GATE U5672 ( .I1(n5462), .O(n5455) );
  NAND_GATE U5673 ( .I1(n5455), .I2(n1332), .O(n4545) );
  NAND_GATE U5674 ( .I1(n4546), .I2(n4545), .O(n4727) );
  NAND3_GATE U5675 ( .I1(n4729), .I2(n4722), .I3(n4727), .O(n4548) );
  NAND_GATE U5676 ( .I1(B[23]), .I2(A[5]), .O(n4730) );
  INV_GATE U5677 ( .I1(n4730), .O(n4723) );
  NAND3_GATE U5678 ( .I1(n4729), .I2(n4722), .I3(n4723), .O(n4547) );
  NAND_GATE U5679 ( .I1(n4723), .I2(n4727), .O(n4736) );
  NAND3_GATE U5680 ( .I1(n4548), .I2(n4547), .I3(n4736), .O(n4791) );
  NAND_GATE U5681 ( .I1(n5399), .I2(n4549), .O(n4554) );
  NAND4_GATE U5682 ( .I1(n4552), .I2(n5399), .I3(n4551), .I4(n4550), .O(n4553)
         );
  NAND3_GATE U5683 ( .I1(n4791), .I2(n4554), .I3(n4553), .O(n4555) );
  NAND_GATE U5684 ( .I1(n4556), .I2(n4555), .O(n4814) );
  NAND3_GATE U5685 ( .I1(n4812), .I2(n4811), .I3(n4814), .O(n4558) );
  NAND_GATE U5686 ( .I1(B[23]), .I2(A[7]), .O(n4817) );
  INV_GATE U5687 ( .I1(n4817), .O(n4807) );
  NAND3_GATE U5688 ( .I1(n4807), .I2(n4812), .I3(n4811), .O(n4557) );
  NAND_GATE U5689 ( .I1(n4807), .I2(n4814), .O(n4803) );
  NAND3_GATE U5690 ( .I1(n4558), .I2(n4557), .I3(n4803), .O(n4823) );
  NAND_GATE U5691 ( .I1(B[23]), .I2(A[8]), .O(n5513) );
  INV_GATE U5692 ( .I1(n4571), .O(n4568) );
  NAND4_GATE U5693 ( .I1(n4560), .I2(n4569), .I3(n4568), .I4(n4559), .O(n4577)
         );
  NAND3_GATE U5694 ( .I1(n3895), .I2(n4561), .I3(n4565), .O(n4562) );
  AND_GATE U5695 ( .I1(n4562), .I2(n4559), .O(n4564) );
  OR_GATE U5696 ( .I1(n4564), .I2(n4563), .O(n4576) );
  NAND_GATE U5697 ( .I1(n1142), .I2(n4565), .O(n4569) );
  NAND3_GATE U5698 ( .I1(n4569), .I2(n4568), .I3(n4559), .O(n4573) );
  NAND_GATE U5699 ( .I1(n4569), .I2(n4559), .O(n4570) );
  NAND_GATE U5700 ( .I1(n4571), .I2(n4570), .O(n4572) );
  NAND3_GATE U5701 ( .I1(n4574), .I2(n4573), .I3(n4572), .O(n4575) );
  NAND3_GATE U5702 ( .I1(n4577), .I2(n4576), .I3(n4575), .O(n4824) );
  NAND_GATE U5703 ( .I1(n5513), .I2(n4824), .O(n4578) );
  NAND_GATE U5704 ( .I1(n4823), .I2(n4578), .O(n4580) );
  INV_GATE U5705 ( .I1(n5513), .O(n4822) );
  NAND_GATE U5706 ( .I1(n4822), .I2(n813), .O(n4579) );
  NAND4_GATE U5707 ( .I1(n4590), .I2(n4584), .I3(n802), .I4(n4581), .O(n4591)
         );
  NAND4_GATE U5708 ( .I1(n4583), .I2(n4590), .I3(n4582), .I4(n802), .O(n4587)
         );
  NAND_GATE U5709 ( .I1(n4590), .I2(n4584), .O(n4586) );
  INV_GATE U5710 ( .I1(n4584), .O(n4589) );
  NAND3_GATE U5711 ( .I1(n4585), .I2(n4589), .I3(n608), .O(n4594) );
  NAND3_GATE U5712 ( .I1(n4585), .I2(n4584), .I3(n1311), .O(n4593) );
  NAND4_GATE U5713 ( .I1(n4587), .I2(n4586), .I3(n4594), .I4(n4593), .O(n4588)
         );
  NAND_GATE U5714 ( .I1(n4591), .I2(n4588), .O(n4833) );
  NAND_GATE U5715 ( .I1(B[23]), .I2(A[9]), .O(n4829) );
  INV_GATE U5716 ( .I1(n4829), .O(n4831) );
  NAND_GATE U5717 ( .I1(n608), .I2(n4589), .O(n4592) );
  NAND3_GATE U5718 ( .I1(n4592), .I2(n4591), .I3(n4590), .O(n4830) );
  NAND3_GATE U5719 ( .I1(n4831), .I2(n4830), .I3(n1156), .O(n4595) );
  NAND3_GATE U5720 ( .I1(n4598), .I2(n4597), .I3(n4842), .O(n4605) );
  INV_GATE U5721 ( .I1(n5375), .O(n4840) );
  AND3_GATE U5722 ( .I1(n4601), .I2(n4600), .I3(n4599), .O(n4603) );
  OR_GATE U5723 ( .I1(n4603), .I2(n4602), .O(n4841) );
  NAND_GATE U5724 ( .I1(n4840), .I2(n706), .O(n4604) );
  NAND_GATE U5725 ( .I1(n4605), .I2(n4604), .O(n5360) );
  NAND_GATE U5726 ( .I1(B[23]), .I2(A[11]), .O(n5364) );
  INV_GATE U5727 ( .I1(n4617), .O(n4619) );
  NAND4_GATE U5728 ( .I1(n4615), .I2(n4473), .I3(n4607), .I4(n4606), .O(n4612)
         );
  NAND4_GATE U5729 ( .I1(n4608), .I2(n4607), .I3(n4615), .I4(n4473), .O(n4611)
         );
  NAND_GATE U5730 ( .I1(n4615), .I2(n4609), .O(n4610) );
  NAND3_GATE U5731 ( .I1(n4612), .I2(n4611), .I3(n4610), .O(n4613) );
  NAND_GATE U5732 ( .I1(n4619), .I2(n4613), .O(n4628) );
  INV_GATE U5733 ( .I1(n4620), .O(n4618) );
  NAND4_GATE U5734 ( .I1(n4615), .I2(n4614), .I3(n1152), .I4(n4618), .O(n4627)
         );
  NAND_GATE U5735 ( .I1(n4628), .I2(n4627), .O(n4616) );
  NAND_GATE U5736 ( .I1(n5364), .I2(n4616), .O(n4622) );
  NAND_GATE U5737 ( .I1(n4618), .I2(n4617), .O(n4625) );
  NAND_GATE U5738 ( .I1(n4620), .I2(n4619), .O(n4624) );
  NAND4_GATE U5739 ( .I1(n4623), .I2(n5364), .I3(n4625), .I4(n4624), .O(n4621)
         );
  NAND3_GATE U5740 ( .I1(n5360), .I2(n4622), .I3(n4621), .O(n4630) );
  INV_GATE U5741 ( .I1(n5364), .O(n4850) );
  NAND3_GATE U5742 ( .I1(n4625), .I2(n4624), .I3(n4623), .O(n4626) );
  NAND_GATE U5743 ( .I1(n4850), .I2(n856), .O(n4629) );
  INV_GATE U5744 ( .I1(n4636), .O(n4638) );
  NAND3_GATE U5745 ( .I1(n4638), .I2(n4631), .I3(n4637), .O(n4634) );
  OR_GATE U5746 ( .I1(n4637), .I2(n4632), .O(n4633) );
  AND_GATE U5747 ( .I1(n4634), .I2(n4633), .O(n4643) );
  INV_GATE U5748 ( .I1(n4637), .O(n4635) );
  NAND_GATE U5749 ( .I1(n4636), .I2(n4635), .O(n4640) );
  NAND_GATE U5750 ( .I1(n4638), .I2(n4637), .O(n4639) );
  NAND3_GATE U5751 ( .I1(n4641), .I2(n4640), .I3(n4639), .O(n4642) );
  NAND_GATE U5752 ( .I1(n4643), .I2(n4642), .O(n4857) );
  NAND_GATE U5753 ( .I1(B[23]), .I2(A[12]), .O(n4856) );
  NAND_GATE U5754 ( .I1(n4857), .I2(n4856), .O(n4644) );
  NAND_GATE U5755 ( .I1(n4860), .I2(n4644), .O(n4646) );
  INV_GATE U5756 ( .I1(n4856), .O(n4864) );
  NAND_GATE U5757 ( .I1(n4859), .I2(n4864), .O(n4645) );
  NAND_GATE U5758 ( .I1(n4646), .I2(n4645), .O(n4719) );
  NAND_GATE U5759 ( .I1(n5326), .I2(n4717), .O(n4647) );
  NAND_GATE U5760 ( .I1(n4719), .I2(n4647), .O(n4648) );
  NAND_GATE U5761 ( .I1(n4649), .I2(n4648), .O(n4875) );
  NAND_GATE U5762 ( .I1(n4878), .I2(n5316), .O(n4650) );
  NAND_GATE U5763 ( .I1(n4875), .I2(n4650), .O(n4651) );
  NAND_GATE U5764 ( .I1(n4873), .I2(n4651), .O(n4888) );
  NAND_GATE U5765 ( .I1(n4890), .I2(n4894), .O(n4652) );
  NAND_GATE U5766 ( .I1(n4888), .I2(n4652), .O(n4653) );
  NAND_GATE U5767 ( .I1(n4884), .I2(n4653), .O(n4904) );
  NAND_GATE U5768 ( .I1(n4907), .I2(n4909), .O(n4654) );
  NAND_GATE U5769 ( .I1(n4904), .I2(n4654), .O(n4655) );
  NAND_GATE U5770 ( .I1(n4901), .I2(n4655), .O(n4920) );
  NAND_GATE U5771 ( .I1(n4922), .I2(n4925), .O(n4656) );
  NAND_GATE U5772 ( .I1(n4920), .I2(n4656), .O(n4657) );
  NAND_GATE U5773 ( .I1(n4916), .I2(n4657), .O(n4936) );
  NAND_GATE U5774 ( .I1(n4938), .I2(n4941), .O(n4658) );
  NAND_GATE U5775 ( .I1(n4936), .I2(n4658), .O(n4659) );
  NAND_GATE U5776 ( .I1(n4932), .I2(n4659), .O(n4951) );
  NAND_GATE U5777 ( .I1(n4953), .I2(n4956), .O(n4660) );
  NAND_GATE U5778 ( .I1(n4951), .I2(n4660), .O(n4661) );
  NAND_GATE U5779 ( .I1(n4947), .I2(n4661), .O(n4967) );
  NAND_GATE U5780 ( .I1(n4965), .I2(n4972), .O(n4662) );
  NAND_GATE U5781 ( .I1(n4967), .I2(n4662), .O(n4663) );
  NAND_GATE U5782 ( .I1(n4963), .I2(n4663), .O(n4983) );
  NAND_GATE U5783 ( .I1(n4981), .I2(n4988), .O(n4664) );
  NAND_GATE U5784 ( .I1(n4983), .I2(n4664), .O(n4665) );
  NAND_GATE U5785 ( .I1(n4979), .I2(n4665), .O(n4705) );
  NAND_GATE U5786 ( .I1(n4703), .I2(n4710), .O(n4666) );
  NAND_GATE U5787 ( .I1(n4705), .I2(n4666), .O(n4667) );
  NAND_GATE U5788 ( .I1(n4701), .I2(n4667), .O(n5001) );
  NAND_GATE U5789 ( .I1(n4999), .I2(n5006), .O(n4668) );
  NAND_GATE U5790 ( .I1(n5001), .I2(n4668), .O(n4669) );
  NAND_GATE U5791 ( .I1(n4997), .I2(n4669), .O(n5018) );
  NAND_GATE U5792 ( .I1(n5016), .I2(n5018), .O(n5013) );
  OR_GATE U5793 ( .I1(n4670), .I2(n4677), .O(n4673) );
  OR_GATE U5794 ( .I1(n4675), .I2(n4671), .O(n4672) );
  AND_GATE U5795 ( .I1(n4673), .I2(n4672), .O(n4682) );
  INV_GATE U5796 ( .I1(n4677), .O(n4674) );
  NAND_GATE U5797 ( .I1(n4674), .I2(n4675), .O(n4680) );
  INV_GATE U5798 ( .I1(n4675), .O(n4676) );
  NAND_GATE U5799 ( .I1(n4677), .I2(n4676), .O(n4679) );
  NAND3_GATE U5800 ( .I1(n4680), .I2(n4679), .I3(n4678), .O(n4681) );
  NAND_GATE U5801 ( .I1(n4682), .I2(n4681), .O(n5014) );
  INV_GATE U5802 ( .I1(n5014), .O(n5017) );
  INV_GATE U5803 ( .I1(n5018), .O(n5015) );
  NAND_GATE U5804 ( .I1(n5022), .I2(n5015), .O(n4683) );
  NAND_GATE U5805 ( .I1(n5017), .I2(n4683), .O(n4684) );
  NAND_GATE U5806 ( .I1(n5013), .I2(n4684), .O(n5033) );
  NAND_GATE U5807 ( .I1(n5031), .I2(n5038), .O(n4685) );
  NAND_GATE U5808 ( .I1(n5033), .I2(n4685), .O(n4686) );
  NAND_GATE U5809 ( .I1(n5029), .I2(n4686), .O(n5050) );
  NAND_GATE U5810 ( .I1(n5048), .I2(n5055), .O(n4687) );
  NAND_GATE U5811 ( .I1(n5050), .I2(n4687), .O(n4688) );
  NAND_GATE U5812 ( .I1(n5045), .I2(n4688), .O(n5067) );
  NAND_GATE U5813 ( .I1(n5065), .I2(n5072), .O(n4689) );
  NAND_GATE U5814 ( .I1(n5067), .I2(n4689), .O(n4690) );
  NAND_GATE U5815 ( .I1(n5062), .I2(n4690), .O(n5083) );
  NAND_GATE U5816 ( .I1(n5081), .I2(n5088), .O(n4691) );
  NAND_GATE U5817 ( .I1(n5083), .I2(n4691), .O(n4692) );
  NAND_GATE U5818 ( .I1(n5079), .I2(n4692), .O(n5100) );
  NAND_GATE U5819 ( .I1(n5098), .I2(n5105), .O(n4693) );
  NAND_GATE U5820 ( .I1(n5100), .I2(n4693), .O(n4694) );
  NAND_GATE U5821 ( .I1(n5095), .I2(n4694), .O(n5116) );
  NAND_GATE U5822 ( .I1(n5114), .I2(n5121), .O(n4695) );
  NAND_GATE U5823 ( .I1(n5116), .I2(n4695), .O(n4696) );
  NAND_GATE U5824 ( .I1(n5112), .I2(n4696), .O(n5132) );
  NAND_GATE U5825 ( .I1(n5130), .I2(n5137), .O(n4697) );
  NAND_GATE U5826 ( .I1(n5132), .I2(n4697), .O(n4698) );
  NAND_GATE U5827 ( .I1(n5128), .I2(n4698), .O(n4699) );
  NAND_GATE U5828 ( .I1(n286), .I2(n4699), .O(n15316) );
  AND_GATE U5829 ( .I1(n15316), .I2(n4700), .O(\A1[53] ) );
  NAND_GATE U5830 ( .I1(B[22]), .I2(A[31]), .O(n5152) );
  INV_GATE U5831 ( .I1(n5152), .O(n5126) );
  NAND_GATE U5832 ( .I1(B[22]), .I2(A[30]), .O(n5163) );
  INV_GATE U5833 ( .I1(n5163), .O(n5110) );
  NAND_GATE U5834 ( .I1(B[22]), .I2(A[29]), .O(n5174) );
  INV_GATE U5835 ( .I1(n5174), .O(n5093) );
  NAND_GATE U5836 ( .I1(B[22]), .I2(A[28]), .O(n5185) );
  INV_GATE U5837 ( .I1(n5185), .O(n5077) );
  NAND_GATE U5838 ( .I1(B[22]), .I2(A[27]), .O(n5196) );
  INV_GATE U5839 ( .I1(n5196), .O(n5060) );
  NAND_GATE U5840 ( .I1(B[22]), .I2(A[26]), .O(n5207) );
  INV_GATE U5841 ( .I1(n5207), .O(n5043) );
  NAND_GATE U5842 ( .I1(B[22]), .I2(A[25]), .O(n5217) );
  INV_GATE U5843 ( .I1(n5217), .O(n5027) );
  NAND_GATE U5844 ( .I1(B[22]), .I2(A[24]), .O(n5228) );
  INV_GATE U5845 ( .I1(n5228), .O(n5011) );
  NAND_GATE U5846 ( .I1(B[22]), .I2(A[23]), .O(n5241) );
  INV_GATE U5847 ( .I1(n5241), .O(n4995) );
  INV_GATE U5848 ( .I1(n4701), .O(n4702) );
  NAND_GATE U5849 ( .I1(n4702), .I2(n4705), .O(n4714) );
  NAND_GATE U5850 ( .I1(n4704), .I2(n4708), .O(n4712) );
  NAND_GATE U5851 ( .I1(n4706), .I2(n4705), .O(n4707) );
  NAND_GATE U5852 ( .I1(n4708), .I2(n4707), .O(n4709) );
  NAND_GATE U5853 ( .I1(n4710), .I2(n4709), .O(n4711) );
  NAND_GATE U5854 ( .I1(n4712), .I2(n4711), .O(n4713) );
  NAND_GATE U5855 ( .I1(n4714), .I2(n4713), .O(n5238) );
  NAND_GATE U5856 ( .I1(n4995), .I2(n5238), .O(n5234) );
  NAND_GATE U5857 ( .I1(B[22]), .I2(A[22]), .O(n5252) );
  INV_GATE U5858 ( .I1(n5252), .O(n4993) );
  NAND_GATE U5859 ( .I1(B[22]), .I2(A[21]), .O(n5590) );
  INV_GATE U5860 ( .I1(n5590), .O(n4977) );
  NAND_GATE U5861 ( .I1(B[22]), .I2(A[20]), .O(n5263) );
  INV_GATE U5862 ( .I1(n5263), .O(n4961) );
  NAND_GATE U5863 ( .I1(B[22]), .I2(A[19]), .O(n5274) );
  INV_GATE U5864 ( .I1(n5274), .O(n4945) );
  NAND_GATE U5865 ( .I1(B[22]), .I2(A[18]), .O(n5285) );
  INV_GATE U5866 ( .I1(n5285), .O(n4930) );
  NAND_GATE U5867 ( .I1(B[22]), .I2(A[17]), .O(n5572) );
  INV_GATE U5868 ( .I1(n5572), .O(n4914) );
  NAND_GATE U5869 ( .I1(B[22]), .I2(A[16]), .O(n5299) );
  INV_GATE U5870 ( .I1(n5299), .O(n4899) );
  NAND_GATE U5871 ( .I1(B[22]), .I2(A[15]), .O(n5321) );
  INV_GATE U5872 ( .I1(n5321), .O(n4882) );
  NAND_GATE U5873 ( .I1(B[22]), .I2(A[14]), .O(n5335) );
  INV_GATE U5874 ( .I1(n5335), .O(n4871) );
  NAND_GATE U5875 ( .I1(n4718), .I2(n4719), .O(n4716) );
  NAND_GATE U5876 ( .I1(n4717), .I2(n710), .O(n4715) );
  NAND_GATE U5877 ( .I1(n4716), .I2(n4715), .O(n5325) );
  NAND_GATE U5878 ( .I1(n4720), .I2(n4715), .O(n5327) );
  NAND_GATE U5879 ( .I1(n5332), .I2(n5327), .O(n4721) );
  NAND3_GATE U5880 ( .I1(n4720), .I2(n4719), .I3(n4718), .O(n5328) );
  NAND_GATE U5881 ( .I1(n4721), .I2(n5328), .O(n5336) );
  NAND_GATE U5882 ( .I1(B[22]), .I2(A[13]), .O(n5350) );
  INV_GATE U5883 ( .I1(n5350), .O(n5344) );
  NAND_GATE U5884 ( .I1(B[22]), .I2(A[11]), .O(n5387) );
  INV_GATE U5885 ( .I1(n5387), .O(n4845) );
  NAND_GATE U5886 ( .I1(B[22]), .I2(A[9]), .O(n5528) );
  INV_GATE U5887 ( .I1(n5528), .O(n5518) );
  NAND_GATE U5888 ( .I1(B[22]), .I2(A[6]), .O(n5752) );
  INV_GATE U5889 ( .I1(n5752), .O(n5743) );
  NAND4_GATE U5890 ( .I1(n676), .I2(n4723), .I3(n4729), .I4(n4722), .O(n5478)
         );
  NAND3_GATE U5891 ( .I1(n4725), .I2(n4737), .I3(n4724), .O(n4728) );
  NAND_GATE U5892 ( .I1(n4734), .I2(n4733), .O(n4729) );
  NAND_GATE U5893 ( .I1(n4728), .I2(n4729), .O(n4726) );
  NAND_GATE U5894 ( .I1(n4727), .I2(n4726), .O(n4732) );
  NAND3_GATE U5895 ( .I1(n4729), .I2(n4728), .I3(n676), .O(n4731) );
  NAND3_GATE U5896 ( .I1(n4732), .I2(n4731), .I3(n4730), .O(n4786) );
  NAND3_GATE U5897 ( .I1(n5478), .I2(n4786), .I3(n4787), .O(n5741) );
  INV_GATE U5898 ( .I1(n5741), .O(n5482) );
  NAND_GATE U5899 ( .I1(n5743), .I2(n5482), .O(n4789) );
  NAND3_GATE U5900 ( .I1(n4752), .I2(n4739), .I3(n4738), .O(n4740) );
  NAND_GATE U5901 ( .I1(n4741), .I2(n4740), .O(n5404) );
  INV_GATE U5902 ( .I1(n5404), .O(n4743) );
  NAND_GATE U5903 ( .I1(n4743), .I2(n5407), .O(n4758) );
  NAND_GATE U5904 ( .I1(B[22]), .I2(A[2]), .O(n5430) );
  INV_GATE U5905 ( .I1(n5430), .O(n5429) );
  NAND_GATE U5906 ( .I1(n1390), .I2(A[1]), .O(n4744) );
  NAND_GATE U5907 ( .I1(n14784), .I2(n4744), .O(n4745) );
  NAND_GATE U5908 ( .I1(B[23]), .I2(n4745), .O(n4749) );
  NAND_GATE U5909 ( .I1(n1389), .I2(A[0]), .O(n4746) );
  NAND_GATE U5910 ( .I1(n14781), .I2(n4746), .O(n4747) );
  NAND_GATE U5911 ( .I1(B[24]), .I2(n4747), .O(n4748) );
  NAND_GATE U5912 ( .I1(n4749), .I2(n4748), .O(n5431) );
  NAND_GATE U5913 ( .I1(n5429), .I2(n5431), .O(n5435) );
  NAND3_GATE U5914 ( .I1(B[22]), .I2(B[23]), .I3(n1196), .O(n5436) );
  NAND_GATE U5915 ( .I1(n5430), .I2(n174), .O(n4750) );
  NAND_GATE U5916 ( .I1(n1199), .I2(n4750), .O(n4751) );
  NAND_GATE U5917 ( .I1(n5435), .I2(n4751), .O(n5414) );
  NAND3_GATE U5918 ( .I1(n4755), .I2(n4752), .I3(n199), .O(n4757) );
  NAND3_GATE U5919 ( .I1(n4755), .I2(n4754), .I3(n4753), .O(n4756) );
  AND_GATE U5920 ( .I1(n4757), .I2(n4756), .O(n5405) );
  NAND3_GATE U5921 ( .I1(n4758), .I2(n5414), .I3(n5405), .O(n4760) );
  NAND_GATE U5922 ( .I1(B[22]), .I2(A[3]), .O(n5417) );
  INV_GATE U5923 ( .I1(n5417), .O(n5409) );
  NAND3_GATE U5924 ( .I1(n4758), .I2(n5409), .I3(n5405), .O(n4759) );
  NAND_GATE U5925 ( .I1(n5414), .I2(n5409), .O(n5408) );
  NAND3_GATE U5926 ( .I1(n4760), .I2(n4759), .I3(n5408), .O(n5443) );
  INV_GATE U5927 ( .I1(n4767), .O(n4765) );
  NAND3_GATE U5928 ( .I1(n4761), .I2(n4766), .I3(n4765), .O(n4764) );
  OR_GATE U5929 ( .I1(n4762), .I2(n4766), .O(n4763) );
  NAND_GATE U5930 ( .I1(n4764), .I2(n4763), .O(n4773) );
  NAND_GATE U5931 ( .I1(B[22]), .I2(A[4]), .O(n5719) );
  NAND_GATE U5932 ( .I1(n4773), .I2(n5719), .O(n4769) );
  NAND_GATE U5933 ( .I1(n4766), .I2(n4765), .O(n4772) );
  NAND4_GATE U5934 ( .I1(n5719), .I2(n4771), .I3(n4772), .I4(n4770), .O(n4768)
         );
  NAND3_GATE U5935 ( .I1(n5443), .I2(n4769), .I3(n4768), .O(n4776) );
  AND3_GATE U5936 ( .I1(n4772), .I2(n4771), .I3(n4770), .O(n4774) );
  OR_GATE U5937 ( .I1(n4774), .I2(n4773), .O(n5444) );
  INV_GATE U5938 ( .I1(n5444), .O(n5442) );
  NAND_GATE U5939 ( .I1(n614), .I2(n5442), .O(n4775) );
  NAND_GATE U5940 ( .I1(n4776), .I2(n4775), .O(n5467) );
  NAND3_GATE U5941 ( .I1(n4782), .I2(n5455), .I3(n1332), .O(n5458) );
  NAND_GATE U5942 ( .I1(n4782), .I2(n5455), .O(n4780) );
  NAND3_GATE U5943 ( .I1(n4778), .I2(n4777), .I3(n5455), .O(n4779) );
  NAND_GATE U5944 ( .I1(n4780), .I2(n4779), .O(n4781) );
  NAND_GATE U5945 ( .I1(n5458), .I2(n4781), .O(n5465) );
  NAND_GATE U5946 ( .I1(n4782), .I2(n1332), .O(n4783) );
  INV_GATE U5947 ( .I1(n4782), .O(n5453) );
  NAND_GATE U5948 ( .I1(n4783), .I2(n5454), .O(n5461) );
  NAND_GATE U5949 ( .I1(n5462), .I2(n5461), .O(n5451) );
  NAND3_GATE U5950 ( .I1(n5467), .I2(n5465), .I3(n5451), .O(n4785) );
  NAND_GATE U5951 ( .I1(B[22]), .I2(A[5]), .O(n5470) );
  INV_GATE U5952 ( .I1(n5470), .O(n5450) );
  NAND3_GATE U5953 ( .I1(n5450), .I2(n5465), .I3(n5451), .O(n4784) );
  NAND_GATE U5954 ( .I1(n5450), .I2(n5467), .O(n5457) );
  NAND3_GATE U5955 ( .I1(n4785), .I2(n4784), .I3(n5457), .O(n5483) );
  NAND3_GATE U5956 ( .I1(n5483), .I2(n5478), .I3(n1157), .O(n4788) );
  NAND_GATE U5957 ( .I1(n5743), .I2(n5483), .O(n5480) );
  NAND3_GATE U5958 ( .I1(n4789), .I2(n4788), .I3(n5480), .O(n5401) );
  INV_GATE U5959 ( .I1(n4791), .O(n4792) );
  NAND_GATE U5960 ( .I1(n4790), .I2(n4794), .O(n5390) );
  NAND3_GATE U5961 ( .I1(n4791), .I2(n854), .I3(n4790), .O(n5397) );
  NAND_GATE U5962 ( .I1(n854), .I2(n4791), .O(n4795) );
  NAND_GATE U5963 ( .I1(n4793), .I2(n4792), .O(n4794) );
  NAND_GATE U5964 ( .I1(n4795), .I2(n4794), .O(n5398) );
  NAND3_GATE U5965 ( .I1(n5401), .I2(n5402), .I3(n5403), .O(n4797) );
  NAND_GATE U5966 ( .I1(B[22]), .I2(A[7]), .O(n5491) );
  INV_GATE U5967 ( .I1(n5491), .O(n5394) );
  NAND3_GATE U5968 ( .I1(n5394), .I2(n5402), .I3(n5403), .O(n4796) );
  NAND_GATE U5969 ( .I1(n5394), .I2(n5401), .O(n5391) );
  NAND3_GATE U5970 ( .I1(n4797), .I2(n4796), .I3(n5391), .O(n5502) );
  NAND_GATE U5971 ( .I1(B[22]), .I2(A[8]), .O(n5503) );
  NAND_GATE U5972 ( .I1(n4799), .I2(n4798), .O(n4802) );
  NAND_GATE U5973 ( .I1(n4802), .I2(n4811), .O(n4806) );
  INV_GATE U5974 ( .I1(n4803), .O(n4804) );
  NAND3_GATE U5975 ( .I1(n4806), .I2(n4805), .I3(n4804), .O(n4809) );
  INV_GATE U5976 ( .I1(n4814), .O(n4810) );
  NAND4_GATE U5977 ( .I1(n4812), .I2(n4810), .I3(n4807), .I4(n4811), .O(n4808)
         );
  NAND3_GATE U5978 ( .I1(n4812), .I2(n4811), .I3(n4810), .O(n4816) );
  NAND_GATE U5979 ( .I1(n4812), .I2(n4811), .O(n4813) );
  NAND_GATE U5980 ( .I1(n4814), .I2(n4813), .O(n4815) );
  NAND3_GATE U5981 ( .I1(n4817), .I2(n4816), .I3(n4815), .O(n5498) );
  NAND_GATE U5982 ( .I1(n1238), .I2(n5498), .O(n5505) );
  NAND_GATE U5983 ( .I1(n5503), .I2(n5505), .O(n4818) );
  NAND_GATE U5984 ( .I1(n5502), .I2(n4818), .O(n4820) );
  INV_GATE U5985 ( .I1(n5503), .O(n5507) );
  INV_GATE U5986 ( .I1(n5505), .O(n5501) );
  NAND_GATE U5987 ( .I1(n5507), .I2(n5501), .O(n4819) );
  NAND_GATE U5988 ( .I1(n4820), .I2(n4819), .O(n5522) );
  INV_GATE U5989 ( .I1(n4823), .O(n4825) );
  NAND_GATE U5990 ( .I1(n4825), .I2(n4824), .O(n4821) );
  NAND_GATE U5991 ( .I1(n4822), .I2(n4821), .O(n5515) );
  NAND3_GATE U5992 ( .I1(n4823), .I2(n4822), .I3(n813), .O(n5516) );
  NAND_GATE U5993 ( .I1(n4823), .I2(n813), .O(n4826) );
  NAND_GATE U5994 ( .I1(n4826), .I2(n4821), .O(n5512) );
  NAND_GATE U5995 ( .I1(B[22]), .I2(A[10]), .O(n5535) );
  NAND_GATE U5996 ( .I1(n277), .I2(n4833), .O(n4827) );
  NAND3_GATE U5997 ( .I1(n4829), .I2(n4828), .I3(n4827), .O(n4836) );
  NAND4_GATE U5998 ( .I1(n4831), .I2(n4830), .I3(n277), .I4(n1156), .O(n4835)
         );
  OR_GATE U5999 ( .I1(n4833), .I2(n4832), .O(n4834) );
  NAND3_GATE U6000 ( .I1(n4836), .I2(n4835), .I3(n4834), .O(n5534) );
  NAND_GATE U6001 ( .I1(n5535), .I2(n5534), .O(n4837) );
  NAND_GATE U6002 ( .I1(n5532), .I2(n4837), .O(n4839) );
  INV_GATE U6003 ( .I1(n5535), .O(n5537) );
  INV_GATE U6004 ( .I1(n5534), .O(n5533) );
  NAND_GATE U6005 ( .I1(n5537), .I2(n5533), .O(n4838) );
  NAND_GATE U6006 ( .I1(n4839), .I2(n4838), .O(n5380) );
  NAND3_GATE U6007 ( .I1(n706), .I2(n4840), .I3(n4842), .O(n5378) );
  NAND_GATE U6008 ( .I1(n258), .I2(n4841), .O(n4844) );
  NAND_GATE U6009 ( .I1(n4842), .I2(n706), .O(n4843) );
  NAND_GATE U6010 ( .I1(n4844), .I2(n4843), .O(n5374) );
  NAND3_GATE U6011 ( .I1(n4845), .I2(n5372), .I3(n4846), .O(n5381) );
  NAND3_GATE U6012 ( .I1(n5380), .I2(n5372), .I3(n4846), .O(n5368) );
  NAND3_GATE U6013 ( .I1(n262), .I2(n5381), .I3(n5368), .O(n5366) );
  NAND3_GATE U6014 ( .I1(n5360), .I2(n4850), .I3(n856), .O(n5359) );
  NAND_GATE U6015 ( .I1(n4850), .I2(n4851), .O(n5358) );
  NAND3_GATE U6016 ( .I1(n5360), .I2(n856), .I3(n5364), .O(n4849) );
  NAND3_GATE U6017 ( .I1(n609), .I2(n600), .I3(n5364), .O(n4848) );
  NAND3_GATE U6018 ( .I1(n5358), .I2(n4849), .I3(n4848), .O(n4847) );
  NAND_GATE U6019 ( .I1(n5359), .I2(n4847), .O(n5355) );
  NAND_GATE U6020 ( .I1(n5366), .I2(n5355), .O(n4855) );
  NAND_GATE U6021 ( .I1(B[22]), .I2(A[12]), .O(n5554) );
  INV_GATE U6022 ( .I1(n5554), .O(n5356) );
  NAND_GATE U6023 ( .I1(n5366), .I2(n5356), .O(n4854) );
  NAND3_GATE U6024 ( .I1(n4851), .I2(n5359), .I3(n4850), .O(n4852) );
  AND_GATE U6025 ( .I1(n5356), .I2(n4852), .O(n5357) );
  NAND_GATE U6026 ( .I1(n1151), .I2(n5357), .O(n4853) );
  NAND3_GATE U6027 ( .I1(n4855), .I2(n4854), .I3(n4853), .O(n5349) );
  NAND_GATE U6028 ( .I1(n5344), .I2(n5349), .O(n4870) );
  NAND_GATE U6029 ( .I1(n740), .I2(n4857), .O(n4863) );
  NAND_GATE U6030 ( .I1(n4864), .I2(n4863), .O(n4858) );
  NAND3_GATE U6031 ( .I1(n4860), .I2(n4859), .I3(n4856), .O(n4866) );
  NAND3_GATE U6032 ( .I1(n740), .I2(n4857), .I3(n4856), .O(n4865) );
  NAND3_GATE U6033 ( .I1(n4858), .I2(n4866), .I3(n4865), .O(n4861) );
  NAND3_GATE U6034 ( .I1(n4860), .I2(n4864), .I3(n4859), .O(n4862) );
  NAND_GATE U6035 ( .I1(n4861), .I2(n4862), .O(n5347) );
  NAND_GATE U6036 ( .I1(n5349), .I2(n5347), .O(n4869) );
  NAND3_GATE U6037 ( .I1(n4864), .I2(n4863), .I3(n4862), .O(n4868) );
  AND_GATE U6038 ( .I1(n4866), .I2(n4865), .O(n4867) );
  NAND3_GATE U6039 ( .I1(n5344), .I2(n4868), .I3(n4867), .O(n5343) );
  NAND3_GATE U6040 ( .I1(n4870), .I2(n4869), .I3(n5343), .O(n5339) );
  NAND_GATE U6041 ( .I1(n5336), .I2(n5339), .O(n4872) );
  NAND_GATE U6042 ( .I1(n4871), .I2(n5339), .O(n5337) );
  NAND3_GATE U6043 ( .I1(n5338), .I2(n4872), .I3(n5337), .O(n5320) );
  NAND_GATE U6044 ( .I1(n4882), .I2(n5320), .O(n5308) );
  INV_GATE U6045 ( .I1(n4875), .O(n4877) );
  NAND_GATE U6046 ( .I1(n4874), .I2(n4879), .O(n5312) );
  NAND_GATE U6047 ( .I1(n4876), .I2(n4875), .O(n4880) );
  NAND_GATE U6048 ( .I1(n4878), .I2(n4877), .O(n4879) );
  NAND_GATE U6049 ( .I1(n4880), .I2(n4879), .O(n5315) );
  NAND_GATE U6050 ( .I1(n5312), .I2(n5317), .O(n4881) );
  NAND_GATE U6051 ( .I1(n5314), .I2(n4881), .O(n5309) );
  NAND_GATE U6052 ( .I1(n4882), .I2(n5309), .O(n5307) );
  NAND_GATE U6053 ( .I1(n5320), .I2(n5309), .O(n4883) );
  NAND_GATE U6054 ( .I1(n4899), .I2(n5298), .O(n5302) );
  INV_GATE U6055 ( .I1(n4884), .O(n4885) );
  NAND_GATE U6056 ( .I1(n4885), .I2(n4888), .O(n4898) );
  INV_GATE U6057 ( .I1(n4888), .O(n4889) );
  NAND_GATE U6058 ( .I1(n4890), .I2(n4889), .O(n4886) );
  NAND_GATE U6059 ( .I1(n4887), .I2(n4886), .O(n4896) );
  NAND_GATE U6060 ( .I1(n17), .I2(n4888), .O(n4892) );
  NAND_GATE U6061 ( .I1(n4892), .I2(n4891), .O(n4893) );
  NAND_GATE U6062 ( .I1(n4894), .I2(n4893), .O(n4895) );
  NAND_GATE U6063 ( .I1(n4896), .I2(n4895), .O(n4897) );
  NAND_GATE U6064 ( .I1(n4898), .I2(n4897), .O(n5303) );
  NAND_GATE U6065 ( .I1(n4899), .I2(n5303), .O(n5297) );
  NAND_GATE U6066 ( .I1(n5298), .I2(n5303), .O(n4900) );
  NAND3_GATE U6067 ( .I1(n5302), .I2(n5297), .I3(n4900), .O(n5290) );
  NAND_GATE U6068 ( .I1(n4914), .I2(n5290), .O(n5292) );
  INV_GATE U6069 ( .I1(n4901), .O(n4902) );
  NAND_GATE U6070 ( .I1(n4902), .I2(n4904), .O(n4913) );
  INV_GATE U6071 ( .I1(n4904), .O(n4906) );
  NAND_GATE U6072 ( .I1(n4903), .I2(n4908), .O(n4911) );
  NAND_GATE U6073 ( .I1(n4907), .I2(n4906), .O(n4908) );
  NAND_GATE U6074 ( .I1(n4911), .I2(n4910), .O(n4912) );
  NAND_GATE U6075 ( .I1(n4913), .I2(n4912), .O(n5291) );
  NAND_GATE U6076 ( .I1(n4914), .I2(n5291), .O(n5295) );
  NAND_GATE U6077 ( .I1(n5290), .I2(n5291), .O(n4915) );
  NAND3_GATE U6078 ( .I1(n5292), .I2(n5295), .I3(n4915), .O(n5284) );
  NAND_GATE U6079 ( .I1(n4930), .I2(n5284), .O(n5280) );
  INV_GATE U6080 ( .I1(n4916), .O(n4917) );
  NAND_GATE U6081 ( .I1(n4917), .I2(n4920), .O(n4929) );
  NAND_GATE U6082 ( .I1(n4919), .I2(n4918), .O(n4927) );
  NAND_GATE U6083 ( .I1(n4921), .I2(n4920), .O(n4923) );
  NAND_GATE U6084 ( .I1(n4923), .I2(n4918), .O(n4924) );
  NAND_GATE U6085 ( .I1(n4925), .I2(n4924), .O(n4926) );
  NAND_GATE U6086 ( .I1(n4927), .I2(n4926), .O(n4928) );
  NAND_GATE U6087 ( .I1(n4929), .I2(n4928), .O(n5283) );
  NAND_GATE U6088 ( .I1(n4930), .I2(n5283), .O(n5279) );
  NAND_GATE U6089 ( .I1(n5284), .I2(n5283), .O(n4931) );
  NAND3_GATE U6090 ( .I1(n5280), .I2(n5279), .I3(n4931), .O(n5273) );
  NAND_GATE U6091 ( .I1(n4945), .I2(n5273), .O(n5269) );
  INV_GATE U6092 ( .I1(n4932), .O(n4933) );
  NAND_GATE U6093 ( .I1(n4933), .I2(n4936), .O(n4944) );
  INV_GATE U6094 ( .I1(n4936), .O(n4937) );
  NAND_GATE U6095 ( .I1(n4938), .I2(n4937), .O(n4934) );
  NAND_GATE U6096 ( .I1(n4935), .I2(n4934), .O(n4943) );
  NAND_GATE U6097 ( .I1(n398), .I2(n4936), .O(n4939) );
  NAND_GATE U6098 ( .I1(n4939), .I2(n4934), .O(n4940) );
  NAND_GATE U6099 ( .I1(n4941), .I2(n4940), .O(n4942) );
  NAND_GATE U6100 ( .I1(n5273), .I2(n5272), .O(n4946) );
  NAND3_GATE U6101 ( .I1(n5269), .I2(n5268), .I3(n4946), .O(n5262) );
  NAND_GATE U6102 ( .I1(n4961), .I2(n5262), .O(n5258) );
  INV_GATE U6103 ( .I1(n4947), .O(n4948) );
  NAND_GATE U6104 ( .I1(n4948), .I2(n4951), .O(n4960) );
  NAND_GATE U6105 ( .I1(n4950), .I2(n4949), .O(n4958) );
  NAND_GATE U6106 ( .I1(n4952), .I2(n4951), .O(n4954) );
  NAND_GATE U6107 ( .I1(n4954), .I2(n4949), .O(n4955) );
  NAND_GATE U6108 ( .I1(n4956), .I2(n4955), .O(n4957) );
  NAND_GATE U6109 ( .I1(n4958), .I2(n4957), .O(n4959) );
  NAND_GATE U6110 ( .I1(n4960), .I2(n4959), .O(n5261) );
  NAND_GATE U6111 ( .I1(n4961), .I2(n5261), .O(n5257) );
  NAND_GATE U6112 ( .I1(n5262), .I2(n5261), .O(n4962) );
  NAND3_GATE U6113 ( .I1(n5258), .I2(n5257), .I3(n4962), .O(n5589) );
  NAND_GATE U6114 ( .I1(n4977), .I2(n5589), .O(n5583) );
  INV_GATE U6115 ( .I1(n4963), .O(n4964) );
  NAND_GATE U6116 ( .I1(n4964), .I2(n4967), .O(n4976) );
  NAND_GATE U6117 ( .I1(n4966), .I2(n4970), .O(n4974) );
  NAND_GATE U6118 ( .I1(n4968), .I2(n4967), .O(n4969) );
  NAND_GATE U6119 ( .I1(n4970), .I2(n4969), .O(n4971) );
  NAND_GATE U6120 ( .I1(n4972), .I2(n4971), .O(n4973) );
  NAND_GATE U6121 ( .I1(n4974), .I2(n4973), .O(n4975) );
  NAND_GATE U6122 ( .I1(n4976), .I2(n4975), .O(n5587) );
  NAND_GATE U6123 ( .I1(n4977), .I2(n5587), .O(n5582) );
  NAND_GATE U6124 ( .I1(n5589), .I2(n5587), .O(n4978) );
  NAND3_GATE U6125 ( .I1(n5583), .I2(n5582), .I3(n4978), .O(n5251) );
  NAND_GATE U6126 ( .I1(n4993), .I2(n5251), .O(n5247) );
  INV_GATE U6127 ( .I1(n4979), .O(n4980) );
  NAND_GATE U6128 ( .I1(n4980), .I2(n4983), .O(n4992) );
  NAND_GATE U6129 ( .I1(n4982), .I2(n4986), .O(n4990) );
  NAND_GATE U6130 ( .I1(n4984), .I2(n4983), .O(n4985) );
  NAND_GATE U6131 ( .I1(n4986), .I2(n4985), .O(n4987) );
  NAND_GATE U6132 ( .I1(n4988), .I2(n4987), .O(n4989) );
  NAND_GATE U6133 ( .I1(n4990), .I2(n4989), .O(n4991) );
  NAND_GATE U6134 ( .I1(n4992), .I2(n4991), .O(n5250) );
  NAND_GATE U6135 ( .I1(n4993), .I2(n5250), .O(n5246) );
  NAND_GATE U6136 ( .I1(n5251), .I2(n5250), .O(n4994) );
  NAND3_GATE U6137 ( .I1(n5247), .I2(n5246), .I3(n4994), .O(n5239) );
  NAND_GATE U6138 ( .I1(n4995), .I2(n5239), .O(n5233) );
  NAND_GATE U6139 ( .I1(n5238), .I2(n5239), .O(n4996) );
  NAND3_GATE U6140 ( .I1(n5234), .I2(n5233), .I3(n4996), .O(n5227) );
  NAND_GATE U6141 ( .I1(n5011), .I2(n5227), .O(n5223) );
  INV_GATE U6142 ( .I1(n4997), .O(n4998) );
  NAND_GATE U6143 ( .I1(n4998), .I2(n5001), .O(n5010) );
  NAND_GATE U6144 ( .I1(n5000), .I2(n5004), .O(n5008) );
  NAND_GATE U6145 ( .I1(n5002), .I2(n5001), .O(n5003) );
  NAND_GATE U6146 ( .I1(n5004), .I2(n5003), .O(n5005) );
  NAND_GATE U6147 ( .I1(n5006), .I2(n5005), .O(n5007) );
  NAND_GATE U6148 ( .I1(n5008), .I2(n5007), .O(n5009) );
  NAND_GATE U6149 ( .I1(n5010), .I2(n5009), .O(n5226) );
  NAND_GATE U6150 ( .I1(n5011), .I2(n5226), .O(n5222) );
  NAND_GATE U6151 ( .I1(n5227), .I2(n5226), .O(n5012) );
  NAND3_GATE U6152 ( .I1(n5223), .I2(n5222), .I3(n5012), .O(n5216) );
  NAND_GATE U6153 ( .I1(n5027), .I2(n5216), .O(n5212) );
  OR_GATE U6154 ( .I1(n5014), .I2(n5013), .O(n5026) );
  NAND_GATE U6155 ( .I1(n5015), .I2(n5014), .O(n5020) );
  NAND_GATE U6156 ( .I1(n5016), .I2(n5020), .O(n5024) );
  NAND_GATE U6157 ( .I1(n5018), .I2(n5017), .O(n5019) );
  NAND_GATE U6158 ( .I1(n5020), .I2(n5019), .O(n5021) );
  NAND_GATE U6159 ( .I1(n5022), .I2(n5021), .O(n5023) );
  NAND_GATE U6160 ( .I1(n5024), .I2(n5023), .O(n5025) );
  NAND_GATE U6161 ( .I1(n5026), .I2(n5025), .O(n5215) );
  NAND_GATE U6162 ( .I1(n5027), .I2(n5215), .O(n5211) );
  NAND_GATE U6163 ( .I1(n5216), .I2(n5215), .O(n5028) );
  NAND3_GATE U6164 ( .I1(n5212), .I2(n5211), .I3(n5028), .O(n5206) );
  NAND_GATE U6165 ( .I1(n5043), .I2(n5206), .O(n5202) );
  INV_GATE U6166 ( .I1(n5029), .O(n5030) );
  NAND_GATE U6167 ( .I1(n5030), .I2(n5033), .O(n5042) );
  NAND_GATE U6168 ( .I1(n5032), .I2(n5036), .O(n5040) );
  NAND_GATE U6169 ( .I1(n5034), .I2(n5033), .O(n5035) );
  NAND_GATE U6170 ( .I1(n5036), .I2(n5035), .O(n5037) );
  NAND_GATE U6171 ( .I1(n5038), .I2(n5037), .O(n5039) );
  NAND_GATE U6172 ( .I1(n5040), .I2(n5039), .O(n5041) );
  NAND_GATE U6173 ( .I1(n5042), .I2(n5041), .O(n5205) );
  NAND_GATE U6174 ( .I1(n5043), .I2(n5205), .O(n5201) );
  NAND_GATE U6175 ( .I1(n5206), .I2(n5205), .O(n5044) );
  NAND3_GATE U6176 ( .I1(n5202), .I2(n5201), .I3(n5044), .O(n5195) );
  NAND_GATE U6177 ( .I1(n5060), .I2(n5195), .O(n5191) );
  INV_GATE U6178 ( .I1(n5045), .O(n5046) );
  NAND_GATE U6179 ( .I1(n5046), .I2(n5050), .O(n5059) );
  INV_GATE U6180 ( .I1(n5050), .O(n5047) );
  NAND_GATE U6181 ( .I1(n5048), .I2(n5047), .O(n5053) );
  NAND_GATE U6182 ( .I1(n5049), .I2(n5053), .O(n5057) );
  NAND_GATE U6183 ( .I1(n5051), .I2(n5050), .O(n5052) );
  NAND_GATE U6184 ( .I1(n5053), .I2(n5052), .O(n5054) );
  NAND_GATE U6185 ( .I1(n5055), .I2(n5054), .O(n5056) );
  NAND_GATE U6186 ( .I1(n5057), .I2(n5056), .O(n5058) );
  NAND_GATE U6187 ( .I1(n5059), .I2(n5058), .O(n5194) );
  NAND_GATE U6188 ( .I1(n5060), .I2(n5194), .O(n5190) );
  NAND_GATE U6189 ( .I1(n5195), .I2(n5194), .O(n5061) );
  NAND3_GATE U6190 ( .I1(n5191), .I2(n5190), .I3(n5061), .O(n5184) );
  NAND_GATE U6191 ( .I1(n5077), .I2(n5184), .O(n5180) );
  INV_GATE U6192 ( .I1(n5062), .O(n5063) );
  NAND_GATE U6193 ( .I1(n5063), .I2(n5067), .O(n5076) );
  INV_GATE U6194 ( .I1(n5067), .O(n5064) );
  NAND_GATE U6195 ( .I1(n5065), .I2(n5064), .O(n5070) );
  NAND_GATE U6196 ( .I1(n5066), .I2(n5070), .O(n5074) );
  NAND_GATE U6197 ( .I1(n5068), .I2(n5067), .O(n5069) );
  NAND_GATE U6198 ( .I1(n5070), .I2(n5069), .O(n5071) );
  NAND_GATE U6199 ( .I1(n5072), .I2(n5071), .O(n5073) );
  NAND_GATE U6200 ( .I1(n5074), .I2(n5073), .O(n5075) );
  NAND_GATE U6201 ( .I1(n5076), .I2(n5075), .O(n5183) );
  NAND_GATE U6202 ( .I1(n5077), .I2(n5183), .O(n5179) );
  NAND_GATE U6203 ( .I1(n5184), .I2(n5183), .O(n5078) );
  NAND3_GATE U6204 ( .I1(n5180), .I2(n5179), .I3(n5078), .O(n5173) );
  NAND_GATE U6205 ( .I1(n5093), .I2(n5173), .O(n5169) );
  INV_GATE U6206 ( .I1(n5079), .O(n5080) );
  NAND_GATE U6207 ( .I1(n5080), .I2(n5083), .O(n5092) );
  NAND_GATE U6208 ( .I1(n5082), .I2(n5086), .O(n5090) );
  NAND_GATE U6209 ( .I1(n5084), .I2(n5083), .O(n5085) );
  NAND_GATE U6210 ( .I1(n5086), .I2(n5085), .O(n5087) );
  NAND_GATE U6211 ( .I1(n5088), .I2(n5087), .O(n5089) );
  NAND_GATE U6212 ( .I1(n5090), .I2(n5089), .O(n5091) );
  NAND_GATE U6213 ( .I1(n5092), .I2(n5091), .O(n5172) );
  NAND_GATE U6214 ( .I1(n5093), .I2(n5172), .O(n5168) );
  NAND_GATE U6215 ( .I1(n5173), .I2(n5172), .O(n5094) );
  NAND3_GATE U6216 ( .I1(n5169), .I2(n5168), .I3(n5094), .O(n5162) );
  NAND_GATE U6217 ( .I1(n5110), .I2(n5162), .O(n5158) );
  INV_GATE U6218 ( .I1(n5095), .O(n5096) );
  NAND_GATE U6219 ( .I1(n5096), .I2(n5100), .O(n5109) );
  INV_GATE U6220 ( .I1(n5100), .O(n5097) );
  NAND_GATE U6221 ( .I1(n5098), .I2(n5097), .O(n5103) );
  NAND_GATE U6222 ( .I1(n5099), .I2(n5103), .O(n5107) );
  NAND_GATE U6223 ( .I1(n5101), .I2(n5100), .O(n5102) );
  NAND_GATE U6224 ( .I1(n5103), .I2(n5102), .O(n5104) );
  NAND_GATE U6225 ( .I1(n5105), .I2(n5104), .O(n5106) );
  NAND_GATE U6226 ( .I1(n5107), .I2(n5106), .O(n5108) );
  NAND_GATE U6227 ( .I1(n5109), .I2(n5108), .O(n5161) );
  NAND_GATE U6228 ( .I1(n5110), .I2(n5161), .O(n5157) );
  NAND_GATE U6229 ( .I1(n5162), .I2(n5161), .O(n5111) );
  NAND3_GATE U6230 ( .I1(n5158), .I2(n5157), .I3(n5111), .O(n5151) );
  NAND_GATE U6231 ( .I1(n5126), .I2(n5151), .O(n5147) );
  INV_GATE U6232 ( .I1(n5112), .O(n5113) );
  NAND_GATE U6233 ( .I1(n5113), .I2(n5116), .O(n5125) );
  NAND_GATE U6234 ( .I1(n5115), .I2(n5119), .O(n5123) );
  NAND_GATE U6235 ( .I1(n5117), .I2(n5116), .O(n5118) );
  NAND_GATE U6236 ( .I1(n5119), .I2(n5118), .O(n5120) );
  NAND_GATE U6237 ( .I1(n5121), .I2(n5120), .O(n5122) );
  NAND_GATE U6238 ( .I1(n5123), .I2(n5122), .O(n5124) );
  NAND_GATE U6239 ( .I1(n5125), .I2(n5124), .O(n5150) );
  NAND_GATE U6240 ( .I1(n5126), .I2(n5150), .O(n5146) );
  NAND_GATE U6241 ( .I1(n5151), .I2(n5150), .O(n5127) );
  NAND3_GATE U6242 ( .I1(n5147), .I2(n5146), .I3(n5127), .O(n15318) );
  INV_GATE U6243 ( .I1(n15318), .O(n5142) );
  INV_GATE U6244 ( .I1(n5128), .O(n5129) );
  NAND_GATE U6245 ( .I1(n5129), .I2(n5132), .O(n5141) );
  NAND_GATE U6246 ( .I1(n5131), .I2(n5135), .O(n5139) );
  NAND_GATE U6247 ( .I1(n5133), .I2(n5132), .O(n5134) );
  NAND_GATE U6248 ( .I1(n5135), .I2(n5134), .O(n5136) );
  NAND_GATE U6249 ( .I1(n5137), .I2(n5136), .O(n5138) );
  NAND_GATE U6250 ( .I1(n5139), .I2(n5138), .O(n5140) );
  NAND_GATE U6251 ( .I1(n5141), .I2(n5140), .O(n15317) );
  NAND_GATE U6252 ( .I1(n5142), .I2(n15317), .O(n5145) );
  INV_GATE U6253 ( .I1(n15317), .O(n5143) );
  NAND_GATE U6254 ( .I1(n15318), .I2(n5143), .O(n5144) );
  NAND_GATE U6255 ( .I1(n5145), .I2(n5144), .O(\A1[52] ) );
  OR_GATE U6256 ( .I1(n5146), .I2(n5151), .O(n5149) );
  OR_GATE U6257 ( .I1(n5150), .I2(n5147), .O(n5148) );
  AND_GATE U6258 ( .I1(n5149), .I2(n5148), .O(n5156) );
  NAND_GATE U6259 ( .I1(n1122), .I2(n5150), .O(n5154) );
  NAND3_GATE U6260 ( .I1(n5154), .I2(n5153), .I3(n5152), .O(n5155) );
  NAND_GATE U6261 ( .I1(n5156), .I2(n5155), .O(n5618) );
  INV_GATE U6262 ( .I1(n5618), .O(n5615) );
  OR_GATE U6263 ( .I1(n5157), .I2(n5162), .O(n5160) );
  OR_GATE U6264 ( .I1(n5161), .I2(n5158), .O(n5159) );
  AND_GATE U6265 ( .I1(n5160), .I2(n5159), .O(n5167) );
  NAND_GATE U6266 ( .I1(n1114), .I2(n5161), .O(n5165) );
  NAND3_GATE U6267 ( .I1(n5165), .I2(n5164), .I3(n5163), .O(n5166) );
  NAND_GATE U6268 ( .I1(n5167), .I2(n5166), .O(n6061) );
  INV_GATE U6269 ( .I1(n6061), .O(n6064) );
  NAND_GATE U6270 ( .I1(B[21]), .I2(A[31]), .O(n6068) );
  INV_GATE U6271 ( .I1(n6068), .O(n6062) );
  NAND_GATE U6272 ( .I1(n6064), .I2(n6062), .O(n6058) );
  OR_GATE U6273 ( .I1(n5168), .I2(n5173), .O(n5171) );
  OR_GATE U6274 ( .I1(n5172), .I2(n5169), .O(n5170) );
  AND_GATE U6275 ( .I1(n5171), .I2(n5170), .O(n5178) );
  NAND_GATE U6276 ( .I1(n1107), .I2(n5172), .O(n5176) );
  NAND3_GATE U6277 ( .I1(n5176), .I2(n5175), .I3(n5174), .O(n5177) );
  NAND_GATE U6278 ( .I1(n5178), .I2(n5177), .O(n6044) );
  INV_GATE U6279 ( .I1(n6044), .O(n6047) );
  NAND_GATE U6280 ( .I1(B[21]), .I2(A[30]), .O(n6051) );
  INV_GATE U6281 ( .I1(n6051), .O(n6045) );
  NAND_GATE U6282 ( .I1(n6047), .I2(n6045), .O(n6041) );
  OR_GATE U6283 ( .I1(n5179), .I2(n5184), .O(n5182) );
  OR_GATE U6284 ( .I1(n5183), .I2(n5180), .O(n5181) );
  AND_GATE U6285 ( .I1(n5182), .I2(n5181), .O(n5189) );
  NAND_GATE U6286 ( .I1(n1101), .I2(n5183), .O(n5187) );
  NAND3_GATE U6287 ( .I1(n5187), .I2(n5186), .I3(n5185), .O(n5188) );
  NAND_GATE U6288 ( .I1(n5189), .I2(n5188), .O(n6027) );
  INV_GATE U6289 ( .I1(n6027), .O(n6030) );
  NAND_GATE U6290 ( .I1(B[21]), .I2(A[29]), .O(n6034) );
  INV_GATE U6291 ( .I1(n6034), .O(n6028) );
  NAND_GATE U6292 ( .I1(n6030), .I2(n6028), .O(n6024) );
  OR_GATE U6293 ( .I1(n5190), .I2(n5195), .O(n5193) );
  OR_GATE U6294 ( .I1(n5194), .I2(n5191), .O(n5192) );
  AND_GATE U6295 ( .I1(n5193), .I2(n5192), .O(n5200) );
  NAND_GATE U6296 ( .I1(n1091), .I2(n5194), .O(n5198) );
  NAND3_GATE U6297 ( .I1(n5198), .I2(n5197), .I3(n5196), .O(n5199) );
  NAND_GATE U6298 ( .I1(n5200), .I2(n5199), .O(n6014) );
  INV_GATE U6299 ( .I1(n6014), .O(n6017) );
  NAND_GATE U6300 ( .I1(B[21]), .I2(A[28]), .O(n6108) );
  INV_GATE U6301 ( .I1(n6108), .O(n6015) );
  NAND_GATE U6302 ( .I1(n6017), .I2(n6015), .O(n6013) );
  OR_GATE U6303 ( .I1(n5201), .I2(n5206), .O(n5204) );
  OR_GATE U6304 ( .I1(n5205), .I2(n5202), .O(n5203) );
  NAND_GATE U6305 ( .I1(n1059), .I2(n5205), .O(n5209) );
  NAND3_GATE U6306 ( .I1(n5209), .I2(n5208), .I3(n5207), .O(n5210) );
  INV_GATE U6307 ( .I1(n5996), .O(n5997) );
  NAND_GATE U6308 ( .I1(B[21]), .I2(A[27]), .O(n6007) );
  INV_GATE U6309 ( .I1(n6007), .O(n6000) );
  NAND_GATE U6310 ( .I1(n5997), .I2(n6000), .O(n6001) );
  OR_GATE U6311 ( .I1(n5211), .I2(n5216), .O(n5214) );
  OR_GATE U6312 ( .I1(n5215), .I2(n5212), .O(n5213) );
  AND_GATE U6313 ( .I1(n5214), .I2(n5213), .O(n5221) );
  NAND_GATE U6314 ( .I1(n5216), .I2(n1075), .O(n5218) );
  NAND3_GATE U6315 ( .I1(n5219), .I2(n5218), .I3(n5217), .O(n5220) );
  NAND_GATE U6316 ( .I1(n5221), .I2(n5220), .O(n5979) );
  INV_GATE U6317 ( .I1(n5979), .O(n5980) );
  NAND_GATE U6318 ( .I1(B[21]), .I2(A[26]), .O(n5990) );
  INV_GATE U6319 ( .I1(n5990), .O(n5983) );
  NAND_GATE U6320 ( .I1(n5980), .I2(n5983), .O(n5984) );
  OR_GATE U6321 ( .I1(n5222), .I2(n5227), .O(n5225) );
  OR_GATE U6322 ( .I1(n5226), .I2(n5223), .O(n5224) );
  AND_GATE U6323 ( .I1(n5225), .I2(n5224), .O(n5232) );
  NAND_GATE U6324 ( .I1(n1076), .I2(n5226), .O(n5230) );
  NAND3_GATE U6325 ( .I1(n5230), .I2(n5229), .I3(n5228), .O(n5231) );
  NAND_GATE U6326 ( .I1(n5232), .I2(n5231), .O(n5962) );
  INV_GATE U6327 ( .I1(n5962), .O(n5963) );
  NAND_GATE U6328 ( .I1(B[21]), .I2(A[25]), .O(n5973) );
  INV_GATE U6329 ( .I1(n5973), .O(n5966) );
  NAND_GATE U6330 ( .I1(n5963), .I2(n5966), .O(n5967) );
  OR_GATE U6331 ( .I1(n5233), .I2(n5238), .O(n5236) );
  OR_GATE U6332 ( .I1(n5239), .I2(n5234), .O(n5235) );
  AND_GATE U6333 ( .I1(n5236), .I2(n5235), .O(n5245) );
  INV_GATE U6334 ( .I1(n5239), .O(n5237) );
  NAND_GATE U6335 ( .I1(n5238), .I2(n5237), .O(n5243) );
  INV_GATE U6336 ( .I1(n5238), .O(n5240) );
  NAND_GATE U6337 ( .I1(n5240), .I2(n5239), .O(n5242) );
  NAND3_GATE U6338 ( .I1(n5243), .I2(n5242), .I3(n5241), .O(n5244) );
  NAND_GATE U6339 ( .I1(n5245), .I2(n5244), .O(n5945) );
  INV_GATE U6340 ( .I1(n5945), .O(n5946) );
  NAND_GATE U6341 ( .I1(B[21]), .I2(A[24]), .O(n5956) );
  INV_GATE U6342 ( .I1(n5956), .O(n5949) );
  NAND_GATE U6343 ( .I1(n5946), .I2(n5949), .O(n5950) );
  OR_GATE U6344 ( .I1(n5246), .I2(n5251), .O(n5249) );
  OR_GATE U6345 ( .I1(n5250), .I2(n5247), .O(n5248) );
  AND_GATE U6346 ( .I1(n5249), .I2(n5248), .O(n5256) );
  NAND_GATE U6347 ( .I1(n1077), .I2(n5250), .O(n5254) );
  NAND3_GATE U6348 ( .I1(n5254), .I2(n5253), .I3(n5252), .O(n5255) );
  NAND_GATE U6349 ( .I1(n5256), .I2(n5255), .O(n5928) );
  INV_GATE U6350 ( .I1(n5928), .O(n5929) );
  NAND_GATE U6351 ( .I1(B[21]), .I2(A[23]), .O(n5940) );
  INV_GATE U6352 ( .I1(n5940), .O(n5932) );
  NAND_GATE U6353 ( .I1(n5929), .I2(n5932), .O(n5933) );
  NAND_GATE U6354 ( .I1(B[21]), .I2(A[22]), .O(n5923) );
  INV_GATE U6355 ( .I1(n5923), .O(n5915) );
  OR_GATE U6356 ( .I1(n5257), .I2(n5262), .O(n5260) );
  OR_GATE U6357 ( .I1(n5261), .I2(n5258), .O(n5259) );
  AND_GATE U6358 ( .I1(n5260), .I2(n5259), .O(n5267) );
  NAND_GATE U6359 ( .I1(n392), .I2(n5261), .O(n5265) );
  NAND3_GATE U6360 ( .I1(n5265), .I2(n5264), .I3(n5263), .O(n5266) );
  NAND_GATE U6361 ( .I1(n5267), .I2(n5266), .O(n5896) );
  NAND_GATE U6362 ( .I1(B[21]), .I2(A[21]), .O(n5905) );
  INV_GATE U6363 ( .I1(n5905), .O(n5898) );
  NAND_GATE U6364 ( .I1(n564), .I2(n5898), .O(n5899) );
  OR_GATE U6365 ( .I1(n5268), .I2(n5273), .O(n5271) );
  OR_GATE U6366 ( .I1(n5272), .I2(n5269), .O(n5270) );
  AND_GATE U6367 ( .I1(n5271), .I2(n5270), .O(n5278) );
  NAND_GATE U6368 ( .I1(n1038), .I2(n5272), .O(n5276) );
  NAND3_GATE U6369 ( .I1(n5276), .I2(n5275), .I3(n5274), .O(n5277) );
  NAND_GATE U6370 ( .I1(B[21]), .I2(A[20]), .O(n5888) );
  INV_GATE U6371 ( .I1(n5888), .O(n5624) );
  NAND_GATE U6372 ( .I1(n583), .I2(n5624), .O(n5625) );
  OR_GATE U6373 ( .I1(n5283), .I2(n5280), .O(n5281) );
  AND_GATE U6374 ( .I1(n5282), .I2(n5281), .O(n5289) );
  NAND_GATE U6375 ( .I1(n1039), .I2(n5283), .O(n5287) );
  NAND3_GATE U6376 ( .I1(n5287), .I2(n5286), .I3(n5285), .O(n5288) );
  NAND_GATE U6377 ( .I1(n5289), .I2(n5288), .O(n5876) );
  INV_GATE U6378 ( .I1(n5876), .O(n5872) );
  NAND_GATE U6379 ( .I1(B[21]), .I2(A[19]), .O(n6212) );
  INV_GATE U6380 ( .I1(n6212), .O(n5877) );
  NAND_GATE U6381 ( .I1(n5872), .I2(n5877), .O(n5878) );
  INV_GATE U6382 ( .I1(n5291), .O(n5293) );
  NAND_GATE U6383 ( .I1(n875), .I2(n5291), .O(n5570) );
  NAND3_GATE U6384 ( .I1(n5572), .I2(n5571), .I3(n5570), .O(n5296) );
  INV_GATE U6385 ( .I1(n5292), .O(n5294) );
  NAND_GATE U6386 ( .I1(n5294), .I2(n5293), .O(n5568) );
  NAND_GATE U6387 ( .I1(B[21]), .I2(A[18]), .O(n5864) );
  INV_GATE U6388 ( .I1(n5864), .O(n5855) );
  NAND_GATE U6389 ( .I1(n788), .I2(n5855), .O(n5856) );
  OR_GATE U6390 ( .I1(n5297), .I2(n5298), .O(n5306) );
  NAND_GATE U6391 ( .I1(n681), .I2(n5303), .O(n5301) );
  NAND3_GATE U6392 ( .I1(n5301), .I2(n5300), .I3(n5299), .O(n5305) );
  OR_GATE U6393 ( .I1(n5303), .I2(n5302), .O(n5304) );
  NAND3_GATE U6394 ( .I1(n5306), .I2(n5305), .I3(n5304), .O(n5846) );
  NAND_GATE U6395 ( .I1(B[21]), .I2(A[17]), .O(n6226) );
  INV_GATE U6396 ( .I1(n6226), .O(n5845) );
  NAND_GATE U6397 ( .I1(n545), .I2(n5845), .O(n5844) );
  OR_GATE U6398 ( .I1(n5309), .I2(n5308), .O(n5310) );
  INV_GATE U6399 ( .I1(n5312), .O(n5313) );
  NAND_GATE U6400 ( .I1(n5314), .I2(n5313), .O(n5318) );
  NAND_GATE U6401 ( .I1(n5316), .I2(n5315), .O(n5317) );
  NAND_GATE U6402 ( .I1(n5318), .I2(n5317), .O(n5319) );
  NAND_GATE U6403 ( .I1(n5320), .I2(n5319), .O(n5322) );
  NAND3_GATE U6404 ( .I1(n5323), .I2(n5322), .I3(n5321), .O(n5324) );
  INV_GATE U6405 ( .I1(n5834), .O(n5833) );
  NAND_GATE U6406 ( .I1(B[21]), .I2(A[16]), .O(n5831) );
  INV_GATE U6407 ( .I1(n5831), .O(n5836) );
  NAND_GATE U6408 ( .I1(B[21]), .I2(A[15]), .O(n6254) );
  INV_GATE U6409 ( .I1(n6254), .O(n5634) );
  NAND_GATE U6410 ( .I1(n5326), .I2(n5325), .O(n5332) );
  NAND_GATE U6411 ( .I1(n5332), .I2(n5331), .O(n5329) );
  NAND_GATE U6412 ( .I1(n5339), .I2(n5329), .O(n5334) );
  INV_GATE U6413 ( .I1(n5339), .O(n5330) );
  NAND3_GATE U6414 ( .I1(n5332), .I2(n5331), .I3(n5330), .O(n5333) );
  NAND3_GATE U6415 ( .I1(n5335), .I2(n5334), .I3(n5333), .O(n5342) );
  OR_GATE U6416 ( .I1(n5337), .I2(n5336), .O(n5341) );
  OR_GATE U6417 ( .I1(n5339), .I2(n5338), .O(n5340) );
  NAND3_GATE U6418 ( .I1(n5342), .I2(n5341), .I3(n5340), .O(n5631) );
  NAND_GATE U6419 ( .I1(n5634), .I2(n709), .O(n5563) );
  OR_GATE U6420 ( .I1(n5343), .I2(n5349), .O(n5346) );
  INV_GATE U6421 ( .I1(n5347), .O(n5348) );
  NAND3_GATE U6422 ( .I1(n5348), .I2(n5349), .I3(n5344), .O(n5345) );
  AND_GATE U6423 ( .I1(n5346), .I2(n5345), .O(n5354) );
  NAND_GATE U6424 ( .I1(n3), .I2(n5347), .O(n5352) );
  NAND_GATE U6425 ( .I1(n5349), .I2(n5348), .O(n5351) );
  NAND3_GATE U6426 ( .I1(n5352), .I2(n5351), .I3(n5350), .O(n5353) );
  NAND_GATE U6427 ( .I1(n5354), .I2(n5353), .O(n5821) );
  INV_GATE U6428 ( .I1(n5821), .O(n5818) );
  NAND_GATE U6429 ( .I1(B[21]), .I2(A[14]), .O(n5819) );
  INV_GATE U6430 ( .I1(n5819), .O(n5816) );
  NAND_GATE U6431 ( .I1(n5818), .I2(n5816), .O(n5814) );
  NAND_GATE U6432 ( .I1(B[21]), .I2(A[13]), .O(n6280) );
  INV_GATE U6433 ( .I1(n6280), .O(n5808) );
  NAND_GATE U6434 ( .I1(n5360), .I2(n856), .O(n5362) );
  NAND_GATE U6435 ( .I1(n609), .I2(n600), .O(n5361) );
  NAND_GATE U6436 ( .I1(n5362), .I2(n5361), .O(n5363) );
  NAND_GATE U6437 ( .I1(n5364), .I2(n5363), .O(n5369) );
  NAND_GATE U6438 ( .I1(n5367), .I2(n5369), .O(n5365) );
  NAND_GATE U6439 ( .I1(n5366), .I2(n5365), .O(n5553) );
  NAND5_GATE U6440 ( .I1(n262), .I2(n5381), .I3(n5369), .I4(n5368), .I5(n5367), 
        .O(n5552) );
  NAND3_GATE U6441 ( .I1(n5554), .I2(n5553), .I3(n5552), .O(n5370) );
  NAND_GATE U6442 ( .I1(n5808), .I2(n5810), .O(n5558) );
  NAND_GATE U6443 ( .I1(B[21]), .I2(A[12]), .O(n6472) );
  INV_GATE U6444 ( .I1(n6472), .O(n5803) );
  NAND_GATE U6445 ( .I1(n634), .I2(n5378), .O(n5372) );
  NAND3_GATE U6446 ( .I1(n5371), .I2(n5372), .I3(n574), .O(n5385) );
  NAND_GATE U6447 ( .I1(n5372), .I2(n5371), .O(n5373) );
  NAND_GATE U6448 ( .I1(n5380), .I2(n5373), .O(n5386) );
  AND3_GATE U6449 ( .I1(n5385), .I2(n5387), .I3(n5386), .O(n5384) );
  NAND_GATE U6450 ( .I1(n5375), .I2(n5374), .O(n5376) );
  NAND_GATE U6451 ( .I1(n5377), .I2(n5376), .O(n5379) );
  NAND3_GATE U6452 ( .I1(n5379), .I2(n1270), .I3(n5378), .O(n5383) );
  OR_GATE U6453 ( .I1(n5381), .I2(n5380), .O(n5382) );
  NAND_GATE U6454 ( .I1(n5383), .I2(n5382), .O(n5388) );
  OR_GATE U6455 ( .I1(n5384), .I2(n5388), .O(n6473) );
  NAND_GATE U6456 ( .I1(n5803), .I2(n619), .O(n5548) );
  NAND4_GATE U6457 ( .I1(n5387), .I2(n6472), .I3(n5386), .I4(n5385), .O(n5546)
         );
  NAND_GATE U6458 ( .I1(n6472), .I2(n5388), .O(n5545) );
  NAND_GATE U6459 ( .I1(B[21]), .I2(A[11]), .O(n5645) );
  INV_GATE U6460 ( .I1(n5645), .O(n5638) );
  NAND_GATE U6461 ( .I1(B[21]), .I2(A[9]), .O(n5785) );
  INV_GATE U6462 ( .I1(n5785), .O(n5654) );
  NAND_GATE U6463 ( .I1(B[21]), .I2(A[8]), .O(n5767) );
  INV_GATE U6464 ( .I1(n5767), .O(n5777) );
  NAND_GATE U6465 ( .I1(n5390), .I2(n5389), .O(n5393) );
  INV_GATE U6466 ( .I1(n5391), .O(n5392) );
  NAND3_GATE U6467 ( .I1(n5397), .I2(n5393), .I3(n5392), .O(n5396) );
  NAND4_GATE U6468 ( .I1(n5394), .I2(n5402), .I3(n675), .I4(n5403), .O(n5395)
         );
  NAND_GATE U6469 ( .I1(n5396), .I2(n5395), .O(n5492) );
  NAND_GATE U6470 ( .I1(n5399), .I2(n5398), .O(n5403) );
  NAND_GATE U6471 ( .I1(n5402), .I2(n5403), .O(n5400) );
  NAND_GATE U6472 ( .I1(n5401), .I2(n5400), .O(n5489) );
  NAND3_GATE U6473 ( .I1(n5403), .I2(n5402), .I3(n675), .O(n5490) );
  NAND3_GATE U6474 ( .I1(n5489), .I2(n5490), .I3(n5491), .O(n5771) );
  NAND_GATE U6475 ( .I1(n5777), .I2(n823), .O(n5496) );
  NAND_GATE U6476 ( .I1(B[21]), .I2(A[5]), .O(n5725) );
  INV_GATE U6477 ( .I1(n5725), .O(n5723) );
  NAND_GATE U6478 ( .I1(B[21]), .I2(A[4]), .O(n5694) );
  NAND_GATE U6479 ( .I1(n5405), .I2(n5404), .O(n5406) );
  NAND_GATE U6480 ( .I1(n5407), .I2(n5406), .O(n5413) );
  OR_GATE U6481 ( .I1(n5413), .I2(n5408), .O(n5411) );
  INV_GATE U6482 ( .I1(n5414), .O(n5412) );
  NAND3_GATE U6483 ( .I1(n5412), .I2(n5409), .I3(n5413), .O(n5410) );
  AND_GATE U6484 ( .I1(n5411), .I2(n5410), .O(n5419) );
  NAND_GATE U6485 ( .I1(n5412), .I2(n5413), .O(n5416) );
  NAND3_GATE U6486 ( .I1(n5417), .I2(n5416), .I3(n5415), .O(n5418) );
  NAND_GATE U6487 ( .I1(n5419), .I2(n5418), .O(n5696) );
  NAND_GATE U6488 ( .I1(B[21]), .I2(A[2]), .O(n5679) );
  INV_GATE U6489 ( .I1(n5679), .O(n5684) );
  NAND_GATE U6490 ( .I1(n1388), .I2(A[0]), .O(n5420) );
  NAND_GATE U6491 ( .I1(n14781), .I2(n5420), .O(n5421) );
  NAND_GATE U6492 ( .I1(B[23]), .I2(n5421), .O(n5425) );
  NAND_GATE U6493 ( .I1(n1389), .I2(A[1]), .O(n5422) );
  NAND_GATE U6494 ( .I1(n14784), .I2(n5422), .O(n5423) );
  NAND_GATE U6495 ( .I1(B[22]), .I2(n5423), .O(n5424) );
  NAND_GATE U6496 ( .I1(n5425), .I2(n5424), .O(n5680) );
  NAND_GATE U6497 ( .I1(n5684), .I2(n5680), .O(n5688) );
  NAND3_GATE U6498 ( .I1(B[21]), .I2(B[22]), .I3(n1196), .O(n5681) );
  INV_GATE U6499 ( .I1(n5681), .O(n5689) );
  NAND_GATE U6500 ( .I1(n5679), .I2(n5682), .O(n5426) );
  NAND_GATE U6501 ( .I1(n5689), .I2(n5426), .O(n5427) );
  NAND_GATE U6502 ( .I1(n5688), .I2(n5427), .O(n5663) );
  NAND_GATE U6503 ( .I1(n5429), .I2(n5428), .O(n5434) );
  NAND3_GATE U6504 ( .I1(n174), .I2(n5430), .I3(n5436), .O(n5433) );
  NAND_GATE U6505 ( .I1(n5431), .I2(n1199), .O(n5432) );
  NAND3_GATE U6506 ( .I1(n5434), .I2(n5433), .I3(n5432), .O(n5438) );
  OR_GATE U6507 ( .I1(n5436), .I2(n5435), .O(n5437) );
  NAND_GATE U6508 ( .I1(n5438), .I2(n5437), .O(n5664) );
  NAND_GATE U6509 ( .I1(n5663), .I2(n5664), .O(n5440) );
  NAND_GATE U6510 ( .I1(B[21]), .I2(A[3]), .O(n5668) );
  INV_GATE U6511 ( .I1(n5668), .O(n5659) );
  NAND_GATE U6512 ( .I1(n5659), .I2(n5664), .O(n5439) );
  NAND_GATE U6513 ( .I1(n5659), .I2(n5663), .O(n5660) );
  NAND3_GATE U6514 ( .I1(n5440), .I2(n5439), .I3(n5660), .O(n5700) );
  NAND_GATE U6515 ( .I1(n5694), .I2(n5696), .O(n5441) );
  NAND_GATE U6516 ( .I1(n5723), .I2(n5710), .O(n5705) );
  NAND3_GATE U6517 ( .I1(n5443), .I2(n614), .I3(n5442), .O(n5721) );
  NAND_GATE U6518 ( .I1(n614), .I2(n5445), .O(n5708) );
  NAND_GATE U6519 ( .I1(n714), .I2(n5444), .O(n5445) );
  NAND_GATE U6520 ( .I1(n5446), .I2(n5445), .O(n5718) );
  NAND_GATE U6521 ( .I1(n5708), .I2(n5447), .O(n5707) );
  NAND_GATE U6522 ( .I1(n5721), .I2(n5707), .O(n5448) );
  NAND_GATE U6523 ( .I1(n5710), .I2(n5448), .O(n5449) );
  NAND_GATE U6524 ( .I1(n5723), .I2(n5448), .O(n5713) );
  NAND_GATE U6525 ( .I1(B[21]), .I2(A[6]), .O(n6306) );
  INV_GATE U6526 ( .I1(n5467), .O(n5463) );
  NAND4_GATE U6527 ( .I1(n5463), .I2(n5451), .I3(n5450), .I4(n5465), .O(n5473)
         );
  NAND_GATE U6528 ( .I1(n5453), .I2(n5452), .O(n5454) );
  NAND_GATE U6529 ( .I1(n5455), .I2(n5454), .O(n5456) );
  NAND_GATE U6530 ( .I1(n5456), .I2(n5451), .O(n5460) );
  INV_GATE U6531 ( .I1(n5457), .O(n5459) );
  NAND3_GATE U6532 ( .I1(n5460), .I2(n5459), .I3(n5458), .O(n5472) );
  NAND3_GATE U6533 ( .I1(n5464), .I2(n5463), .I3(n5465), .O(n5469) );
  NAND_GATE U6534 ( .I1(n5465), .I2(n5464), .O(n5466) );
  NAND_GATE U6535 ( .I1(n5467), .I2(n5466), .O(n5468) );
  NAND3_GATE U6536 ( .I1(n5470), .I2(n5469), .I3(n5468), .O(n5471) );
  NAND3_GATE U6537 ( .I1(n5473), .I2(n5472), .I3(n5471), .O(n5736) );
  NAND_GATE U6538 ( .I1(n6306), .I2(n5736), .O(n5474) );
  NAND_GATE U6539 ( .I1(n5735), .I2(n5474), .O(n5476) );
  INV_GATE U6540 ( .I1(n6306), .O(n5733) );
  INV_GATE U6541 ( .I1(n5736), .O(n5734) );
  NAND_GATE U6542 ( .I1(n5733), .I2(n5734), .O(n5475) );
  NAND_GATE U6543 ( .I1(n5476), .I2(n5475), .O(n5756) );
  INV_GATE U6544 ( .I1(n5480), .O(n5477) );
  NAND_GATE U6545 ( .I1(n5477), .I2(n5482), .O(n5754) );
  NAND3_GATE U6546 ( .I1(n5743), .I2(n5478), .I3(n1157), .O(n5479) );
  NAND_GATE U6547 ( .I1(n5480), .I2(n5479), .O(n5481) );
  NAND_GATE U6548 ( .I1(n5754), .I2(n5481), .O(n5747) );
  INV_GATE U6549 ( .I1(n5483), .O(n5742) );
  NAND_GATE U6550 ( .I1(n5742), .I2(n5741), .O(n5485) );
  NAND_GATE U6551 ( .I1(n5483), .I2(n5482), .O(n5484) );
  NAND_GATE U6552 ( .I1(n5485), .I2(n5484), .O(n5751) );
  NAND3_GATE U6553 ( .I1(n5756), .I2(n5747), .I3(n5744), .O(n5488) );
  NAND_GATE U6554 ( .I1(B[21]), .I2(A[7]), .O(n5763) );
  INV_GATE U6555 ( .I1(n5763), .O(n5748) );
  NAND3_GATE U6556 ( .I1(n5748), .I2(n5747), .I3(n5744), .O(n5487) );
  NAND_GATE U6557 ( .I1(n5748), .I2(n5756), .O(n5486) );
  NAND3_GATE U6558 ( .I1(n5488), .I2(n5487), .I3(n5486), .O(n5766) );
  NAND4_GATE U6559 ( .I1(n5491), .I2(n5767), .I3(n5490), .I4(n5489), .O(n5494)
         );
  NAND_GATE U6560 ( .I1(n5767), .I2(n5492), .O(n5493) );
  NAND3_GATE U6561 ( .I1(n5766), .I2(n5494), .I3(n5493), .O(n5495) );
  NAND_GATE U6562 ( .I1(n5496), .I2(n5495), .O(n5651) );
  NAND_GATE U6563 ( .I1(n5654), .I2(n5651), .O(n5652) );
  NAND_GATE U6564 ( .I1(n5502), .I2(n5507), .O(n5500) );
  INV_GATE U6565 ( .I1(n5500), .O(n5497) );
  NAND3_GATE U6566 ( .I1(n1238), .I2(n5498), .I3(n5497), .O(n5650) );
  NAND3_GATE U6567 ( .I1(n5498), .I2(n1238), .I3(n5507), .O(n5499) );
  NAND_GATE U6568 ( .I1(n5500), .I2(n5499), .O(n5648) );
  NAND_GATE U6569 ( .I1(n5650), .I2(n5648), .O(n5504) );
  NAND3_GATE U6570 ( .I1(n783), .I2(n5503), .I3(n5505), .O(n5508) );
  NAND_GATE U6571 ( .I1(n5509), .I2(n5508), .O(n5647) );
  NAND3_GATE U6572 ( .I1(n5504), .I2(n1162), .I3(n5651), .O(n5511) );
  NAND_GATE U6573 ( .I1(n783), .I2(n5505), .O(n5506) );
  NAND3_GATE U6574 ( .I1(n5507), .I2(n5506), .I3(n5650), .O(n5656) );
  NAND3_GATE U6575 ( .I1(n5654), .I2(n5656), .I3(n1162), .O(n5510) );
  NAND3_GATE U6576 ( .I1(n5652), .I2(n5511), .I3(n5510), .O(n5793) );
  NAND_GATE U6577 ( .I1(B[21]), .I2(A[10]), .O(n5791) );
  NAND_GATE U6578 ( .I1(n5513), .I2(n5512), .O(n5514) );
  NAND_GATE U6579 ( .I1(n5515), .I2(n5514), .O(n5517) );
  NAND3_GATE U6580 ( .I1(n5517), .I2(n1363), .I3(n5516), .O(n5520) );
  NAND4_GATE U6581 ( .I1(n5518), .I2(n5524), .I3(n5525), .I4(n5523), .O(n5519)
         );
  AND_GATE U6582 ( .I1(n5520), .I2(n5519), .O(n6431) );
  NAND_GATE U6583 ( .I1(n5524), .I2(n5523), .O(n5521) );
  NAND_GATE U6584 ( .I1(n5522), .I2(n5521), .O(n5527) );
  NAND3_GATE U6585 ( .I1(n5525), .I2(n5524), .I3(n5523), .O(n5526) );
  NAND3_GATE U6586 ( .I1(n5528), .I2(n5527), .I3(n5526), .O(n6430) );
  NAND_GATE U6587 ( .I1(n5791), .I2(n5792), .O(n5529) );
  NAND_GATE U6588 ( .I1(n5793), .I2(n5529), .O(n5531) );
  INV_GATE U6589 ( .I1(n5791), .O(n6429) );
  NAND_GATE U6590 ( .I1(n6429), .I2(n817), .O(n5530) );
  NAND_GATE U6591 ( .I1(n5531), .I2(n5530), .O(n5641) );
  NAND_GATE U6592 ( .I1(n5638), .I2(n5641), .O(n5636) );
  NAND_GATE U6593 ( .I1(n1244), .I2(n5534), .O(n5536) );
  NAND3_GATE U6594 ( .I1(n5532), .I2(n5537), .I3(n5533), .O(n5542) );
  NAND3_GATE U6595 ( .I1(n5537), .I2(n5536), .I3(n5542), .O(n5637) );
  NAND3_GATE U6596 ( .I1(n5535), .I2(n5533), .I3(n5532), .O(n5538) );
  NAND3_GATE U6597 ( .I1(n5535), .I2(n5534), .I3(n1244), .O(n5539) );
  NAND3_GATE U6598 ( .I1(n5638), .I2(n5637), .I3(n1141), .O(n5544) );
  NAND_GATE U6599 ( .I1(n5537), .I2(n5536), .O(n5540) );
  NAND3_GATE U6600 ( .I1(n5540), .I2(n5539), .I3(n5538), .O(n5541) );
  NAND_GATE U6601 ( .I1(n5542), .I2(n5541), .O(n5642) );
  NAND_GATE U6602 ( .I1(n5641), .I2(n5642), .O(n5543) );
  NAND3_GATE U6603 ( .I1(n5636), .I2(n5544), .I3(n5543), .O(n6471) );
  NAND3_GATE U6604 ( .I1(n5546), .I2(n5545), .I3(n6471), .O(n5547) );
  NAND_GATE U6605 ( .I1(n5548), .I2(n5547), .O(n5809) );
  NAND_GATE U6606 ( .I1(n5550), .I2(n5549), .O(n5551) );
  NAND_GATE U6607 ( .I1(n6280), .I2(n5551), .O(n5556) );
  NAND4_GATE U6608 ( .I1(n5554), .I2(n5553), .I3(n6280), .I4(n5552), .O(n5555)
         );
  NAND3_GATE U6609 ( .I1(n5809), .I2(n5556), .I3(n5555), .O(n5557) );
  NAND_GATE U6610 ( .I1(n5558), .I2(n5557), .O(n5817) );
  NAND_GATE U6611 ( .I1(n5821), .I2(n5819), .O(n5559) );
  NAND_GATE U6612 ( .I1(n5817), .I2(n5559), .O(n5560) );
  NAND_GATE U6613 ( .I1(n5814), .I2(n5560), .O(n5633) );
  NAND_GATE U6614 ( .I1(n6254), .I2(n5631), .O(n5561) );
  NAND_GATE U6615 ( .I1(n5633), .I2(n5561), .O(n5562) );
  NAND_GATE U6616 ( .I1(n5834), .I2(n5831), .O(n5564) );
  NAND_GATE U6617 ( .I1(n5846), .I2(n6226), .O(n5565) );
  NAND_GATE U6618 ( .I1(n779), .I2(n5565), .O(n5566) );
  NAND_GATE U6619 ( .I1(n5844), .I2(n5566), .O(n5857) );
  NAND_GATE U6620 ( .I1(n5568), .I2(n5567), .O(n5569) );
  NAND_GATE U6621 ( .I1(n5864), .I2(n5569), .O(n5574) );
  NAND4_GATE U6622 ( .I1(n5572), .I2(n5571), .I3(n5570), .I4(n5864), .O(n5573)
         );
  NAND3_GATE U6623 ( .I1(n5857), .I2(n5574), .I3(n5573), .O(n5575) );
  NAND_GATE U6624 ( .I1(n5856), .I2(n5575), .O(n5879) );
  NAND_GATE U6625 ( .I1(n5876), .I2(n6212), .O(n5576) );
  NAND_GATE U6626 ( .I1(n5879), .I2(n5576), .O(n5577) );
  NAND_GATE U6627 ( .I1(n5878), .I2(n5577), .O(n5626) );
  NAND_GATE U6628 ( .I1(n5622), .I2(n5888), .O(n5578) );
  NAND_GATE U6629 ( .I1(n5626), .I2(n5578), .O(n5579) );
  NAND_GATE U6630 ( .I1(n5625), .I2(n5579), .O(n5900) );
  NAND_GATE U6631 ( .I1(n5896), .I2(n5905), .O(n5580) );
  NAND_GATE U6632 ( .I1(n5900), .I2(n5580), .O(n5581) );
  NAND_GATE U6633 ( .I1(n5899), .I2(n5581), .O(n5912) );
  NAND_GATE U6634 ( .I1(n5915), .I2(n5912), .O(n5916) );
  OR_GATE U6635 ( .I1(n5582), .I2(n5589), .O(n5585) );
  OR_GATE U6636 ( .I1(n5587), .I2(n5583), .O(n5584) );
  AND_GATE U6637 ( .I1(n5585), .I2(n5584), .O(n5594) );
  INV_GATE U6638 ( .I1(n5589), .O(n5586) );
  NAND_GATE U6639 ( .I1(n5586), .I2(n5587), .O(n5592) );
  INV_GATE U6640 ( .I1(n5587), .O(n5588) );
  NAND_GATE U6641 ( .I1(n5589), .I2(n5588), .O(n5591) );
  NAND3_GATE U6642 ( .I1(n5592), .I2(n5591), .I3(n5590), .O(n5593) );
  NAND_GATE U6643 ( .I1(n5594), .I2(n5593), .O(n5911) );
  INV_GATE U6644 ( .I1(n5911), .O(n5917) );
  NAND_GATE U6645 ( .I1(n5923), .I2(n798), .O(n5595) );
  NAND_GATE U6646 ( .I1(n5917), .I2(n5595), .O(n5596) );
  NAND_GATE U6647 ( .I1(n5916), .I2(n5596), .O(n5934) );
  NAND_GATE U6648 ( .I1(n5928), .I2(n5940), .O(n5597) );
  NAND_GATE U6649 ( .I1(n5934), .I2(n5597), .O(n5598) );
  NAND_GATE U6650 ( .I1(n5933), .I2(n5598), .O(n5951) );
  NAND_GATE U6651 ( .I1(n5945), .I2(n5956), .O(n5599) );
  NAND_GATE U6652 ( .I1(n5951), .I2(n5599), .O(n5600) );
  NAND_GATE U6653 ( .I1(n5950), .I2(n5600), .O(n5968) );
  NAND_GATE U6654 ( .I1(n5962), .I2(n5973), .O(n5601) );
  NAND_GATE U6655 ( .I1(n5968), .I2(n5601), .O(n5602) );
  NAND_GATE U6656 ( .I1(n5967), .I2(n5602), .O(n5985) );
  NAND_GATE U6657 ( .I1(n5979), .I2(n5990), .O(n5603) );
  NAND_GATE U6658 ( .I1(n5985), .I2(n5603), .O(n5604) );
  NAND_GATE U6659 ( .I1(n5984), .I2(n5604), .O(n6002) );
  NAND_GATE U6660 ( .I1(n5996), .I2(n6007), .O(n5605) );
  NAND_GATE U6661 ( .I1(n6002), .I2(n5605), .O(n5606) );
  NAND_GATE U6662 ( .I1(n6001), .I2(n5606), .O(n6016) );
  NAND_GATE U6663 ( .I1(n6014), .I2(n6108), .O(n5607) );
  NAND_GATE U6664 ( .I1(n6016), .I2(n5607), .O(n5608) );
  NAND_GATE U6665 ( .I1(n6013), .I2(n5608), .O(n6029) );
  NAND_GATE U6666 ( .I1(n6027), .I2(n6034), .O(n5609) );
  NAND_GATE U6667 ( .I1(n6029), .I2(n5609), .O(n5610) );
  NAND_GATE U6668 ( .I1(n6024), .I2(n5610), .O(n6046) );
  NAND_GATE U6669 ( .I1(n6044), .I2(n6051), .O(n5611) );
  NAND_GATE U6670 ( .I1(n6046), .I2(n5611), .O(n5612) );
  NAND_GATE U6671 ( .I1(n6041), .I2(n5612), .O(n6063) );
  NAND_GATE U6672 ( .I1(n6061), .I2(n6068), .O(n5613) );
  NAND_GATE U6673 ( .I1(n6063), .I2(n5613), .O(n5614) );
  NAND_GATE U6674 ( .I1(n6058), .I2(n5614), .O(n5616) );
  NAND_GATE U6675 ( .I1(n5615), .I2(n5616), .O(n15319) );
  INV_GATE U6676 ( .I1(n5616), .O(n5617) );
  NAND_GATE U6677 ( .I1(n5618), .I2(n5617), .O(n5619) );
  AND_GATE U6678 ( .I1(n15319), .I2(n5619), .O(\A1[51] ) );
  NAND_GATE U6679 ( .I1(B[20]), .I2(A[31]), .O(n6083) );
  INV_GATE U6680 ( .I1(n6083), .O(n6056) );
  NAND_GATE U6681 ( .I1(B[20]), .I2(A[30]), .O(n6094) );
  INV_GATE U6682 ( .I1(n6094), .O(n6039) );
  NAND_GATE U6683 ( .I1(B[20]), .I2(A[29]), .O(n6112) );
  INV_GATE U6684 ( .I1(n6112), .O(n6022) );
  NAND_GATE U6685 ( .I1(B[20]), .I2(A[28]), .O(n6118) );
  INV_GATE U6686 ( .I1(n6118), .O(n6004) );
  NAND_GATE U6687 ( .I1(B[20]), .I2(A[27]), .O(n6135) );
  INV_GATE U6688 ( .I1(n6135), .O(n5987) );
  NAND_GATE U6689 ( .I1(B[20]), .I2(A[26]), .O(n6146) );
  INV_GATE U6690 ( .I1(n6146), .O(n5970) );
  NAND_GATE U6691 ( .I1(B[20]), .I2(A[25]), .O(n6157) );
  INV_GATE U6692 ( .I1(n6157), .O(n5953) );
  NAND_GATE U6693 ( .I1(B[20]), .I2(A[24]), .O(n6168) );
  INV_GATE U6694 ( .I1(n6168), .O(n5936) );
  NAND_GATE U6695 ( .I1(B[20]), .I2(A[23]), .O(n6179) );
  INV_GATE U6696 ( .I1(n6179), .O(n5919) );
  NAND_GATE U6697 ( .I1(B[20]), .I2(A[22]), .O(n6190) );
  INV_GATE U6698 ( .I1(n6190), .O(n5902) );
  NAND_GATE U6699 ( .I1(n583), .I2(n5626), .O(n5620) );
  INV_GATE U6700 ( .I1(n5626), .O(n5621) );
  NAND_GATE U6701 ( .I1(n5620), .I2(n5623), .O(n5887) );
  NAND_GATE U6702 ( .I1(n5622), .I2(n5621), .O(n5623) );
  NAND_GATE U6703 ( .I1(n5624), .I2(n5623), .O(n5890) );
  INV_GATE U6704 ( .I1(n5890), .O(n5627) );
  NAND_GATE U6705 ( .I1(n5627), .I2(n5892), .O(n5628) );
  NAND_GATE U6706 ( .I1(B[20]), .I2(A[21]), .O(n6201) );
  INV_GATE U6707 ( .I1(n6201), .O(n5886) );
  NAND3_GATE U6708 ( .I1(n5889), .I2(n5628), .I3(n5886), .O(n6196) );
  NAND_GATE U6709 ( .I1(B[20]), .I2(A[20]), .O(n6216) );
  INV_GATE U6710 ( .I1(n6216), .O(n5880) );
  NAND_GATE U6711 ( .I1(B[20]), .I2(A[17]), .O(n6241) );
  INV_GATE U6712 ( .I1(n6241), .O(n5842) );
  NAND_GATE U6713 ( .I1(B[20]), .I2(A[16]), .O(n6259) );
  INV_GATE U6714 ( .I1(n6259), .O(n5829) );
  NAND_GATE U6715 ( .I1(n709), .I2(n5633), .O(n5629) );
  INV_GATE U6716 ( .I1(n5633), .O(n5630) );
  NAND_GATE U6717 ( .I1(n5629), .I2(n5632), .O(n6253) );
  NAND_GATE U6718 ( .I1(n5631), .I2(n5630), .O(n5632) );
  NAND_GATE U6719 ( .I1(n5634), .I2(n5632), .O(n6251) );
  NAND_GATE U6720 ( .I1(n6257), .I2(n6251), .O(n5635) );
  NAND3_GATE U6721 ( .I1(n5634), .I2(n5633), .I3(n709), .O(n6252) );
  NAND_GATE U6722 ( .I1(n5635), .I2(n6252), .O(n6262) );
  NAND_GATE U6723 ( .I1(B[20]), .I2(A[15]), .O(n6269) );
  INV_GATE U6724 ( .I1(n6269), .O(n5827) );
  NAND_GATE U6725 ( .I1(B[20]), .I2(A[14]), .O(n6285) );
  INV_GATE U6726 ( .I1(n6285), .O(n5812) );
  NAND_GATE U6727 ( .I1(B[20]), .I2(A[13]), .O(n6482) );
  INV_GATE U6728 ( .I1(n6482), .O(n6470) );
  NAND_GATE U6729 ( .I1(B[20]), .I2(A[12]), .O(n6456) );
  INV_GATE U6730 ( .I1(n6456), .O(n6457) );
  OR_GATE U6731 ( .I1(n5642), .I2(n5636), .O(n5640) );
  NAND4_GATE U6732 ( .I1(n5638), .I2(n5637), .I3(n1141), .I4(n811), .O(n5639)
         );
  NAND_GATE U6733 ( .I1(n5640), .I2(n5639), .O(n5646) );
  INV_GATE U6734 ( .I1(n5646), .O(n6459) );
  NAND_GATE U6735 ( .I1(n5641), .I2(n1228), .O(n5643) );
  NAND_GATE U6736 ( .I1(n811), .I2(n5642), .O(n5644) );
  NAND3_GATE U6737 ( .I1(n5643), .I2(n5644), .I3(n5645), .O(n6458) );
  NAND_GATE U6738 ( .I1(n6457), .I2(n1241), .O(n5801) );
  NAND4_GATE U6739 ( .I1(n5645), .I2(n6456), .I3(n5644), .I4(n5643), .O(n5799)
         );
  NAND_GATE U6740 ( .I1(n6456), .I2(n5646), .O(n5798) );
  NAND_GATE U6741 ( .I1(B[20]), .I2(A[11]), .O(n6445) );
  INV_GATE U6742 ( .I1(n6445), .O(n6428) );
  NAND_GATE U6743 ( .I1(B[20]), .I2(A[10]), .O(n6558) );
  INV_GATE U6744 ( .I1(n5651), .O(n5655) );
  OR_GATE U6745 ( .I1(n5648), .I2(n5647), .O(n5649) );
  NAND_GATE U6746 ( .I1(n5650), .I2(n5649), .O(n5653) );
  NAND_GATE U6747 ( .I1(n5655), .I2(n5653), .O(n5786) );
  NAND4_GATE U6748 ( .I1(n5785), .I2(n6558), .I3(n5786), .I4(n5784), .O(n5783)
         );
  OR_GATE U6749 ( .I1(n5653), .I2(n5652), .O(n5658) );
  NAND4_GATE U6750 ( .I1(n5656), .I2(n5655), .I3(n5654), .I4(n1162), .O(n5657)
         );
  NAND_GATE U6751 ( .I1(n5658), .I2(n5657), .O(n5787) );
  NAND_GATE U6752 ( .I1(n6558), .I2(n5787), .O(n5782) );
  NAND_GATE U6753 ( .I1(B[20]), .I2(A[9]), .O(n6414) );
  INV_GATE U6754 ( .I1(n6414), .O(n6407) );
  NAND_GATE U6755 ( .I1(B[20]), .I2(A[7]), .O(n6314) );
  INV_GATE U6756 ( .I1(n6314), .O(n6301) );
  NAND_GATE U6757 ( .I1(B[20]), .I2(A[5]), .O(n6375) );
  INV_GATE U6758 ( .I1(n6375), .O(n6366) );
  NAND_GATE U6759 ( .I1(B[20]), .I2(A[4]), .O(n6319) );
  INV_GATE U6760 ( .I1(n6319), .O(n6316) );
  INV_GATE U6761 ( .I1(n5663), .O(n5665) );
  NAND3_GATE U6762 ( .I1(n5665), .I2(n5659), .I3(n5664), .O(n5662) );
  OR_GATE U6763 ( .I1(n5664), .I2(n5660), .O(n5661) );
  AND_GATE U6764 ( .I1(n5662), .I2(n5661), .O(n5670) );
  NAND_GATE U6765 ( .I1(n5665), .I2(n5664), .O(n5666) );
  NAND3_GATE U6766 ( .I1(n5668), .I2(n5667), .I3(n5666), .O(n5669) );
  NAND_GATE U6767 ( .I1(n5670), .I2(n5669), .O(n6318) );
  NAND_GATE U6768 ( .I1(n6316), .I2(n169), .O(n6322) );
  NAND_GATE U6769 ( .I1(B[20]), .I2(A[3]), .O(n6338) );
  INV_GATE U6770 ( .I1(n6338), .O(n5690) );
  NAND_GATE U6771 ( .I1(B[20]), .I2(A[2]), .O(n6355) );
  INV_GATE U6772 ( .I1(n6355), .O(n6350) );
  NAND_GATE U6773 ( .I1(n1387), .I2(A[0]), .O(n5671) );
  NAND_GATE U6774 ( .I1(n14781), .I2(n5671), .O(n5672) );
  NAND_GATE U6775 ( .I1(B[22]), .I2(n5672), .O(n5675) );
  NAND_GATE U6776 ( .I1(n1388), .I2(A[1]), .O(n5673) );
  NAND_GATE U6777 ( .I1(n14784), .I2(n5673), .O(n5674) );
  NAND_GATE U6778 ( .I1(B[21]), .I2(n5674), .O(n5676) );
  NAND_GATE U6779 ( .I1(n5675), .I2(n5676), .O(n6351) );
  NAND_GATE U6780 ( .I1(n6350), .I2(n6351), .O(n6358) );
  NAND3_GATE U6781 ( .I1(B[20]), .I2(B[21]), .I3(n1196), .O(n6349) );
  INV_GATE U6782 ( .I1(n6349), .O(n6359) );
  NAND_GATE U6783 ( .I1(n6355), .I2(n5676), .O(n5677) );
  NAND_GATE U6784 ( .I1(n6359), .I2(n5677), .O(n5678) );
  NAND_GATE U6785 ( .I1(n6358), .I2(n5678), .O(n6333) );
  NAND_GATE U6786 ( .I1(n5690), .I2(n6333), .O(n6328) );
  NAND3_GATE U6787 ( .I1(n5681), .I2(n5682), .I3(n5679), .O(n5687) );
  NAND_GATE U6788 ( .I1(n5680), .I2(n5689), .O(n5686) );
  NAND_GATE U6789 ( .I1(n5682), .I2(n5681), .O(n5683) );
  NAND_GATE U6790 ( .I1(n5684), .I2(n5683), .O(n5685) );
  NAND3_GATE U6791 ( .I1(n5687), .I2(n5686), .I3(n5685), .O(n6331) );
  NAND_GATE U6792 ( .I1(n6331), .I2(n6332), .O(n6334) );
  NAND_GATE U6793 ( .I1(n6333), .I2(n6334), .O(n5691) );
  NAND_GATE U6794 ( .I1(n5690), .I2(n6334), .O(n6327) );
  NAND3_GATE U6795 ( .I1(n6328), .I2(n5691), .I3(n6327), .O(n6323) );
  NAND_GATE U6796 ( .I1(n6319), .I2(n6318), .O(n5692) );
  NAND_GATE U6797 ( .I1(n6323), .I2(n5692), .O(n5693) );
  NAND_GATE U6798 ( .I1(n6322), .I2(n5693), .O(n6370) );
  NAND_GATE U6799 ( .I1(n6366), .I2(n6370), .O(n6367) );
  INV_GATE U6800 ( .I1(n5700), .O(n5695) );
  NAND3_GATE U6801 ( .I1(n5696), .I2(n5695), .I3(n5694), .O(n5698) );
  NAND3_GATE U6802 ( .I1(n5699), .I2(n5698), .I3(n5697), .O(n5702) );
  NAND_GATE U6803 ( .I1(n1351), .I2(n5700), .O(n5701) );
  NAND_GATE U6804 ( .I1(n5702), .I2(n5701), .O(n6371) );
  NAND_GATE U6805 ( .I1(n6370), .I2(n6371), .O(n5704) );
  NAND_GATE U6806 ( .I1(n6366), .I2(n6371), .O(n5703) );
  NAND3_GATE U6807 ( .I1(n6367), .I2(n5704), .I3(n5703), .O(n6588) );
  INV_GATE U6808 ( .I1(n5705), .O(n5706) );
  NAND3_GATE U6809 ( .I1(n5707), .I2(n5721), .I3(n5706), .O(n5730) );
  NAND_GATE U6810 ( .I1(B[20]), .I2(A[6]), .O(n6589) );
  NAND_GATE U6811 ( .I1(n5719), .I2(n5718), .O(n5712) );
  INV_GATE U6812 ( .I1(n5708), .O(n5720) );
  NAND_GATE U6813 ( .I1(n5712), .I2(n5711), .O(n5709) );
  NAND_GATE U6814 ( .I1(n5710), .I2(n5709), .O(n5726) );
  INV_GATE U6815 ( .I1(n5710), .O(n5724) );
  NAND3_GATE U6816 ( .I1(n5712), .I2(n5711), .I3(n5724), .O(n5727) );
  NAND4_GATE U6817 ( .I1(n5725), .I2(n5726), .I3(n6589), .I4(n5727), .O(n5716)
         );
  INV_GATE U6818 ( .I1(n5713), .O(n5714) );
  NAND3_GATE U6819 ( .I1(n5724), .I2(n5714), .I3(n6589), .O(n5715) );
  NAND4_GATE U6820 ( .I1(n6588), .I2(n5717), .I3(n5716), .I4(n5715), .O(n5732)
         );
  NAND_GATE U6821 ( .I1(n5721), .I2(n5720), .O(n5722) );
  NAND4_GATE U6822 ( .I1(n5724), .I2(n5723), .I3(n5712), .I4(n5722), .O(n5729)
         );
  NAND3_GATE U6823 ( .I1(n5727), .I2(n5726), .I3(n5725), .O(n5728) );
  NAND3_GATE U6824 ( .I1(n5730), .I2(n5729), .I3(n5728), .O(n6590) );
  NAND_GATE U6825 ( .I1(n1067), .I2(n1206), .O(n5731) );
  NAND_GATE U6826 ( .I1(n5732), .I2(n5731), .O(n6311) );
  NAND_GATE U6827 ( .I1(n6301), .I2(n6311), .O(n6298) );
  NAND3_GATE U6828 ( .I1(n5735), .I2(n5733), .I3(n5734), .O(n6304) );
  NAND_GATE U6829 ( .I1(n1361), .I2(n5736), .O(n5737) );
  NAND_GATE U6830 ( .I1(n5738), .I2(n5737), .O(n6305) );
  NAND3_GATE U6831 ( .I1(n6311), .I2(n6309), .I3(n6308), .O(n5740) );
  NAND3_GATE U6832 ( .I1(n6301), .I2(n6309), .I3(n6308), .O(n5739) );
  NAND3_GATE U6833 ( .I1(n6298), .I2(n5740), .I3(n5739), .O(n6391) );
  NAND_GATE U6834 ( .I1(B[20]), .I2(A[8]), .O(n6390) );
  AND3_GATE U6835 ( .I1(n5754), .I2(n5756), .I3(n5748), .O(n5746) );
  NAND_GATE U6836 ( .I1(n5743), .I2(n5485), .O(n5753) );
  NAND_GATE U6837 ( .I1(n5752), .I2(n5751), .O(n5744) );
  NAND_GATE U6838 ( .I1(n5753), .I2(n5744), .O(n5745) );
  NAND_GATE U6839 ( .I1(n5746), .I2(n5745), .O(n5750) );
  INV_GATE U6840 ( .I1(n5756), .O(n5758) );
  NAND4_GATE U6841 ( .I1(n5748), .I2(n5747), .I3(n5758), .I4(n5744), .O(n5749)
         );
  NAND_GATE U6842 ( .I1(n5744), .I2(n5757), .O(n5755) );
  NAND_GATE U6843 ( .I1(n5756), .I2(n5755), .O(n5762) );
  NAND3_GATE U6844 ( .I1(n5758), .I2(n5757), .I3(n5744), .O(n5761) );
  NAND4_GATE U6845 ( .I1(n5763), .I2(n5762), .I3(n6390), .I4(n5761), .O(n5759)
         );
  NAND3_GATE U6846 ( .I1(n6391), .I2(n5760), .I3(n5759), .O(n5765) );
  INV_GATE U6847 ( .I1(n6390), .O(n6399) );
  NAND3_GATE U6848 ( .I1(n5763), .I2(n5762), .I3(n5761), .O(n6392) );
  NAND_GATE U6849 ( .I1(n794), .I2(n6392), .O(n6398) );
  NAND_GATE U6850 ( .I1(n5765), .I2(n5764), .O(n6409) );
  NAND_GATE U6851 ( .I1(n6407), .I2(n6409), .O(n6408) );
  NAND_GATE U6852 ( .I1(n5777), .I2(n5766), .O(n5769) );
  NAND3_GATE U6853 ( .I1(n5777), .I2(n5772), .I3(n5771), .O(n5768) );
  INV_GATE U6854 ( .I1(n5766), .O(n5774) );
  NAND3_GATE U6855 ( .I1(n5767), .I2(n5774), .I3(n764), .O(n5778) );
  NAND4_GATE U6856 ( .I1(n5769), .I2(n5768), .I3(n5779), .I4(n5778), .O(n5773)
         );
  INV_GATE U6857 ( .I1(n5769), .O(n5770) );
  NAND3_GATE U6858 ( .I1(n5772), .I2(n5771), .I3(n5770), .O(n5775) );
  NAND_GATE U6859 ( .I1(n5773), .I2(n5775), .O(n6410) );
  NAND_GATE U6860 ( .I1(n6409), .I2(n6410), .O(n5781) );
  NAND_GATE U6861 ( .I1(n764), .I2(n5774), .O(n5776) );
  NAND3_GATE U6862 ( .I1(n5777), .I2(n5776), .I3(n5775), .O(n6406) );
  NAND3_GATE U6863 ( .I1(n6407), .I2(n6406), .I3(n1161), .O(n5780) );
  NAND3_GATE U6864 ( .I1(n6408), .I2(n5781), .I3(n5780), .O(n6423) );
  NAND3_GATE U6865 ( .I1(n5783), .I2(n5782), .I3(n6423), .O(n5790) );
  INV_GATE U6866 ( .I1(n6558), .O(n6422) );
  AND3_GATE U6867 ( .I1(n5786), .I2(n5785), .I3(n5784), .O(n5788) );
  NAND_GATE U6868 ( .I1(n6422), .I2(n784), .O(n5789) );
  NAND_GATE U6869 ( .I1(n5790), .I2(n5789), .O(n6442) );
  NAND_GATE U6870 ( .I1(n6428), .I2(n6442), .O(n6438) );
  NAND3_GATE U6871 ( .I1(n855), .I2(n5791), .I3(n5792), .O(n6433) );
  NAND_GATE U6872 ( .I1(n855), .I2(n5792), .O(n5795) );
  NAND_GATE U6873 ( .I1(n5793), .I2(n6429), .O(n6435) );
  INV_GATE U6874 ( .I1(n6435), .O(n5794) );
  NAND_GATE U6875 ( .I1(n817), .I2(n5794), .O(n6437) );
  NAND3_GATE U6876 ( .I1(n6429), .I2(n5795), .I3(n6437), .O(n6427) );
  NAND3_GATE U6877 ( .I1(n6442), .I2(n1165), .I3(n6427), .O(n5797) );
  NAND3_GATE U6878 ( .I1(n6428), .I2(n6427), .I3(n1165), .O(n5796) );
  NAND3_GATE U6879 ( .I1(n6438), .I2(n5797), .I3(n5796), .O(n6454) );
  NAND3_GATE U6880 ( .I1(n5799), .I2(n5798), .I3(n6454), .O(n5800) );
  NAND_GATE U6881 ( .I1(n5801), .I2(n5800), .O(n6479) );
  NAND_GATE U6882 ( .I1(n6470), .I2(n6479), .O(n6476) );
  NAND_GATE U6883 ( .I1(n6473), .I2(n595), .O(n5802) );
  NAND_GATE U6884 ( .I1(n5803), .I2(n5802), .O(n6474) );
  NAND_GATE U6885 ( .I1(n619), .I2(n6471), .O(n5804) );
  NAND_GATE U6886 ( .I1(n5804), .I2(n5802), .O(n5805) );
  NAND_GATE U6887 ( .I1(n6472), .I2(n5805), .O(n6468) );
  NAND3_GATE U6888 ( .I1(n6469), .I2(n6468), .I3(n6470), .O(n5806) );
  AND_GATE U6889 ( .I1(n6476), .I2(n5806), .O(n6282) );
  NAND3_GATE U6890 ( .I1(n6479), .I2(n6469), .I3(n6468), .O(n6281) );
  NAND_GATE U6891 ( .I1(n6282), .I2(n6281), .O(n6288) );
  NAND_GATE U6892 ( .I1(n5808), .I2(n5807), .O(n6291) );
  NAND3_GATE U6893 ( .I1(n5808), .I2(n5809), .I3(n5810), .O(n6293) );
  NAND_GATE U6894 ( .I1(n5810), .I2(n5809), .O(n5811) );
  NAND_GATE U6895 ( .I1(n5811), .I2(n5807), .O(n6279) );
  NAND_GATE U6896 ( .I1(n6280), .I2(n6279), .O(n6290) );
  NAND3_GATE U6897 ( .I1(n5812), .I2(n6283), .I3(n6290), .O(n6289) );
  NAND3_GATE U6898 ( .I1(n6288), .I2(n6283), .I3(n6290), .O(n5813) );
  NAND3_GATE U6899 ( .I1(n219), .I2(n6289), .I3(n5813), .O(n6272) );
  NAND_GATE U6900 ( .I1(n5827), .I2(n6272), .O(n6274) );
  INV_GATE U6901 ( .I1(n5817), .O(n5820) );
  NAND_GATE U6902 ( .I1(n5821), .I2(n5820), .O(n5815) );
  NAND_GATE U6903 ( .I1(n5816), .I2(n5815), .O(n5824) );
  NAND_GATE U6904 ( .I1(n5818), .I2(n5817), .O(n5823) );
  NAND3_GATE U6905 ( .I1(n5821), .I2(n5820), .I3(n5819), .O(n5822) );
  NAND3_GATE U6906 ( .I1(n5824), .I2(n5823), .I3(n5822), .O(n5825) );
  NAND_GATE U6907 ( .I1(n5826), .I2(n5825), .O(n6275) );
  NAND_GATE U6908 ( .I1(n5827), .I2(n6275), .O(n6273) );
  NAND_GATE U6909 ( .I1(n6272), .I2(n6275), .O(n5828) );
  NAND3_GATE U6910 ( .I1(n6274), .I2(n6273), .I3(n5828), .O(n6265) );
  NAND_GATE U6911 ( .I1(n6262), .I2(n6265), .O(n5830) );
  NAND_GATE U6912 ( .I1(n5829), .I2(n6265), .O(n6263) );
  NAND3_GATE U6913 ( .I1(n6264), .I2(n5830), .I3(n6263), .O(n6244) );
  NAND_GATE U6914 ( .I1(n5842), .I2(n6244), .O(n6246) );
  NAND_GATE U6915 ( .I1(n801), .I2(n5832), .O(n5841) );
  NAND3_GATE U6916 ( .I1(n5831), .I2(n756), .I3(n5834), .O(n5839) );
  NAND_GATE U6917 ( .I1(n5833), .I2(n5832), .O(n5838) );
  NAND_GATE U6918 ( .I1(n5834), .I2(n756), .O(n5835) );
  NAND_GATE U6919 ( .I1(n5836), .I2(n5835), .O(n5837) );
  NAND3_GATE U6920 ( .I1(n5839), .I2(n5838), .I3(n5837), .O(n5840) );
  NAND_GATE U6921 ( .I1(n5841), .I2(n5840), .O(n6247) );
  NAND_GATE U6922 ( .I1(n5842), .I2(n6247), .O(n6245) );
  NAND_GATE U6923 ( .I1(n6244), .I2(n6247), .O(n5843) );
  NAND3_GATE U6924 ( .I1(n6246), .I2(n6245), .I3(n5843), .O(n6230) );
  NAND_GATE U6925 ( .I1(n5845), .I2(n5847), .O(n6222) );
  NAND_GATE U6926 ( .I1(n545), .I2(n779), .O(n5848) );
  NAND_GATE U6927 ( .I1(n5846), .I2(n872), .O(n5847) );
  NAND_GATE U6928 ( .I1(n5848), .I2(n5847), .O(n6225) );
  NAND_GATE U6929 ( .I1(n6222), .I2(n6227), .O(n5849) );
  NAND_GATE U6930 ( .I1(n6224), .I2(n5849), .O(n6232) );
  NAND_GATE U6931 ( .I1(n6230), .I2(n6232), .O(n5862) );
  NAND_GATE U6932 ( .I1(B[20]), .I2(A[19]), .O(n6508) );
  OR_GATE U6933 ( .I1(n5862), .I2(n6508), .O(n5871) );
  INV_GATE U6934 ( .I1(n6508), .O(n6503) );
  NAND_GATE U6935 ( .I1(B[20]), .I2(A[18]), .O(n6237) );
  INV_GATE U6936 ( .I1(n6237), .O(n5850) );
  NAND_GATE U6937 ( .I1(n6230), .I2(n5850), .O(n6233) );
  NAND_GATE U6938 ( .I1(n6232), .I2(n5850), .O(n6221) );
  NAND_GATE U6939 ( .I1(n6233), .I2(n6221), .O(n5861) );
  NAND_GATE U6940 ( .I1(n6503), .I2(n5861), .O(n5870) );
  NAND_GATE U6941 ( .I1(n788), .I2(n5857), .O(n5852) );
  NAND_GATE U6942 ( .I1(n5852), .I2(n5851), .O(n5863) );
  NAND_GATE U6943 ( .I1(n5864), .I2(n5863), .O(n5860) );
  NAND_GATE U6944 ( .I1(n5853), .I2(n541), .O(n5854) );
  NAND_GATE U6945 ( .I1(n5855), .I2(n5854), .O(n5866) );
  INV_GATE U6946 ( .I1(n5866), .O(n5858) );
  NAND_GATE U6947 ( .I1(n5858), .I2(n5868), .O(n5859) );
  NAND3_GATE U6948 ( .I1(n5860), .I2(n5859), .I3(n6503), .O(n6502) );
  NAND_GATE U6949 ( .I1(n5866), .I2(n5865), .O(n5867) );
  NAND_GATE U6950 ( .I1(n6507), .I2(n6506), .O(n5869) );
  NAND_GATE U6951 ( .I1(n5880), .I2(n6215), .O(n6207) );
  NAND_GATE U6952 ( .I1(n5872), .I2(n5879), .O(n5874) );
  INV_GATE U6953 ( .I1(n5879), .O(n5875) );
  NAND_GATE U6954 ( .I1(n5876), .I2(n5875), .O(n5873) );
  NAND_GATE U6955 ( .I1(n5874), .I2(n5873), .O(n6211) );
  NAND_GATE U6956 ( .I1(n6212), .I2(n6211), .O(n5881) );
  NAND_GATE U6957 ( .I1(n5877), .I2(n5873), .O(n5882) );
  NAND3_GATE U6958 ( .I1(n5881), .I2(n6213), .I3(n5880), .O(n6206) );
  NAND_GATE U6959 ( .I1(n5882), .I2(n5881), .O(n5883) );
  NAND_GATE U6960 ( .I1(n5884), .I2(n5883), .O(n6210) );
  NAND_GATE U6961 ( .I1(n6215), .I2(n6210), .O(n5885) );
  NAND3_GATE U6962 ( .I1(n6207), .I2(n6206), .I3(n5885), .O(n6200) );
  NAND_GATE U6963 ( .I1(n5886), .I2(n6200), .O(n6195) );
  NAND_GATE U6964 ( .I1(n5888), .I2(n5887), .O(n5889) );
  NAND_GATE U6965 ( .I1(n5890), .I2(n5889), .O(n5891) );
  NAND_GATE U6966 ( .I1(n5892), .I2(n5891), .O(n6199) );
  NAND_GATE U6967 ( .I1(n6200), .I2(n6199), .O(n5893) );
  NAND3_GATE U6968 ( .I1(n6196), .I2(n6195), .I3(n5893), .O(n6189) );
  NAND_GATE U6969 ( .I1(n5902), .I2(n6189), .O(n6185) );
  NAND_GATE U6970 ( .I1(n564), .I2(n5900), .O(n5894) );
  INV_GATE U6971 ( .I1(n5900), .O(n5895) );
  NAND_GATE U6972 ( .I1(n5894), .I2(n5897), .O(n5904) );
  NAND_GATE U6973 ( .I1(n5896), .I2(n5895), .O(n5897) );
  NAND_GATE U6974 ( .I1(n5898), .I2(n5897), .O(n5907) );
  INV_GATE U6975 ( .I1(n5907), .O(n5901) );
  NAND_GATE U6976 ( .I1(n5901), .I2(n5909), .O(n5903) );
  NAND3_GATE U6977 ( .I1(n5906), .I2(n5903), .I3(n5902), .O(n6184) );
  NAND_GATE U6978 ( .I1(n5905), .I2(n5904), .O(n5906) );
  NAND_GATE U6979 ( .I1(n5907), .I2(n5906), .O(n5908) );
  NAND_GATE U6980 ( .I1(n5909), .I2(n5908), .O(n6188) );
  NAND_GATE U6981 ( .I1(n6189), .I2(n6188), .O(n5910) );
  NAND3_GATE U6982 ( .I1(n6185), .I2(n6184), .I3(n5910), .O(n6178) );
  NAND_GATE U6983 ( .I1(n5919), .I2(n6178), .O(n6174) );
  NAND_GATE U6984 ( .I1(n798), .I2(n5911), .O(n5914) );
  NAND_GATE U6985 ( .I1(n5912), .I2(n5917), .O(n5913) );
  NAND_GATE U6986 ( .I1(n5914), .I2(n5913), .O(n5922) );
  NAND_GATE U6987 ( .I1(n5923), .I2(n5922), .O(n5921) );
  NAND_GATE U6988 ( .I1(n5915), .I2(n5914), .O(n5924) );
  INV_GATE U6989 ( .I1(n5924), .O(n5918) );
  NAND_GATE U6990 ( .I1(n5918), .I2(n5926), .O(n5920) );
  NAND3_GATE U6991 ( .I1(n5921), .I2(n5920), .I3(n5919), .O(n6173) );
  NAND_GATE U6992 ( .I1(n5924), .I2(n5921), .O(n5925) );
  NAND_GATE U6993 ( .I1(n5926), .I2(n5925), .O(n6177) );
  NAND_GATE U6994 ( .I1(n6178), .I2(n6177), .O(n5927) );
  NAND3_GATE U6995 ( .I1(n6174), .I2(n6173), .I3(n5927), .O(n6167) );
  NAND_GATE U6996 ( .I1(n5936), .I2(n6167), .O(n6163) );
  NAND_GATE U6997 ( .I1(n5929), .I2(n5934), .O(n5930) );
  NAND_GATE U6998 ( .I1(n5931), .I2(n5930), .O(n5939) );
  NAND_GATE U6999 ( .I1(n5940), .I2(n5939), .O(n5938) );
  NAND_GATE U7000 ( .I1(n5932), .I2(n5931), .O(n5941) );
  INV_GATE U7001 ( .I1(n5933), .O(n5935) );
  NAND_GATE U7002 ( .I1(n5935), .I2(n5934), .O(n5943) );
  NAND3_GATE U7003 ( .I1(n5938), .I2(n5937), .I3(n5936), .O(n6162) );
  NAND_GATE U7004 ( .I1(n5941), .I2(n5938), .O(n5942) );
  NAND_GATE U7005 ( .I1(n5943), .I2(n5942), .O(n6166) );
  NAND_GATE U7006 ( .I1(n6167), .I2(n6166), .O(n5944) );
  NAND3_GATE U7007 ( .I1(n6163), .I2(n6162), .I3(n5944), .O(n6156) );
  NAND_GATE U7008 ( .I1(n5953), .I2(n6156), .O(n6152) );
  NAND_GATE U7009 ( .I1(n5946), .I2(n5951), .O(n5947) );
  NAND_GATE U7010 ( .I1(n5948), .I2(n5947), .O(n5955) );
  NAND_GATE U7011 ( .I1(n5949), .I2(n5948), .O(n5958) );
  INV_GATE U7012 ( .I1(n5950), .O(n5952) );
  NAND_GATE U7013 ( .I1(n5952), .I2(n5951), .O(n5960) );
  NAND3_GATE U7014 ( .I1(n5957), .I2(n5954), .I3(n5953), .O(n6151) );
  NAND_GATE U7015 ( .I1(n5956), .I2(n5955), .O(n5957) );
  NAND_GATE U7016 ( .I1(n5958), .I2(n5957), .O(n5959) );
  NAND_GATE U7017 ( .I1(n5960), .I2(n5959), .O(n6155) );
  NAND_GATE U7018 ( .I1(n6156), .I2(n6155), .O(n5961) );
  NAND3_GATE U7019 ( .I1(n6152), .I2(n6151), .I3(n5961), .O(n6145) );
  NAND_GATE U7020 ( .I1(n5970), .I2(n6145), .O(n6141) );
  NAND_GATE U7021 ( .I1(n5963), .I2(n5968), .O(n5964) );
  NAND_GATE U7022 ( .I1(n5965), .I2(n5964), .O(n5972) );
  NAND_GATE U7023 ( .I1(n5966), .I2(n5965), .O(n5975) );
  INV_GATE U7024 ( .I1(n5967), .O(n5969) );
  NAND_GATE U7025 ( .I1(n5969), .I2(n5968), .O(n5977) );
  NAND3_GATE U7026 ( .I1(n5974), .I2(n5971), .I3(n5970), .O(n6140) );
  NAND_GATE U7027 ( .I1(n5973), .I2(n5972), .O(n5974) );
  NAND_GATE U7028 ( .I1(n5975), .I2(n5974), .O(n5976) );
  NAND_GATE U7029 ( .I1(n5977), .I2(n5976), .O(n6144) );
  NAND_GATE U7030 ( .I1(n6145), .I2(n6144), .O(n5978) );
  NAND3_GATE U7031 ( .I1(n6141), .I2(n6140), .I3(n5978), .O(n6134) );
  NAND_GATE U7032 ( .I1(n5987), .I2(n6134), .O(n6130) );
  NAND_GATE U7033 ( .I1(n5980), .I2(n5985), .O(n5981) );
  NAND_GATE U7034 ( .I1(n5982), .I2(n5981), .O(n5989) );
  NAND_GATE U7035 ( .I1(n5983), .I2(n5982), .O(n5992) );
  INV_GATE U7036 ( .I1(n5984), .O(n5986) );
  NAND_GATE U7037 ( .I1(n5986), .I2(n5985), .O(n5994) );
  NAND3_GATE U7038 ( .I1(n5991), .I2(n5988), .I3(n5987), .O(n6129) );
  NAND_GATE U7039 ( .I1(n5990), .I2(n5989), .O(n5991) );
  NAND_GATE U7040 ( .I1(n5992), .I2(n5991), .O(n5993) );
  NAND_GATE U7041 ( .I1(n5994), .I2(n5993), .O(n6133) );
  NAND_GATE U7042 ( .I1(n6134), .I2(n6133), .O(n5995) );
  NAND3_GATE U7043 ( .I1(n6130), .I2(n6129), .I3(n5995), .O(n6117) );
  NAND_GATE U7044 ( .I1(n6004), .I2(n6117), .O(n6121) );
  NAND_GATE U7045 ( .I1(n5997), .I2(n6002), .O(n5998) );
  NAND_GATE U7046 ( .I1(n5999), .I2(n5998), .O(n6006) );
  NAND_GATE U7047 ( .I1(n6000), .I2(n5999), .O(n6009) );
  INV_GATE U7048 ( .I1(n6009), .O(n6003) );
  NAND_GATE U7049 ( .I1(n6003), .I2(n6011), .O(n6005) );
  NAND3_GATE U7050 ( .I1(n6008), .I2(n6005), .I3(n6004), .O(n6125) );
  NAND_GATE U7051 ( .I1(n6007), .I2(n6006), .O(n6008) );
  NAND_GATE U7052 ( .I1(n6009), .I2(n6008), .O(n6010) );
  NAND_GATE U7053 ( .I1(n6011), .I2(n6010), .O(n6122) );
  NAND_GATE U7054 ( .I1(n6117), .I2(n6122), .O(n6012) );
  NAND3_GATE U7055 ( .I1(n6121), .I2(n6125), .I3(n6012), .O(n6111) );
  NAND_GATE U7056 ( .I1(n6022), .I2(n6111), .O(n6099) );
  NAND_GATE U7057 ( .I1(n6015), .I2(n6019), .O(n6104) );
  NAND_GATE U7058 ( .I1(n6017), .I2(n6016), .O(n6018) );
  NAND_GATE U7059 ( .I1(n6019), .I2(n6018), .O(n6107) );
  NAND_GATE U7060 ( .I1(n6108), .I2(n6107), .O(n6020) );
  NAND_GATE U7061 ( .I1(n6104), .I2(n6020), .O(n6021) );
  NAND_GATE U7062 ( .I1(n6106), .I2(n6021), .O(n6102) );
  NAND_GATE U7063 ( .I1(n6022), .I2(n6102), .O(n6098) );
  NAND_GATE U7064 ( .I1(n6111), .I2(n6102), .O(n6023) );
  NAND3_GATE U7065 ( .I1(n6099), .I2(n6098), .I3(n6023), .O(n6093) );
  NAND_GATE U7066 ( .I1(n6039), .I2(n6093), .O(n6089) );
  INV_GATE U7067 ( .I1(n6024), .O(n6025) );
  NAND_GATE U7068 ( .I1(n6025), .I2(n6029), .O(n6038) );
  INV_GATE U7069 ( .I1(n6029), .O(n6026) );
  NAND_GATE U7070 ( .I1(n6027), .I2(n6026), .O(n6032) );
  NAND_GATE U7071 ( .I1(n6028), .I2(n6032), .O(n6036) );
  NAND_GATE U7072 ( .I1(n6030), .I2(n6029), .O(n6031) );
  NAND_GATE U7073 ( .I1(n6032), .I2(n6031), .O(n6033) );
  NAND_GATE U7074 ( .I1(n6034), .I2(n6033), .O(n6035) );
  NAND_GATE U7075 ( .I1(n6036), .I2(n6035), .O(n6037) );
  NAND_GATE U7076 ( .I1(n6038), .I2(n6037), .O(n6092) );
  NAND_GATE U7077 ( .I1(n6039), .I2(n6092), .O(n6088) );
  NAND_GATE U7078 ( .I1(n6093), .I2(n6092), .O(n6040) );
  NAND3_GATE U7079 ( .I1(n6089), .I2(n6088), .I3(n6040), .O(n6082) );
  NAND_GATE U7080 ( .I1(n6056), .I2(n6082), .O(n6078) );
  INV_GATE U7081 ( .I1(n6041), .O(n6042) );
  NAND_GATE U7082 ( .I1(n6042), .I2(n6046), .O(n6055) );
  INV_GATE U7083 ( .I1(n6046), .O(n6043) );
  NAND_GATE U7084 ( .I1(n6044), .I2(n6043), .O(n6049) );
  NAND_GATE U7085 ( .I1(n6045), .I2(n6049), .O(n6053) );
  NAND_GATE U7086 ( .I1(n6047), .I2(n6046), .O(n6048) );
  NAND_GATE U7087 ( .I1(n6049), .I2(n6048), .O(n6050) );
  NAND_GATE U7088 ( .I1(n6051), .I2(n6050), .O(n6052) );
  NAND_GATE U7089 ( .I1(n6053), .I2(n6052), .O(n6054) );
  NAND_GATE U7090 ( .I1(n6055), .I2(n6054), .O(n6081) );
  NAND_GATE U7091 ( .I1(n6056), .I2(n6081), .O(n6077) );
  NAND_GATE U7092 ( .I1(n6082), .I2(n6081), .O(n6057) );
  NAND3_GATE U7093 ( .I1(n6078), .I2(n6077), .I3(n6057), .O(n15321) );
  INV_GATE U7094 ( .I1(n15321), .O(n6073) );
  INV_GATE U7095 ( .I1(n6058), .O(n6059) );
  NAND_GATE U7096 ( .I1(n6059), .I2(n6063), .O(n6072) );
  INV_GATE U7097 ( .I1(n6063), .O(n6060) );
  NAND_GATE U7098 ( .I1(n6061), .I2(n6060), .O(n6066) );
  NAND_GATE U7099 ( .I1(n6062), .I2(n6066), .O(n6070) );
  NAND_GATE U7100 ( .I1(n6064), .I2(n6063), .O(n6065) );
  NAND_GATE U7101 ( .I1(n6066), .I2(n6065), .O(n6067) );
  NAND_GATE U7102 ( .I1(n6068), .I2(n6067), .O(n6069) );
  NAND_GATE U7103 ( .I1(n6070), .I2(n6069), .O(n6071) );
  NAND_GATE U7104 ( .I1(n6072), .I2(n6071), .O(n15320) );
  NAND_GATE U7105 ( .I1(n6073), .I2(n15320), .O(n6076) );
  INV_GATE U7106 ( .I1(n15320), .O(n6074) );
  NAND_GATE U7107 ( .I1(n15321), .I2(n6074), .O(n6075) );
  NAND_GATE U7108 ( .I1(n6076), .I2(n6075), .O(\A1[50] ) );
  OR_GATE U7109 ( .I1(n6077), .I2(n6082), .O(n6080) );
  OR_GATE U7110 ( .I1(n6081), .I2(n6078), .O(n6079) );
  AND_GATE U7111 ( .I1(n6080), .I2(n6079), .O(n6087) );
  NAND_GATE U7112 ( .I1(n1108), .I2(n6081), .O(n6085) );
  NAND3_GATE U7113 ( .I1(n6085), .I2(n6084), .I3(n6083), .O(n6086) );
  OR_GATE U7114 ( .I1(n6088), .I2(n6093), .O(n6091) );
  OR_GATE U7115 ( .I1(n6092), .I2(n6089), .O(n6090) );
  NAND_GATE U7116 ( .I1(n1102), .I2(n6092), .O(n6096) );
  NAND3_GATE U7117 ( .I1(n6096), .I2(n6095), .I3(n6094), .O(n6097) );
  INV_GATE U7118 ( .I1(n6970), .O(n6973) );
  NAND_GATE U7119 ( .I1(B[19]), .I2(A[31]), .O(n6977) );
  INV_GATE U7120 ( .I1(n6977), .O(n6971) );
  NAND_GATE U7121 ( .I1(n6973), .I2(n6971), .O(n6968) );
  NAND_GATE U7122 ( .I1(B[19]), .I2(A[30]), .O(n6994) );
  INV_GATE U7123 ( .I1(n6994), .O(n6959) );
  OR_GATE U7124 ( .I1(n6098), .I2(n6111), .O(n6101) );
  OR_GATE U7125 ( .I1(n6102), .I2(n6099), .O(n6100) );
  INV_GATE U7126 ( .I1(n6111), .O(n6103) );
  NAND_GATE U7127 ( .I1(n6103), .I2(n6102), .O(n6114) );
  INV_GATE U7128 ( .I1(n6104), .O(n6105) );
  NAND_GATE U7129 ( .I1(n6106), .I2(n6105), .O(n6109) );
  NAND_GATE U7130 ( .I1(n6109), .I2(n6020), .O(n6110) );
  NAND_GATE U7131 ( .I1(n6111), .I2(n6110), .O(n6113) );
  NAND3_GATE U7132 ( .I1(n6114), .I2(n6113), .I3(n6112), .O(n6115) );
  INV_GATE U7133 ( .I1(n6958), .O(n6961) );
  NAND_GATE U7134 ( .I1(n6959), .I2(n6961), .O(n6535) );
  NAND_GATE U7135 ( .I1(B[19]), .I2(A[29]), .O(n7006) );
  INV_GATE U7136 ( .I1(n7006), .O(n6949) );
  INV_GATE U7137 ( .I1(n6117), .O(n6127) );
  NAND_GATE U7138 ( .I1(n6127), .I2(n6122), .O(n6120) );
  INV_GATE U7139 ( .I1(n6122), .O(n6116) );
  NAND_GATE U7140 ( .I1(n6117), .I2(n6116), .O(n6119) );
  NAND3_GATE U7141 ( .I1(n6120), .I2(n6119), .I3(n6118), .O(n6124) );
  OR_GATE U7142 ( .I1(n6122), .I2(n6121), .O(n6123) );
  NAND_GATE U7143 ( .I1(n6124), .I2(n6123), .O(n6128) );
  INV_GATE U7144 ( .I1(n6125), .O(n6126) );
  INV_GATE U7145 ( .I1(n6945), .O(n6946) );
  NAND_GATE U7146 ( .I1(n6949), .I2(n6946), .O(n6950) );
  NAND_GATE U7147 ( .I1(n7006), .I2(n6128), .O(n6531) );
  NAND_GATE U7148 ( .I1(n7006), .I2(n283), .O(n6530) );
  OR_GATE U7149 ( .I1(n6129), .I2(n6134), .O(n6132) );
  OR_GATE U7150 ( .I1(n6133), .I2(n6130), .O(n6131) );
  AND_GATE U7151 ( .I1(n6132), .I2(n6131), .O(n6139) );
  NAND_GATE U7152 ( .I1(n6134), .I2(n1159), .O(n6136) );
  NAND3_GATE U7153 ( .I1(n6137), .I2(n6136), .I3(n6135), .O(n6138) );
  NAND_GATE U7154 ( .I1(n6139), .I2(n6138), .O(n6927) );
  INV_GATE U7155 ( .I1(n6927), .O(n6928) );
  NAND_GATE U7156 ( .I1(B[19]), .I2(A[28]), .O(n6938) );
  INV_GATE U7157 ( .I1(n6938), .O(n6931) );
  NAND_GATE U7158 ( .I1(n6928), .I2(n6931), .O(n6932) );
  OR_GATE U7159 ( .I1(n6140), .I2(n6145), .O(n6143) );
  OR_GATE U7160 ( .I1(n6144), .I2(n6141), .O(n6142) );
  AND_GATE U7161 ( .I1(n6143), .I2(n6142), .O(n6150) );
  NAND_GATE U7162 ( .I1(n6145), .I2(n1147), .O(n6147) );
  NAND3_GATE U7163 ( .I1(n6148), .I2(n6147), .I3(n6146), .O(n6149) );
  NAND_GATE U7164 ( .I1(n6150), .I2(n6149), .O(n6910) );
  INV_GATE U7165 ( .I1(n6910), .O(n6911) );
  NAND_GATE U7166 ( .I1(B[19]), .I2(A[27]), .O(n6921) );
  INV_GATE U7167 ( .I1(n6921), .O(n6914) );
  NAND_GATE U7168 ( .I1(n6911), .I2(n6914), .O(n6915) );
  NAND_GATE U7169 ( .I1(B[19]), .I2(A[26]), .O(n6905) );
  INV_GATE U7170 ( .I1(n6905), .O(n6897) );
  OR_GATE U7171 ( .I1(n6151), .I2(n6156), .O(n6154) );
  OR_GATE U7172 ( .I1(n6155), .I2(n6152), .O(n6153) );
  AND_GATE U7173 ( .I1(n6154), .I2(n6153), .O(n6161) );
  NAND_GATE U7174 ( .I1(n6156), .I2(n1146), .O(n6158) );
  NAND3_GATE U7175 ( .I1(n6159), .I2(n6158), .I3(n6157), .O(n6160) );
  NAND_GATE U7176 ( .I1(n6161), .I2(n6160), .O(n6893) );
  INV_GATE U7177 ( .I1(n6893), .O(n6894) );
  NAND_GATE U7178 ( .I1(n6897), .I2(n6894), .O(n6898) );
  OR_GATE U7179 ( .I1(n6162), .I2(n6167), .O(n6165) );
  OR_GATE U7180 ( .I1(n6166), .I2(n6163), .O(n6164) );
  AND_GATE U7181 ( .I1(n6165), .I2(n6164), .O(n6172) );
  NAND_GATE U7182 ( .I1(n1145), .I2(n6166), .O(n6170) );
  NAND3_GATE U7183 ( .I1(n6170), .I2(n6169), .I3(n6168), .O(n6171) );
  NAND_GATE U7184 ( .I1(n6172), .I2(n6171), .O(n6876) );
  INV_GATE U7185 ( .I1(n6876), .O(n6877) );
  NAND_GATE U7186 ( .I1(B[19]), .I2(A[25]), .O(n6888) );
  INV_GATE U7187 ( .I1(n6888), .O(n6880) );
  NAND_GATE U7188 ( .I1(n6877), .I2(n6880), .O(n6881) );
  OR_GATE U7189 ( .I1(n6173), .I2(n6178), .O(n6176) );
  OR_GATE U7190 ( .I1(n6177), .I2(n6174), .O(n6175) );
  AND_GATE U7191 ( .I1(n6176), .I2(n6175), .O(n6183) );
  NAND_GATE U7192 ( .I1(n1164), .I2(n6177), .O(n6181) );
  NAND3_GATE U7193 ( .I1(n6181), .I2(n6180), .I3(n6179), .O(n6182) );
  NAND_GATE U7194 ( .I1(n6183), .I2(n6182), .O(n6861) );
  INV_GATE U7195 ( .I1(n6861), .O(n6862) );
  NAND_GATE U7196 ( .I1(B[19]), .I2(A[24]), .O(n6872) );
  INV_GATE U7197 ( .I1(n6872), .O(n6865) );
  NAND_GATE U7198 ( .I1(B[19]), .I2(A[23]), .O(n6856) );
  INV_GATE U7199 ( .I1(n6856), .O(n6849) );
  OR_GATE U7200 ( .I1(n6184), .I2(n6189), .O(n6187) );
  OR_GATE U7201 ( .I1(n6188), .I2(n6185), .O(n6186) );
  AND_GATE U7202 ( .I1(n6187), .I2(n6186), .O(n6194) );
  NAND_GATE U7203 ( .I1(n1158), .I2(n6188), .O(n6192) );
  NAND3_GATE U7204 ( .I1(n6192), .I2(n6191), .I3(n6190), .O(n6193) );
  NAND_GATE U7205 ( .I1(n6194), .I2(n6193), .O(n6848) );
  INV_GATE U7206 ( .I1(n6848), .O(n6844) );
  OR_GATE U7207 ( .I1(n6199), .I2(n6195), .O(n6198) );
  OR_GATE U7208 ( .I1(n6200), .I2(n6196), .O(n6197) );
  AND_GATE U7209 ( .I1(n6198), .I2(n6197), .O(n6205) );
  NAND_GATE U7210 ( .I1(n1144), .I2(n6199), .O(n6203) );
  NAND3_GATE U7211 ( .I1(n6203), .I2(n6202), .I3(n6201), .O(n6204) );
  NAND_GATE U7212 ( .I1(n6205), .I2(n6204), .O(n6831) );
  NAND_GATE U7213 ( .I1(B[19]), .I2(A[22]), .O(n6839) );
  INV_GATE U7214 ( .I1(n6839), .O(n6832) );
  NAND_GATE U7215 ( .I1(n6828), .I2(n6832), .O(n6833) );
  OR_GATE U7216 ( .I1(n6206), .I2(n6215), .O(n6209) );
  OR_GATE U7217 ( .I1(n6210), .I2(n6207), .O(n6208) );
  AND_GATE U7218 ( .I1(n6209), .I2(n6208), .O(n6220) );
  NAND_GATE U7219 ( .I1(n6213), .I2(n5881), .O(n6214) );
  NAND_GATE U7220 ( .I1(n6215), .I2(n6214), .O(n6217) );
  NAND3_GATE U7221 ( .I1(n6218), .I2(n6217), .I3(n6216), .O(n6219) );
  NAND_GATE U7222 ( .I1(n6220), .I2(n6219), .O(n6813) );
  NAND_GATE U7223 ( .I1(B[19]), .I2(A[21]), .O(n6823) );
  INV_GATE U7224 ( .I1(n6823), .O(n6815) );
  NAND_GATE U7225 ( .I1(n778), .I2(n6815), .O(n6816) );
  NAND_GATE U7226 ( .I1(B[19]), .I2(A[20]), .O(n6804) );
  INV_GATE U7227 ( .I1(n6804), .O(n6799) );
  NAND_GATE U7228 ( .I1(B[19]), .I2(A[19]), .O(n6791) );
  INV_GATE U7229 ( .I1(n6791), .O(n6785) );
  INV_GATE U7230 ( .I1(n6230), .O(n6231) );
  INV_GATE U7231 ( .I1(n6222), .O(n6223) );
  NAND_GATE U7232 ( .I1(n6224), .I2(n6223), .O(n6228) );
  NAND_GATE U7233 ( .I1(n6226), .I2(n6225), .O(n6227) );
  NAND_GATE U7234 ( .I1(n6228), .I2(n6227), .O(n6229) );
  NAND_GATE U7235 ( .I1(n6230), .I2(n6229), .O(n6236) );
  NAND_GATE U7236 ( .I1(n6231), .I2(n6232), .O(n6235) );
  NAND3_GATE U7237 ( .I1(n6237), .I2(n6236), .I3(n6235), .O(n6234) );
  NAND3_GATE U7238 ( .I1(n6238), .I2(n6234), .I3(n6239), .O(n6783) );
  NAND4_GATE U7239 ( .I1(n6237), .I2(n6236), .I3(n6235), .I4(n6791), .O(n6500)
         );
  NAND_GATE U7240 ( .I1(n6239), .I2(n6238), .O(n6240) );
  NAND_GATE U7241 ( .I1(n6791), .I2(n6240), .O(n6499) );
  NAND_GATE U7242 ( .I1(n6244), .I2(n1148), .O(n6242) );
  NAND3_GATE U7243 ( .I1(n6243), .I2(n6242), .I3(n6241), .O(n6250) );
  OR_GATE U7244 ( .I1(n6245), .I2(n6244), .O(n6249) );
  OR_GATE U7245 ( .I1(n6247), .I2(n6246), .O(n6248) );
  NAND3_GATE U7246 ( .I1(n6250), .I2(n6249), .I3(n6248), .O(n6774) );
  INV_GATE U7247 ( .I1(n6774), .O(n6772) );
  NAND_GATE U7248 ( .I1(B[19]), .I2(A[18]), .O(n6773) );
  INV_GATE U7249 ( .I1(n6773), .O(n6770) );
  NAND_GATE U7250 ( .I1(B[19]), .I2(A[17]), .O(n7149) );
  INV_GATE U7251 ( .I1(n7149), .O(n6759) );
  INV_GATE U7252 ( .I1(n6265), .O(n6255) );
  NAND_GATE U7253 ( .I1(n6254), .I2(n6253), .O(n6257) );
  NAND3_GATE U7254 ( .I1(n6256), .I2(n6255), .I3(n6257), .O(n6261) );
  NAND_GATE U7255 ( .I1(n6257), .I2(n6256), .O(n6258) );
  NAND_GATE U7256 ( .I1(n6265), .I2(n6258), .O(n6260) );
  NAND3_GATE U7257 ( .I1(n6261), .I2(n6260), .I3(n6259), .O(n6268) );
  OR_GATE U7258 ( .I1(n6263), .I2(n6262), .O(n6267) );
  OR_GATE U7259 ( .I1(n6265), .I2(n6264), .O(n6266) );
  NAND3_GATE U7260 ( .I1(n6268), .I2(n6267), .I3(n6266), .O(n6762) );
  NAND_GATE U7261 ( .I1(n6759), .I2(n708), .O(n6496) );
  NAND_GATE U7262 ( .I1(B[19]), .I2(A[16]), .O(n7429) );
  INV_GATE U7263 ( .I1(n7429), .O(n6754) );
  NAND_GATE U7264 ( .I1(n1040), .I2(n6275), .O(n6271) );
  NAND3_GATE U7265 ( .I1(n6271), .I2(n6270), .I3(n6269), .O(n6278) );
  OR_GATE U7266 ( .I1(n6273), .I2(n6272), .O(n6277) );
  OR_GATE U7267 ( .I1(n6275), .I2(n6274), .O(n6276) );
  NAND3_GATE U7268 ( .I1(n6278), .I2(n6277), .I3(n6276), .O(n7425) );
  INV_GATE U7269 ( .I1(n7425), .O(n7424) );
  NAND_GATE U7270 ( .I1(n6754), .I2(n7424), .O(n6753) );
  NAND_GATE U7271 ( .I1(B[19]), .I2(A[15]), .O(n6748) );
  INV_GATE U7272 ( .I1(n6748), .O(n7167) );
  NAND4_GATE U7273 ( .I1(n6282), .I2(n6283), .I3(n6281), .I4(n6290), .O(n6287)
         );
  NAND_GATE U7274 ( .I1(n6283), .I2(n6290), .O(n6284) );
  NAND_GATE U7275 ( .I1(n6288), .I2(n6284), .O(n6286) );
  NAND3_GATE U7276 ( .I1(n6287), .I2(n6286), .I3(n6285), .O(n6296) );
  OR_GATE U7277 ( .I1(n6289), .I2(n6288), .O(n6295) );
  NAND_GATE U7278 ( .I1(n6291), .I2(n6290), .O(n6292) );
  NAND3_GATE U7279 ( .I1(n6293), .I2(n6292), .I3(n259), .O(n6294) );
  NAND3_GATE U7280 ( .I1(n6296), .I2(n6295), .I3(n6294), .O(n6750) );
  INV_GATE U7281 ( .I1(n6750), .O(n6751) );
  NAND_GATE U7282 ( .I1(n7167), .I2(n6751), .O(n6491) );
  NAND_GATE U7283 ( .I1(B[19]), .I2(A[13]), .O(n6547) );
  INV_GATE U7284 ( .I1(n6547), .O(n6541) );
  NAND_GATE U7285 ( .I1(B[19]), .I2(A[11]), .O(n6564) );
  INV_GATE U7286 ( .I1(n6564), .O(n6552) );
  NAND_GATE U7287 ( .I1(B[19]), .I2(A[9]), .O(n6692) );
  INV_GATE U7288 ( .I1(n6692), .O(n6403) );
  NAND_GATE U7289 ( .I1(B[19]), .I2(A[8]), .O(n6570) );
  INV_GATE U7290 ( .I1(n6570), .O(n6581) );
  NAND_GATE U7291 ( .I1(n6297), .I2(n6308), .O(n6300) );
  INV_GATE U7292 ( .I1(n6298), .O(n6299) );
  NAND3_GATE U7293 ( .I1(n6300), .I2(n6299), .I3(n6304), .O(n6303) );
  INV_GATE U7294 ( .I1(n6311), .O(n6307) );
  NAND4_GATE U7295 ( .I1(n6301), .I2(n6309), .I3(n6307), .I4(n6308), .O(n6302)
         );
  AND_GATE U7296 ( .I1(n6303), .I2(n6302), .O(n6573) );
  NAND_GATE U7297 ( .I1(n713), .I2(n6304), .O(n6309) );
  NAND_GATE U7298 ( .I1(n6306), .I2(n6305), .O(n6308) );
  NAND3_GATE U7299 ( .I1(n6307), .I2(n6309), .I3(n6308), .O(n6313) );
  NAND_GATE U7300 ( .I1(n6309), .I2(n6308), .O(n6310) );
  NAND_GATE U7301 ( .I1(n6311), .I2(n6310), .O(n6312) );
  NAND3_GATE U7302 ( .I1(n6314), .I2(n6313), .I3(n6312), .O(n6571) );
  NAND_GATE U7303 ( .I1(n6573), .I2(n6571), .O(n6575) );
  NAND_GATE U7304 ( .I1(n6581), .I2(n1331), .O(n6388) );
  NAND_GATE U7305 ( .I1(B[19]), .I2(A[7]), .O(n6602) );
  INV_GATE U7306 ( .I1(n6602), .O(n6587) );
  INV_GATE U7307 ( .I1(n6323), .O(n6317) );
  NAND_GATE U7308 ( .I1(n6318), .I2(n6317), .O(n6315) );
  NAND_GATE U7309 ( .I1(n6316), .I2(n6315), .O(n6321) );
  NAND_GATE U7310 ( .I1(n6321), .I2(n6320), .O(n6326) );
  INV_GATE U7311 ( .I1(n6322), .O(n6324) );
  NAND_GATE U7312 ( .I1(n6324), .I2(n6323), .O(n6325) );
  NAND_GATE U7313 ( .I1(n6326), .I2(n6325), .O(n6612) );
  OR_GATE U7314 ( .I1(n6334), .I2(n6328), .O(n6329) );
  AND_GATE U7315 ( .I1(n6330), .I2(n6329), .O(n6340) );
  NAND3_GATE U7316 ( .I1(n6333), .I2(n6332), .I3(n6331), .O(n6337) );
  INV_GATE U7317 ( .I1(n6333), .O(n6335) );
  NAND_GATE U7318 ( .I1(n6335), .I2(n6334), .O(n6336) );
  NAND3_GATE U7319 ( .I1(n6338), .I2(n6337), .I3(n6336), .O(n6339) );
  NAND_GATE U7320 ( .I1(n6340), .I2(n6339), .O(n6660) );
  INV_GATE U7321 ( .I1(n6660), .O(n6662) );
  NAND_GATE U7322 ( .I1(B[19]), .I2(A[4]), .O(n6666) );
  INV_GATE U7323 ( .I1(n6666), .O(n6658) );
  NAND_GATE U7324 ( .I1(n6662), .I2(n6658), .O(n6656) );
  NAND_GATE U7325 ( .I1(B[19]), .I2(A[3]), .O(n6627) );
  INV_GATE U7326 ( .I1(n6627), .O(n6360) );
  NAND_GATE U7327 ( .I1(B[19]), .I2(A[2]), .O(n6647) );
  INV_GATE U7328 ( .I1(n6647), .O(n6641) );
  NAND_GATE U7329 ( .I1(n1386), .I2(A[0]), .O(n6341) );
  NAND_GATE U7330 ( .I1(n14781), .I2(n6341), .O(n6342) );
  NAND_GATE U7331 ( .I1(B[21]), .I2(n6342), .O(n6346) );
  NAND_GATE U7332 ( .I1(n1387), .I2(A[1]), .O(n6343) );
  NAND_GATE U7333 ( .I1(n14784), .I2(n6343), .O(n6344) );
  NAND_GATE U7334 ( .I1(B[20]), .I2(n6344), .O(n6345) );
  NAND_GATE U7335 ( .I1(n6346), .I2(n6345), .O(n6643) );
  NAND_GATE U7336 ( .I1(n6641), .I2(n6643), .O(n6638) );
  NAND3_GATE U7337 ( .I1(B[19]), .I2(B[20]), .I3(n1196), .O(n6639) );
  INV_GATE U7338 ( .I1(n6639), .O(n6642) );
  INV_GATE U7339 ( .I1(n6643), .O(n6640) );
  NAND_GATE U7340 ( .I1(n6647), .I2(n6640), .O(n6347) );
  NAND_GATE U7341 ( .I1(n6642), .I2(n6347), .O(n6348) );
  NAND_GATE U7342 ( .I1(n6638), .I2(n6348), .O(n6622) );
  NAND_GATE U7343 ( .I1(n6360), .I2(n6622), .O(n6617) );
  NAND_GATE U7344 ( .I1(n6350), .I2(n6353), .O(n6357) );
  NAND_GATE U7345 ( .I1(n6351), .I2(n6359), .O(n6352) );
  NAND_GATE U7346 ( .I1(n6353), .I2(n6352), .O(n6354) );
  NAND_GATE U7347 ( .I1(n6355), .I2(n6354), .O(n6356) );
  NAND_GATE U7348 ( .I1(n6357), .I2(n6356), .O(n6620) );
  NAND_GATE U7349 ( .I1(n6620), .I2(n6621), .O(n6623) );
  NAND_GATE U7350 ( .I1(n6622), .I2(n6623), .O(n6361) );
  NAND_GATE U7351 ( .I1(n6360), .I2(n6623), .O(n6616) );
  NAND3_GATE U7352 ( .I1(n6617), .I2(n6361), .I3(n6616), .O(n6661) );
  NAND_GATE U7353 ( .I1(n6660), .I2(n6666), .O(n6362) );
  NAND_GATE U7354 ( .I1(n6661), .I2(n6362), .O(n6363) );
  NAND_GATE U7355 ( .I1(n6656), .I2(n6363), .O(n6609) );
  NAND_GATE U7356 ( .I1(n6612), .I2(n6609), .O(n6365) );
  NAND_GATE U7357 ( .I1(B[19]), .I2(A[5]), .O(n6613) );
  INV_GATE U7358 ( .I1(n6613), .O(n6364) );
  NAND_GATE U7359 ( .I1(n6364), .I2(n6609), .O(n6607) );
  NAND_GATE U7360 ( .I1(n6364), .I2(n6612), .O(n6606) );
  NAND3_GATE U7361 ( .I1(n6365), .I2(n6607), .I3(n6606), .O(n6681) );
  INV_GATE U7362 ( .I1(n6370), .O(n6372) );
  NAND3_GATE U7363 ( .I1(n6372), .I2(n6366), .I3(n6371), .O(n6369) );
  OR_GATE U7364 ( .I1(n6371), .I2(n6367), .O(n6368) );
  AND_GATE U7365 ( .I1(n6369), .I2(n6368), .O(n6377) );
  NAND_GATE U7366 ( .I1(n6372), .I2(n6371), .O(n6373) );
  NAND3_GATE U7367 ( .I1(n6375), .I2(n6374), .I3(n6373), .O(n6376) );
  NAND_GATE U7368 ( .I1(n6377), .I2(n6376), .O(n6678) );
  NAND_GATE U7369 ( .I1(B[19]), .I2(A[6]), .O(n7248) );
  NAND_GATE U7370 ( .I1(n6678), .I2(n7248), .O(n6378) );
  NAND_GATE U7371 ( .I1(n6681), .I2(n6378), .O(n6380) );
  INV_GATE U7372 ( .I1(n7248), .O(n6677) );
  NAND_GATE U7373 ( .I1(n6680), .I2(n6677), .O(n6379) );
  NAND_GATE U7374 ( .I1(n6380), .I2(n6379), .O(n6597) );
  NAND_GATE U7375 ( .I1(n6587), .I2(n6597), .O(n6596) );
  INV_GATE U7376 ( .I1(n6588), .O(n6591) );
  NAND_GATE U7377 ( .I1(n1067), .I2(n6382), .O(n6592) );
  NAND3_GATE U7378 ( .I1(n6588), .I2(n1067), .I3(n1206), .O(n6595) );
  NAND_GATE U7379 ( .I1(n6591), .I2(n6590), .O(n6382) );
  NAND_GATE U7380 ( .I1(n6588), .I2(n1206), .O(n6381) );
  NAND_GATE U7381 ( .I1(n6382), .I2(n6381), .O(n6383) );
  NAND_GATE U7382 ( .I1(n6589), .I2(n6383), .O(n6585) );
  NAND3_GATE U7383 ( .I1(n6587), .I2(n6586), .I3(n6585), .O(n6385) );
  NAND3_GATE U7384 ( .I1(n6597), .I2(n6586), .I3(n6585), .O(n6384) );
  NAND3_GATE U7385 ( .I1(n6596), .I2(n6385), .I3(n6384), .O(n6572) );
  NAND_GATE U7386 ( .I1(n6570), .I2(n6575), .O(n6386) );
  NAND_GATE U7387 ( .I1(n6572), .I2(n6386), .O(n6387) );
  NAND_GATE U7388 ( .I1(n6403), .I2(n518), .O(n6696) );
  NAND_GATE U7389 ( .I1(n6391), .I2(n6399), .O(n6394) );
  INV_GATE U7390 ( .I1(n6394), .O(n6389) );
  NAND3_GATE U7391 ( .I1(n794), .I2(n6392), .I3(n6389), .O(n6401) );
  NAND3_GATE U7392 ( .I1(n735), .I2(n6390), .I3(n6398), .O(n6397) );
  NAND3_GATE U7393 ( .I1(n794), .I2(n6392), .I3(n6399), .O(n6393) );
  NAND4_GATE U7394 ( .I1(n6397), .I2(n6396), .I3(n6394), .I4(n6393), .O(n6395)
         );
  NAND_GATE U7395 ( .I1(n6401), .I2(n6395), .O(n6697) );
  NAND_GATE U7396 ( .I1(n518), .I2(n6697), .O(n6405) );
  NAND_GATE U7397 ( .I1(n735), .I2(n6398), .O(n6400) );
  NAND3_GATE U7398 ( .I1(n6401), .I2(n6400), .I3(n6399), .O(n6402) );
  AND_GATE U7399 ( .I1(n6403), .I2(n6402), .O(n6695) );
  NAND_GATE U7400 ( .I1(n991), .I2(n6695), .O(n6404) );
  NAND3_GATE U7401 ( .I1(n6696), .I2(n6405), .I3(n6404), .O(n6705) );
  NAND_GATE U7402 ( .I1(B[19]), .I2(A[10]), .O(n7200) );
  INV_GATE U7403 ( .I1(n6409), .O(n6411) );
  NAND4_GATE U7404 ( .I1(n6407), .I2(n6411), .I3(n1161), .I4(n6406), .O(n6417)
         );
  OR_GATE U7405 ( .I1(n6410), .I2(n6408), .O(n6416) );
  NAND_GATE U7406 ( .I1(n6411), .I2(n6410), .O(n6412) );
  NAND3_GATE U7407 ( .I1(n6414), .I2(n6413), .I3(n6412), .O(n6415) );
  NAND3_GATE U7408 ( .I1(n6417), .I2(n6416), .I3(n6415), .O(n6706) );
  NAND_GATE U7409 ( .I1(n7200), .I2(n6706), .O(n6418) );
  NAND_GATE U7410 ( .I1(n6705), .I2(n6418), .O(n6420) );
  INV_GATE U7411 ( .I1(n7200), .O(n7204) );
  NAND_GATE U7412 ( .I1(n7204), .I2(n674), .O(n6419) );
  NAND_GATE U7413 ( .I1(n6420), .I2(n6419), .O(n6563) );
  NAND_GATE U7414 ( .I1(n6552), .I2(n6563), .O(n6554) );
  NAND3_GATE U7415 ( .I1(n6423), .I2(n6422), .I3(n784), .O(n6559) );
  NAND_GATE U7416 ( .I1(n785), .I2(n6559), .O(n6551) );
  NAND_GATE U7417 ( .I1(n6423), .I2(n784), .O(n6424) );
  NAND_GATE U7418 ( .I1(n6424), .I2(n6421), .O(n6557) );
  NAND3_GATE U7419 ( .I1(n6563), .I2(n6551), .I3(n6561), .O(n6426) );
  NAND3_GATE U7420 ( .I1(n6552), .I2(n6551), .I3(n6561), .O(n6425) );
  NAND_GATE U7421 ( .I1(B[19]), .I2(A[12]), .O(n7366) );
  INV_GATE U7422 ( .I1(n6442), .O(n6439) );
  NAND4_GATE U7423 ( .I1(n6428), .I2(n6439), .I3(n1165), .I4(n6427), .O(n6448)
         );
  NAND3_GATE U7424 ( .I1(n6431), .I2(n6430), .I3(n6429), .O(n6434) );
  NAND4_GATE U7425 ( .I1(n6435), .I2(n6434), .I3(n6433), .I4(n6432), .O(n6436)
         );
  NAND_GATE U7426 ( .I1(n6437), .I2(n6436), .O(n6440) );
  OR_GATE U7427 ( .I1(n6440), .I2(n6438), .O(n6447) );
  NAND_GATE U7428 ( .I1(n6439), .I2(n6440), .O(n6444) );
  INV_GATE U7429 ( .I1(n6440), .O(n6441) );
  NAND_GATE U7430 ( .I1(n6442), .I2(n6441), .O(n6443) );
  NAND3_GATE U7431 ( .I1(n6445), .I2(n6444), .I3(n6443), .O(n6446) );
  NAND3_GATE U7432 ( .I1(n6448), .I2(n6447), .I3(n6446), .O(n6721) );
  NAND_GATE U7433 ( .I1(n7366), .I2(n6721), .O(n6449) );
  NAND_GATE U7434 ( .I1(n7365), .I2(n6449), .O(n6451) );
  INV_GATE U7435 ( .I1(n7366), .O(n6719) );
  NAND_GATE U7436 ( .I1(n6719), .I2(n208), .O(n6450) );
  NAND_GATE U7437 ( .I1(n6541), .I2(n6544), .O(n6542) );
  INV_GATE U7438 ( .I1(n6454), .O(n6455) );
  NAND_GATE U7439 ( .I1(n812), .I2(n6455), .O(n6453) );
  NAND_GATE U7440 ( .I1(n6457), .I2(n6454), .O(n6461) );
  INV_GATE U7441 ( .I1(n6461), .O(n6452) );
  NAND_GATE U7442 ( .I1(n1241), .I2(n6452), .O(n6465) );
  NAND3_GATE U7443 ( .I1(n6457), .I2(n6453), .I3(n6465), .O(n6540) );
  NAND3_GATE U7444 ( .I1(n6456), .I2(n6454), .I3(n1241), .O(n6463) );
  NAND3_GATE U7445 ( .I1(n6456), .I2(n6455), .I3(n812), .O(n6462) );
  NAND3_GATE U7446 ( .I1(n6541), .I2(n6540), .I3(n951), .O(n6467) );
  NAND3_GATE U7447 ( .I1(n6459), .I2(n6458), .I3(n6457), .O(n6460) );
  NAND4_GATE U7448 ( .I1(n6463), .I2(n6462), .I3(n6461), .I4(n6460), .O(n6464)
         );
  NAND_GATE U7449 ( .I1(n6465), .I2(n6464), .O(n6543) );
  NAND_GATE U7450 ( .I1(n6544), .I2(n6543), .O(n6466) );
  NAND_GATE U7451 ( .I1(B[19]), .I2(A[14]), .O(n6745) );
  INV_GATE U7452 ( .I1(n6479), .O(n6477) );
  NAND4_GATE U7453 ( .I1(n6470), .I2(n6469), .I3(n6477), .I4(n6468), .O(n6485)
         );
  NAND3_GATE U7454 ( .I1(n6473), .I2(n595), .I3(n6472), .O(n6475) );
  OR_GATE U7455 ( .I1(n6478), .I2(n6476), .O(n6484) );
  NAND_GATE U7456 ( .I1(n6477), .I2(n6478), .O(n6481) );
  NAND3_GATE U7457 ( .I1(n6482), .I2(n6481), .I3(n6480), .O(n6483) );
  NAND3_GATE U7458 ( .I1(n6485), .I2(n6484), .I3(n6483), .O(n6731) );
  NAND_GATE U7459 ( .I1(n6745), .I2(n6731), .O(n6486) );
  NAND_GATE U7460 ( .I1(n6742), .I2(n6486), .O(n6488) );
  INV_GATE U7461 ( .I1(n6745), .O(n6734) );
  INV_GATE U7462 ( .I1(n6731), .O(n6741) );
  NAND_GATE U7463 ( .I1(n6734), .I2(n6741), .O(n6487) );
  NAND_GATE U7464 ( .I1(n6488), .I2(n6487), .O(n6752) );
  NAND_GATE U7465 ( .I1(n6748), .I2(n6750), .O(n6489) );
  NAND_GATE U7466 ( .I1(n6752), .I2(n6489), .O(n6490) );
  NAND_GATE U7467 ( .I1(n7429), .I2(n7425), .O(n6492) );
  NAND_GATE U7468 ( .I1(n7423), .I2(n6492), .O(n6493) );
  NAND_GATE U7469 ( .I1(n6753), .I2(n6493), .O(n6760) );
  NAND_GATE U7470 ( .I1(n7149), .I2(n6762), .O(n6494) );
  NAND_GATE U7471 ( .I1(n6760), .I2(n6494), .O(n6495) );
  NAND_GATE U7472 ( .I1(n6774), .I2(n6773), .O(n6497) );
  NAND_GATE U7473 ( .I1(n6771), .I2(n6497), .O(n6498) );
  NAND3_GATE U7474 ( .I1(n6500), .I2(n6499), .I3(n6787), .O(n6501) );
  NAND_GATE U7475 ( .I1(n6799), .I2(n664), .O(n6797) );
  OR_GATE U7476 ( .I1(n6507), .I2(n6502), .O(n6505) );
  NAND3_GATE U7477 ( .I1(n6507), .I2(n1268), .I3(n6503), .O(n6504) );
  NAND_GATE U7478 ( .I1(n6507), .I2(n1268), .O(n6509) );
  NAND3_GATE U7479 ( .I1(n6510), .I2(n6509), .I3(n6508), .O(n6511) );
  INV_GATE U7480 ( .I1(n6801), .O(n6800) );
  NAND_GATE U7481 ( .I1(n6804), .I2(n824), .O(n6512) );
  NAND_GATE U7482 ( .I1(n6800), .I2(n6512), .O(n6513) );
  NAND_GATE U7483 ( .I1(n6797), .I2(n6513), .O(n6817) );
  NAND_GATE U7484 ( .I1(n6813), .I2(n6823), .O(n6514) );
  NAND_GATE U7485 ( .I1(n6817), .I2(n6514), .O(n6515) );
  NAND_GATE U7486 ( .I1(n6831), .I2(n6839), .O(n6516) );
  NAND_GATE U7487 ( .I1(n618), .I2(n6516), .O(n6517) );
  NAND_GATE U7488 ( .I1(n6833), .I2(n6517), .O(n6851) );
  NAND_GATE U7489 ( .I1(n6856), .I2(n6848), .O(n6518) );
  NAND_GATE U7490 ( .I1(n6851), .I2(n6518), .O(n6519) );
  NAND_GATE U7491 ( .I1(n6850), .I2(n6519), .O(n6867) );
  NAND_GATE U7492 ( .I1(n6861), .I2(n6872), .O(n6520) );
  NAND_GATE U7493 ( .I1(n6867), .I2(n6520), .O(n6521) );
  NAND_GATE U7494 ( .I1(n6866), .I2(n6521), .O(n6882) );
  NAND_GATE U7495 ( .I1(n6876), .I2(n6888), .O(n6522) );
  NAND_GATE U7496 ( .I1(n6882), .I2(n6522), .O(n6523) );
  NAND_GATE U7497 ( .I1(n6881), .I2(n6523), .O(n6899) );
  NAND_GATE U7498 ( .I1(n6905), .I2(n6893), .O(n6524) );
  NAND_GATE U7499 ( .I1(n6899), .I2(n6524), .O(n6525) );
  NAND_GATE U7500 ( .I1(n6898), .I2(n6525), .O(n6916) );
  NAND_GATE U7501 ( .I1(n6910), .I2(n6921), .O(n6526) );
  NAND_GATE U7502 ( .I1(n6916), .I2(n6526), .O(n6527) );
  NAND_GATE U7503 ( .I1(n6915), .I2(n6527), .O(n6933) );
  NAND_GATE U7504 ( .I1(n6927), .I2(n6938), .O(n6528) );
  NAND_GATE U7505 ( .I1(n6933), .I2(n6528), .O(n6529) );
  NAND_GATE U7506 ( .I1(n6932), .I2(n6529), .O(n6951) );
  NAND3_GATE U7507 ( .I1(n6531), .I2(n6530), .I3(n6951), .O(n6532) );
  NAND_GATE U7508 ( .I1(n6950), .I2(n6532), .O(n6960) );
  NAND_GATE U7509 ( .I1(n6994), .I2(n6958), .O(n6533) );
  NAND_GATE U7510 ( .I1(n6960), .I2(n6533), .O(n6534) );
  NAND_GATE U7511 ( .I1(n6535), .I2(n6534), .O(n6972) );
  NAND_GATE U7512 ( .I1(n6970), .I2(n6977), .O(n6536) );
  NAND_GATE U7513 ( .I1(n6972), .I2(n6536), .O(n6537) );
  NAND_GATE U7514 ( .I1(n6968), .I2(n6537), .O(n6538) );
  NAND_GATE U7515 ( .I1(n156), .I2(n6538), .O(n15322) );
  AND_GATE U7516 ( .I1(n15322), .I2(n6539), .O(\A1[49] ) );
  NAND_GATE U7517 ( .I1(B[18]), .I2(A[31]), .O(n6998) );
  INV_GATE U7518 ( .I1(n6998), .O(n6966) );
  NAND_GATE U7519 ( .I1(B[18]), .I2(A[30]), .O(n7010) );
  INV_GATE U7520 ( .I1(n7010), .O(n6952) );
  NAND_GATE U7521 ( .I1(B[18]), .I2(A[29]), .O(n7021) );
  INV_GATE U7522 ( .I1(n7021), .O(n6935) );
  NAND_GATE U7523 ( .I1(B[18]), .I2(A[28]), .O(n7039) );
  INV_GATE U7524 ( .I1(n7039), .O(n6918) );
  NAND_GATE U7525 ( .I1(B[18]), .I2(A[27]), .O(n7050) );
  INV_GATE U7526 ( .I1(n7050), .O(n6901) );
  NAND_GATE U7527 ( .I1(B[18]), .I2(A[26]), .O(n7061) );
  INV_GATE U7528 ( .I1(n7061), .O(n6884) );
  NAND_GATE U7529 ( .I1(B[18]), .I2(A[25]), .O(n7072) );
  INV_GATE U7530 ( .I1(n7072), .O(n6868) );
  NAND_GATE U7531 ( .I1(B[18]), .I2(A[24]), .O(n7083) );
  INV_GATE U7532 ( .I1(n7083), .O(n6852) );
  NAND_GATE U7533 ( .I1(B[18]), .I2(A[23]), .O(n7094) );
  INV_GATE U7534 ( .I1(n7094), .O(n6835) );
  NAND_GATE U7535 ( .I1(B[18]), .I2(A[22]), .O(n7105) );
  INV_GATE U7536 ( .I1(n7105), .O(n6819) );
  NAND_GATE U7537 ( .I1(B[18]), .I2(A[21]), .O(n7116) );
  INV_GATE U7538 ( .I1(n7116), .O(n6809) );
  NAND_GATE U7539 ( .I1(B[18]), .I2(A[20]), .O(n7132) );
  INV_GATE U7540 ( .I1(n7132), .O(n6789) );
  NAND_GATE U7541 ( .I1(B[18]), .I2(A[19]), .O(n7136) );
  INV_GATE U7542 ( .I1(n7136), .O(n7140) );
  NAND_GATE U7543 ( .I1(B[18]), .I2(A[18]), .O(n7154) );
  INV_GATE U7544 ( .I1(n7154), .O(n7158) );
  NAND_GATE U7545 ( .I1(B[18]), .I2(A[17]), .O(n7437) );
  INV_GATE U7546 ( .I1(n7437), .O(n6757) );
  NAND_GATE U7547 ( .I1(B[18]), .I2(A[16]), .O(n7177) );
  INV_GATE U7548 ( .I1(n7177), .O(n7165) );
  NAND_GATE U7549 ( .I1(B[18]), .I2(A[15]), .O(n7406) );
  INV_GATE U7550 ( .I1(n7406), .O(n6740) );
  NAND_GATE U7551 ( .I1(B[18]), .I2(A[14]), .O(n7388) );
  INV_GATE U7552 ( .I1(n7388), .O(n7181) );
  NAND4_GATE U7553 ( .I1(n6541), .I2(n20), .I3(n951), .I4(n6540), .O(n6550) );
  OR_GATE U7554 ( .I1(n6543), .I2(n6542), .O(n6549) );
  NAND_GATE U7555 ( .I1(n20), .I2(n6543), .O(n6546) );
  NAND3_GATE U7556 ( .I1(n6547), .I2(n6546), .I3(n6545), .O(n6548) );
  NAND3_GATE U7557 ( .I1(n6550), .I2(n6549), .I3(n6548), .O(n7389) );
  NAND_GATE U7558 ( .I1(n7181), .I2(n816), .O(n6730) );
  NAND_GATE U7559 ( .I1(B[18]), .I2(A[13]), .O(n7375) );
  INV_GATE U7560 ( .I1(n7375), .O(n6724) );
  NAND_GATE U7561 ( .I1(B[18]), .I2(A[12]), .O(n7187) );
  INV_GATE U7562 ( .I1(n7187), .O(n7194) );
  INV_GATE U7563 ( .I1(n6563), .O(n6560) );
  NAND4_GATE U7564 ( .I1(n6552), .I2(n6551), .I3(n6560), .I4(n6561), .O(n6569)
         );
  NAND_GATE U7565 ( .I1(n6553), .I2(n6561), .O(n6556) );
  INV_GATE U7566 ( .I1(n6554), .O(n6555) );
  NAND3_GATE U7567 ( .I1(n6556), .I2(n6555), .I3(n6559), .O(n6568) );
  NAND_GATE U7568 ( .I1(n6558), .I2(n6557), .O(n6561) );
  NAND3_GATE U7569 ( .I1(n6561), .I2(n6560), .I3(n6551), .O(n6566) );
  NAND_GATE U7570 ( .I1(n6551), .I2(n6561), .O(n6562) );
  NAND_GATE U7571 ( .I1(n6563), .I2(n6562), .O(n6565) );
  NAND3_GATE U7572 ( .I1(n6566), .I2(n6565), .I3(n6564), .O(n6567) );
  NAND3_GATE U7573 ( .I1(n6569), .I2(n6568), .I3(n6567), .O(n7190) );
  NAND_GATE U7574 ( .I1(n7194), .I2(n7188), .O(n6717) );
  NAND_GATE U7575 ( .I1(B[18]), .I2(A[11]), .O(n7210) );
  INV_GATE U7576 ( .I1(n7210), .O(n6712) );
  NAND3_GATE U7577 ( .I1(n6570), .I2(n6572), .I3(n1331), .O(n6579) );
  INV_GATE U7578 ( .I1(n6572), .O(n6574) );
  NAND3_GATE U7579 ( .I1(n6570), .I2(n6574), .I3(n6575), .O(n6578) );
  AND_GATE U7580 ( .I1(n6579), .I2(n6578), .O(n6577) );
  NAND4_GATE U7581 ( .I1(n6573), .I2(n6581), .I3(n6572), .I4(n6571), .O(n6584)
         );
  NAND_GATE U7582 ( .I1(n6575), .I2(n6574), .O(n6580) );
  NAND3_GATE U7583 ( .I1(n6584), .I2(n6580), .I3(n6581), .O(n6576) );
  NAND_GATE U7584 ( .I1(B[18]), .I2(A[9]), .O(n7229) );
  INV_GATE U7585 ( .I1(n7229), .O(n6690) );
  NAND3_GATE U7586 ( .I1(n6577), .I2(n6576), .I3(n6690), .O(n7220) );
  NAND_GATE U7587 ( .I1(n6581), .I2(n6580), .O(n6582) );
  NAND_GATE U7588 ( .I1(n6577), .I2(n6582), .O(n6583) );
  NAND_GATE U7589 ( .I1(n6584), .I2(n6583), .O(n7226) );
  NAND_GATE U7590 ( .I1(B[18]), .I2(A[8]), .O(n7235) );
  INV_GATE U7591 ( .I1(n7235), .O(n7233) );
  INV_GATE U7592 ( .I1(n6597), .O(n6599) );
  NAND4_GATE U7593 ( .I1(n6587), .I2(n6586), .I3(n6599), .I4(n6585), .O(n6605)
         );
  NAND3_GATE U7594 ( .I1(n6591), .I2(n6590), .I3(n6589), .O(n6593) );
  NAND3_GATE U7595 ( .I1(n6381), .I2(n6593), .I3(n6592), .O(n6594) );
  NAND_GATE U7596 ( .I1(n6595), .I2(n6594), .O(n6598) );
  OR_GATE U7597 ( .I1(n6598), .I2(n6596), .O(n6604) );
  NAND_GATE U7598 ( .I1(n6599), .I2(n6598), .O(n6600) );
  NAND3_GATE U7599 ( .I1(n6602), .I2(n6601), .I3(n6600), .O(n6603) );
  NAND3_GATE U7600 ( .I1(n6605), .I2(n6604), .I3(n6603), .O(n7236) );
  INV_GATE U7601 ( .I1(n7236), .O(n7234) );
  NAND_GATE U7602 ( .I1(n7233), .I2(n7234), .O(n7240) );
  INV_GATE U7603 ( .I1(n6609), .O(n6611) );
  INV_GATE U7604 ( .I1(n6612), .O(n6610) );
  INV_GATE U7605 ( .I1(n6607), .O(n6608) );
  NAND_GATE U7606 ( .I1(n6610), .I2(n6608), .O(n7330) );
  NAND_GATE U7607 ( .I1(B[18]), .I2(A[6]), .O(n7333) );
  INV_GATE U7608 ( .I1(n7333), .O(n7339) );
  NAND_GATE U7609 ( .I1(n6610), .I2(n6609), .O(n6615) );
  NAND_GATE U7610 ( .I1(n6612), .I2(n6611), .O(n6614) );
  NAND3_GATE U7611 ( .I1(n6615), .I2(n6614), .I3(n6613), .O(n7329) );
  NAND4_GATE U7612 ( .I1(n7331), .I2(n7330), .I3(n7339), .I4(n7329), .O(n6675)
         );
  NAND_GATE U7613 ( .I1(B[18]), .I2(A[5]), .O(n7263) );
  INV_GATE U7614 ( .I1(n7263), .O(n6671) );
  OR_GATE U7615 ( .I1(n6616), .I2(n6622), .O(n6619) );
  OR_GATE U7616 ( .I1(n6623), .I2(n6617), .O(n6618) );
  AND_GATE U7617 ( .I1(n6619), .I2(n6618), .O(n6629) );
  NAND3_GATE U7618 ( .I1(n6622), .I2(n6621), .I3(n6620), .O(n6626) );
  INV_GATE U7619 ( .I1(n6622), .O(n6624) );
  NAND_GATE U7620 ( .I1(n6624), .I2(n6623), .O(n6625) );
  NAND3_GATE U7621 ( .I1(n6627), .I2(n6626), .I3(n6625), .O(n6628) );
  NAND_GATE U7622 ( .I1(n6629), .I2(n6628), .O(n7314) );
  NAND_GATE U7623 ( .I1(B[18]), .I2(A[4]), .O(n7320) );
  INV_GATE U7624 ( .I1(n7320), .O(n7315) );
  NAND_GATE U7625 ( .I1(n553), .I2(n7315), .O(n7311) );
  NAND_GATE U7626 ( .I1(B[18]), .I2(A[3]), .O(n7280) );
  INV_GATE U7627 ( .I1(n7280), .O(n6652) );
  NAND_GATE U7628 ( .I1(B[18]), .I2(A[2]), .O(n7302) );
  INV_GATE U7629 ( .I1(n7302), .O(n7296) );
  NAND_GATE U7630 ( .I1(n1385), .I2(A[0]), .O(n6630) );
  NAND_GATE U7631 ( .I1(n14781), .I2(n6630), .O(n6631) );
  NAND_GATE U7632 ( .I1(B[20]), .I2(n6631), .O(n6635) );
  NAND_GATE U7633 ( .I1(n1386), .I2(A[1]), .O(n6632) );
  NAND_GATE U7634 ( .I1(n14784), .I2(n6632), .O(n6633) );
  NAND_GATE U7635 ( .I1(B[19]), .I2(n6633), .O(n6634) );
  NAND_GATE U7636 ( .I1(n6635), .I2(n6634), .O(n7298) );
  NAND_GATE U7637 ( .I1(n7296), .I2(n7298), .O(n7293) );
  NAND3_GATE U7638 ( .I1(B[18]), .I2(B[19]), .I3(n1196), .O(n7294) );
  INV_GATE U7639 ( .I1(n7294), .O(n7297) );
  INV_GATE U7640 ( .I1(n7298), .O(n7295) );
  NAND_GATE U7641 ( .I1(n7302), .I2(n7295), .O(n6636) );
  NAND_GATE U7642 ( .I1(n7297), .I2(n6636), .O(n6637) );
  NAND_GATE U7643 ( .I1(n7293), .I2(n6637), .O(n7279) );
  NAND_GATE U7644 ( .I1(n6652), .I2(n7279), .O(n7274) );
  OR_GATE U7645 ( .I1(n6639), .I2(n6638), .O(n6651) );
  NAND_GATE U7646 ( .I1(n6640), .I2(n6639), .O(n6645) );
  NAND_GATE U7647 ( .I1(n6641), .I2(n6645), .O(n6649) );
  NAND_GATE U7648 ( .I1(n6643), .I2(n6642), .O(n6644) );
  NAND_GATE U7649 ( .I1(n6645), .I2(n6644), .O(n6646) );
  NAND_GATE U7650 ( .I1(n6647), .I2(n6646), .O(n6648) );
  NAND_GATE U7651 ( .I1(n6649), .I2(n6648), .O(n6650) );
  NAND_GATE U7652 ( .I1(n6651), .I2(n6650), .O(n7278) );
  NAND_GATE U7653 ( .I1(n7279), .I2(n7278), .O(n6653) );
  NAND_GATE U7654 ( .I1(n6652), .I2(n7278), .O(n7273) );
  NAND3_GATE U7655 ( .I1(n7274), .I2(n6653), .I3(n7273), .O(n7316) );
  NAND_GATE U7656 ( .I1(n7314), .I2(n7320), .O(n6654) );
  NAND_GATE U7657 ( .I1(n7316), .I2(n6654), .O(n6655) );
  NAND_GATE U7658 ( .I1(n7311), .I2(n6655), .O(n7266) );
  NAND_GATE U7659 ( .I1(n6671), .I2(n7266), .O(n7268) );
  INV_GATE U7660 ( .I1(n6656), .O(n6657) );
  NAND_GATE U7661 ( .I1(n6657), .I2(n6661), .O(n6670) );
  INV_GATE U7662 ( .I1(n6661), .O(n6659) );
  NAND_GATE U7663 ( .I1(n6658), .I2(n6664), .O(n6668) );
  NAND_GATE U7664 ( .I1(n6660), .I2(n6659), .O(n6664) );
  NAND_GATE U7665 ( .I1(n6662), .I2(n6661), .O(n6663) );
  NAND_GATE U7666 ( .I1(n6664), .I2(n6663), .O(n6665) );
  NAND_GATE U7667 ( .I1(n6666), .I2(n6665), .O(n6667) );
  NAND_GATE U7668 ( .I1(n6668), .I2(n6667), .O(n6669) );
  NAND_GATE U7669 ( .I1(n6670), .I2(n6669), .O(n7269) );
  NAND_GATE U7670 ( .I1(n7266), .I2(n7269), .O(n6672) );
  NAND_GATE U7671 ( .I1(n6671), .I2(n7269), .O(n7267) );
  NAND3_GATE U7672 ( .I1(n7268), .I2(n6672), .I3(n7267), .O(n7340) );
  NAND4_GATE U7673 ( .I1(n7330), .I2(n7329), .I3(n7331), .I4(n7340), .O(n6674)
         );
  NAND_GATE U7674 ( .I1(n7339), .I2(n7340), .O(n6673) );
  NAND3_GATE U7675 ( .I1(n6675), .I2(n6674), .I3(n6673), .O(n7253) );
  NAND3_GATE U7676 ( .I1(n6681), .I2(n6677), .I3(n6680), .O(n7251) );
  INV_GATE U7677 ( .I1(n6681), .O(n6679) );
  NAND_GATE U7678 ( .I1(n6679), .I2(n6678), .O(n6676) );
  NAND_GATE U7679 ( .I1(n6677), .I2(n6676), .O(n7249) );
  NAND_GATE U7680 ( .I1(n6681), .I2(n6680), .O(n6682) );
  NAND_GATE U7681 ( .I1(n6676), .I2(n6682), .O(n7247) );
  NAND_GATE U7682 ( .I1(n7249), .I2(n6683), .O(n6684) );
  NAND_GATE U7683 ( .I1(n7251), .I2(n6684), .O(n7246) );
  NAND_GATE U7684 ( .I1(n7253), .I2(n7246), .O(n6687) );
  NAND_GATE U7685 ( .I1(B[18]), .I2(A[7]), .O(n7257) );
  INV_GATE U7686 ( .I1(n7257), .O(n7245) );
  NAND_GATE U7687 ( .I1(n7245), .I2(n7246), .O(n6686) );
  NAND_GATE U7688 ( .I1(n7245), .I2(n7253), .O(n6685) );
  NAND_GATE U7689 ( .I1(n7235), .I2(n7236), .O(n6688) );
  NAND_GATE U7690 ( .I1(n7241), .I2(n6688), .O(n6689) );
  NAND_GATE U7691 ( .I1(n7240), .I2(n6689), .O(n7224) );
  NAND_GATE U7692 ( .I1(n7226), .I2(n7224), .O(n6691) );
  NAND_GATE U7693 ( .I1(n6690), .I2(n7224), .O(n7221) );
  NAND3_GATE U7694 ( .I1(n7220), .I2(n6691), .I3(n7221), .O(n7354) );
  NAND_GATE U7695 ( .I1(B[18]), .I2(A[10]), .O(n7650) );
  NAND_GATE U7696 ( .I1(n527), .I2(n6697), .O(n6694) );
  NAND3_GATE U7697 ( .I1(n6694), .I2(n6693), .I3(n6692), .O(n6700) );
  NAND3_GATE U7698 ( .I1(n991), .I2(n6695), .I3(n527), .O(n6699) );
  OR_GATE U7699 ( .I1(n6697), .I2(n6696), .O(n6698) );
  NAND3_GATE U7700 ( .I1(n6700), .I2(n6699), .I3(n6698), .O(n7351) );
  NAND_GATE U7701 ( .I1(n7650), .I2(n7351), .O(n6701) );
  NAND_GATE U7702 ( .I1(n7354), .I2(n6701), .O(n6703) );
  INV_GATE U7703 ( .I1(n7650), .O(n7350) );
  NAND_GATE U7704 ( .I1(n7350), .I2(n7353), .O(n6702) );
  NAND_GATE U7705 ( .I1(n6703), .I2(n6702), .O(n7213) );
  NAND_GATE U7706 ( .I1(n6712), .I2(n7213), .O(n7215) );
  NAND3_GATE U7707 ( .I1(n6705), .I2(n7204), .I3(n674), .O(n7202) );
  INV_GATE U7708 ( .I1(n6705), .O(n6707) );
  NAND_GATE U7709 ( .I1(n6707), .I2(n6706), .O(n6704) );
  NAND_GATE U7710 ( .I1(n7204), .I2(n6704), .O(n6711) );
  NAND_GATE U7711 ( .I1(n6705), .I2(n674), .O(n6708) );
  NAND_GATE U7712 ( .I1(n6708), .I2(n6704), .O(n7205) );
  NAND_GATE U7713 ( .I1(n7200), .I2(n7205), .O(n6709) );
  NAND_GATE U7714 ( .I1(n6711), .I2(n6709), .O(n6710) );
  NAND_GATE U7715 ( .I1(n7202), .I2(n6710), .O(n7216) );
  NAND_GATE U7716 ( .I1(n7213), .I2(n7216), .O(n6715) );
  NAND_GATE U7717 ( .I1(n7200), .I2(n7205), .O(n6714) );
  INV_GATE U7718 ( .I1(n6711), .O(n7201) );
  NAND_GATE U7719 ( .I1(n7202), .I2(n7201), .O(n6713) );
  NAND3_GATE U7720 ( .I1(n6714), .I2(n6713), .I3(n6712), .O(n7214) );
  NAND_GATE U7721 ( .I1(n6717), .I2(n6716), .O(n7372) );
  NAND_GATE U7722 ( .I1(n6724), .I2(n7372), .O(n7378) );
  NAND_GATE U7723 ( .I1(n1343), .I2(n6721), .O(n6718) );
  NAND_GATE U7724 ( .I1(n6719), .I2(n6718), .O(n7369) );
  INV_GATE U7725 ( .I1(n7369), .O(n6720) );
  NAND3_GATE U7726 ( .I1(n7365), .I2(n6719), .I3(n208), .O(n7371) );
  NAND_GATE U7727 ( .I1(n6720), .I2(n7371), .O(n6723) );
  NAND_GATE U7728 ( .I1(n7366), .I2(n6722), .O(n7376) );
  NAND3_GATE U7729 ( .I1(n7372), .I2(n6723), .I3(n7376), .O(n6727) );
  NAND_GATE U7730 ( .I1(n6724), .I2(n6723), .O(n6725) );
  INV_GATE U7731 ( .I1(n6725), .O(n7377) );
  NAND_GATE U7732 ( .I1(n7388), .I2(n7389), .O(n6728) );
  NAND_GATE U7733 ( .I1(n7387), .I2(n6728), .O(n6729) );
  NAND_GATE U7734 ( .I1(n6730), .I2(n6729), .O(n7401) );
  NAND_GATE U7735 ( .I1(n6740), .I2(n7401), .O(n7398) );
  NAND_GATE U7736 ( .I1(n6734), .I2(n6743), .O(n6736) );
  NAND_GATE U7737 ( .I1(n6742), .I2(n6741), .O(n6733) );
  NAND_GATE U7738 ( .I1(n1247), .I2(n6731), .O(n6743) );
  NAND3_GATE U7739 ( .I1(n6736), .I2(n6733), .I3(n6732), .O(n6735) );
  NAND3_GATE U7740 ( .I1(n6742), .I2(n6734), .I3(n6741), .O(n6737) );
  NAND_GATE U7741 ( .I1(n6735), .I2(n6737), .O(n7402) );
  NAND_GATE U7742 ( .I1(n7401), .I2(n7402), .O(n6747) );
  INV_GATE U7743 ( .I1(n6736), .O(n6738) );
  NAND_GATE U7744 ( .I1(n6738), .I2(n6737), .O(n6739) );
  AND_GATE U7745 ( .I1(n6740), .I2(n6739), .O(n7397) );
  NAND_GATE U7746 ( .I1(n6743), .I2(n6733), .O(n6744) );
  NAND_GATE U7747 ( .I1(n6745), .I2(n6744), .O(n7396) );
  NAND_GATE U7748 ( .I1(n7397), .I2(n7396), .O(n6746) );
  NAND_GATE U7749 ( .I1(n7165), .I2(n7174), .O(n7431) );
  NAND3_GATE U7750 ( .I1(n6751), .I2(n6752), .I3(n6748), .O(n7168) );
  INV_GATE U7751 ( .I1(n6752), .O(n6749) );
  NAND3_GATE U7752 ( .I1(n6750), .I2(n6749), .I3(n6748), .O(n7169) );
  NAND3_GATE U7753 ( .I1(n7167), .I2(n6752), .I3(n6751), .O(n7172) );
  NAND3_GATE U7754 ( .I1(n7174), .I2(n989), .I3(n7164), .O(n7432) );
  NAND3_GATE U7755 ( .I1(n7167), .I2(n7166), .I3(n7172), .O(n7164) );
  NAND3_GATE U7756 ( .I1(n7165), .I2(n7164), .I3(n989), .O(n7430) );
  NAND3_GATE U7757 ( .I1(n7431), .I2(n7432), .I3(n7430), .O(n7436) );
  NAND_GATE U7758 ( .I1(n6757), .I2(n7436), .O(n7416) );
  NAND_GATE U7759 ( .I1(n6754), .I2(n7426), .O(n7420) );
  NAND_GATE U7760 ( .I1(n7429), .I2(n209), .O(n6755) );
  NAND3_GATE U7761 ( .I1(n7420), .I2(n7427), .I3(n6755), .O(n6756) );
  NAND_GATE U7762 ( .I1(n7422), .I2(n6756), .O(n7417) );
  NAND_GATE U7763 ( .I1(n6757), .I2(n7417), .O(n7415) );
  NAND_GATE U7764 ( .I1(n7436), .I2(n7417), .O(n6758) );
  NAND3_GATE U7765 ( .I1(n7416), .I2(n7415), .I3(n6758), .O(n7153) );
  NAND_GATE U7766 ( .I1(n7158), .I2(n7153), .O(n7159) );
  NAND3_GATE U7767 ( .I1(n6759), .I2(n6760), .I3(n708), .O(n7147) );
  INV_GATE U7768 ( .I1(n6760), .O(n6761) );
  NAND_GATE U7769 ( .I1(n6759), .I2(n6763), .O(n7146) );
  NAND_GATE U7770 ( .I1(n708), .I2(n6760), .O(n6764) );
  NAND_GATE U7771 ( .I1(n6762), .I2(n6761), .O(n6763) );
  NAND_GATE U7772 ( .I1(n6764), .I2(n6763), .O(n7148) );
  NAND_GATE U7773 ( .I1(n7146), .I2(n7151), .O(n6765) );
  NAND_GATE U7774 ( .I1(n7147), .I2(n6765), .O(n7160) );
  NAND_GATE U7775 ( .I1(n7158), .I2(n7160), .O(n6767) );
  NAND_GATE U7776 ( .I1(n7153), .I2(n7160), .O(n6766) );
  NAND3_GATE U7777 ( .I1(n7159), .I2(n6767), .I3(n6766), .O(n7135) );
  NAND_GATE U7778 ( .I1(n7140), .I2(n7135), .O(n7139) );
  NAND_GATE U7779 ( .I1(n753), .I2(n6771), .O(n6779) );
  NAND_GATE U7780 ( .I1(n6774), .I2(n790), .O(n6769) );
  NAND_GATE U7781 ( .I1(n6770), .I2(n6769), .O(n6777) );
  NAND_GATE U7782 ( .I1(n6772), .I2(n6771), .O(n6776) );
  NAND3_GATE U7783 ( .I1(n6774), .I2(n790), .I3(n6773), .O(n6775) );
  NAND3_GATE U7784 ( .I1(n6777), .I2(n6776), .I3(n6775), .O(n6778) );
  NAND_GATE U7785 ( .I1(n7140), .I2(n7141), .O(n6781) );
  NAND_GATE U7786 ( .I1(n7135), .I2(n7141), .O(n6780) );
  NAND3_GATE U7787 ( .I1(n7139), .I2(n6781), .I3(n6780), .O(n7127) );
  NAND_GATE U7788 ( .I1(n6789), .I2(n7127), .O(n7121) );
  NAND_GATE U7789 ( .I1(n6782), .I2(n6784), .O(n6790) );
  NAND_GATE U7790 ( .I1(n6791), .I2(n6790), .O(n7124) );
  NAND_GATE U7791 ( .I1(n6783), .I2(n1257), .O(n6784) );
  NAND_GATE U7792 ( .I1(n6785), .I2(n6784), .O(n6792) );
  INV_GATE U7793 ( .I1(n6792), .O(n6788) );
  NAND_GATE U7794 ( .I1(n6788), .I2(n6794), .O(n7125) );
  NAND3_GATE U7795 ( .I1(n7124), .I2(n7125), .I3(n6789), .O(n7120) );
  AND_GATE U7796 ( .I1(n7121), .I2(n7120), .O(n6796) );
  NAND_GATE U7797 ( .I1(n6792), .I2(n7124), .O(n6793) );
  NAND_GATE U7798 ( .I1(n6794), .I2(n6793), .O(n7128) );
  NAND_GATE U7799 ( .I1(n7127), .I2(n7128), .O(n6795) );
  NAND_GATE U7800 ( .I1(n6796), .I2(n6795), .O(n7115) );
  NAND_GATE U7801 ( .I1(n6809), .I2(n7115), .O(n7111) );
  OR_GATE U7802 ( .I1(n6801), .I2(n6797), .O(n6808) );
  NAND_GATE U7803 ( .I1(n824), .I2(n6801), .O(n6798) );
  NAND_GATE U7804 ( .I1(n6799), .I2(n6798), .O(n6806) );
  NAND_GATE U7805 ( .I1(n6802), .I2(n6798), .O(n6803) );
  NAND_GATE U7806 ( .I1(n6804), .I2(n6803), .O(n6805) );
  NAND_GATE U7807 ( .I1(n6806), .I2(n6805), .O(n6807) );
  NAND_GATE U7808 ( .I1(n6808), .I2(n6807), .O(n7114) );
  NAND_GATE U7809 ( .I1(n6809), .I2(n7114), .O(n7110) );
  NAND_GATE U7810 ( .I1(n7115), .I2(n7114), .O(n6810) );
  NAND3_GATE U7811 ( .I1(n7111), .I2(n7110), .I3(n6810), .O(n7104) );
  NAND_GATE U7812 ( .I1(n6819), .I2(n7104), .O(n7100) );
  NAND_GATE U7813 ( .I1(n778), .I2(n6817), .O(n6811) );
  INV_GATE U7814 ( .I1(n6817), .O(n6812) );
  NAND_GATE U7815 ( .I1(n6811), .I2(n6814), .O(n6822) );
  NAND_GATE U7816 ( .I1(n6823), .I2(n6822), .O(n6821) );
  NAND_GATE U7817 ( .I1(n6813), .I2(n6812), .O(n6814) );
  NAND_GATE U7818 ( .I1(n6815), .I2(n6814), .O(n6824) );
  INV_GATE U7819 ( .I1(n6824), .O(n6818) );
  NAND_GATE U7820 ( .I1(n6818), .I2(n6826), .O(n6820) );
  NAND3_GATE U7821 ( .I1(n6821), .I2(n6820), .I3(n6819), .O(n7099) );
  NAND_GATE U7822 ( .I1(n6826), .I2(n6825), .O(n7103) );
  NAND_GATE U7823 ( .I1(n7104), .I2(n7103), .O(n6827) );
  NAND3_GATE U7824 ( .I1(n7100), .I2(n7099), .I3(n6827), .O(n7093) );
  NAND_GATE U7825 ( .I1(n6835), .I2(n7093), .O(n7089) );
  NAND_GATE U7826 ( .I1(n6828), .I2(n618), .O(n6830) );
  NAND_GATE U7827 ( .I1(n6831), .I2(n789), .O(n6829) );
  NAND_GATE U7828 ( .I1(n6830), .I2(n6829), .O(n6838) );
  NAND_GATE U7829 ( .I1(n6839), .I2(n6838), .O(n6837) );
  NAND_GATE U7830 ( .I1(n6832), .I2(n6829), .O(n6840) );
  INV_GATE U7831 ( .I1(n6840), .O(n6834) );
  NAND_GATE U7832 ( .I1(n6834), .I2(n6842), .O(n6836) );
  NAND3_GATE U7833 ( .I1(n6837), .I2(n6836), .I3(n6835), .O(n7088) );
  NAND_GATE U7834 ( .I1(n6840), .I2(n6837), .O(n6841) );
  NAND_GATE U7835 ( .I1(n6842), .I2(n6841), .O(n7092) );
  NAND_GATE U7836 ( .I1(n7093), .I2(n7092), .O(n6843) );
  NAND3_GATE U7837 ( .I1(n7089), .I2(n7088), .I3(n6843), .O(n7082) );
  NAND_GATE U7838 ( .I1(n6852), .I2(n7082), .O(n7078) );
  NAND_GATE U7839 ( .I1(n6844), .I2(n6851), .O(n6846) );
  INV_GATE U7840 ( .I1(n6851), .O(n6847) );
  NAND_GATE U7841 ( .I1(n6848), .I2(n6847), .O(n6845) );
  NAND_GATE U7842 ( .I1(n6846), .I2(n6845), .O(n6855) );
  NAND_GATE U7843 ( .I1(n6856), .I2(n6855), .O(n6854) );
  NAND_GATE U7844 ( .I1(n6849), .I2(n6845), .O(n6857) );
  NAND3_GATE U7845 ( .I1(n6854), .I2(n6853), .I3(n6852), .O(n7077) );
  NAND_GATE U7846 ( .I1(n7082), .I2(n7081), .O(n6859) );
  NAND3_GATE U7847 ( .I1(n7078), .I2(n7077), .I3(n6859), .O(n7071) );
  NAND_GATE U7848 ( .I1(n6868), .I2(n7071), .O(n7067) );
  INV_GATE U7849 ( .I1(n6867), .O(n6860) );
  NAND_GATE U7850 ( .I1(n6861), .I2(n6860), .O(n6864) );
  NAND_GATE U7851 ( .I1(n6862), .I2(n6867), .O(n6863) );
  NAND_GATE U7852 ( .I1(n6864), .I2(n6863), .O(n6871) );
  NAND_GATE U7853 ( .I1(n6872), .I2(n6871), .O(n6870) );
  NAND_GATE U7854 ( .I1(n6865), .I2(n6864), .O(n6873) );
  NAND3_GATE U7855 ( .I1(n6870), .I2(n6869), .I3(n6868), .O(n7066) );
  NAND_GATE U7856 ( .I1(n7071), .I2(n7070), .O(n6875) );
  NAND3_GATE U7857 ( .I1(n7067), .I2(n7066), .I3(n6875), .O(n7060) );
  NAND_GATE U7858 ( .I1(n6884), .I2(n7060), .O(n7056) );
  NAND_GATE U7859 ( .I1(n6877), .I2(n6882), .O(n6878) );
  NAND_GATE U7860 ( .I1(n6879), .I2(n6878), .O(n6887) );
  NAND_GATE U7861 ( .I1(n6888), .I2(n6887), .O(n6886) );
  NAND_GATE U7862 ( .I1(n6880), .I2(n6879), .O(n6889) );
  INV_GATE U7863 ( .I1(n6889), .O(n6883) );
  NAND_GATE U7864 ( .I1(n6883), .I2(n6891), .O(n6885) );
  NAND3_GATE U7865 ( .I1(n6886), .I2(n6885), .I3(n6884), .O(n7055) );
  NAND_GATE U7866 ( .I1(n6889), .I2(n6886), .O(n6890) );
  NAND_GATE U7867 ( .I1(n6891), .I2(n6890), .O(n7059) );
  NAND_GATE U7868 ( .I1(n7060), .I2(n7059), .O(n6892) );
  NAND3_GATE U7869 ( .I1(n7056), .I2(n7055), .I3(n6892), .O(n7049) );
  NAND_GATE U7870 ( .I1(n6901), .I2(n7049), .O(n7045) );
  NAND_GATE U7871 ( .I1(n6894), .I2(n6899), .O(n6895) );
  NAND_GATE U7872 ( .I1(n6896), .I2(n6895), .O(n6904) );
  NAND_GATE U7873 ( .I1(n6905), .I2(n6904), .O(n6903) );
  NAND_GATE U7874 ( .I1(n6897), .I2(n6896), .O(n6906) );
  INV_GATE U7875 ( .I1(n6906), .O(n6900) );
  NAND_GATE U7876 ( .I1(n6900), .I2(n6908), .O(n6902) );
  NAND3_GATE U7877 ( .I1(n6903), .I2(n6902), .I3(n6901), .O(n7044) );
  NAND_GATE U7878 ( .I1(n6906), .I2(n6903), .O(n6907) );
  NAND_GATE U7879 ( .I1(n6908), .I2(n6907), .O(n7048) );
  NAND_GATE U7880 ( .I1(n7049), .I2(n7048), .O(n6909) );
  NAND3_GATE U7881 ( .I1(n7045), .I2(n7044), .I3(n6909), .O(n7038) );
  NAND_GATE U7882 ( .I1(n6918), .I2(n7038), .O(n7032) );
  NAND_GATE U7883 ( .I1(n6911), .I2(n6916), .O(n6912) );
  NAND_GATE U7884 ( .I1(n6913), .I2(n6912), .O(n6920) );
  NAND_GATE U7885 ( .I1(n6914), .I2(n6913), .O(n6923) );
  INV_GATE U7886 ( .I1(n6923), .O(n6917) );
  NAND_GATE U7887 ( .I1(n6917), .I2(n6925), .O(n6919) );
  NAND3_GATE U7888 ( .I1(n6922), .I2(n6919), .I3(n6918), .O(n7031) );
  NAND_GATE U7889 ( .I1(n6921), .I2(n6920), .O(n6922) );
  NAND_GATE U7890 ( .I1(n6923), .I2(n6922), .O(n6924) );
  NAND_GATE U7891 ( .I1(n6925), .I2(n6924), .O(n7036) );
  NAND_GATE U7892 ( .I1(n7038), .I2(n7036), .O(n6926) );
  NAND3_GATE U7893 ( .I1(n7032), .I2(n7031), .I3(n6926), .O(n7020) );
  NAND_GATE U7894 ( .I1(n6935), .I2(n7020), .O(n7024) );
  NAND_GATE U7895 ( .I1(n6928), .I2(n6933), .O(n6929) );
  NAND_GATE U7896 ( .I1(n6930), .I2(n6929), .O(n6937) );
  NAND_GATE U7897 ( .I1(n6931), .I2(n6930), .O(n6940) );
  INV_GATE U7898 ( .I1(n6940), .O(n6934) );
  NAND_GATE U7899 ( .I1(n6934), .I2(n6942), .O(n6936) );
  NAND3_GATE U7900 ( .I1(n6939), .I2(n6936), .I3(n6935), .O(n7028) );
  NAND_GATE U7901 ( .I1(n6938), .I2(n6937), .O(n6939) );
  NAND_GATE U7902 ( .I1(n6940), .I2(n6939), .O(n6941) );
  NAND_GATE U7903 ( .I1(n6942), .I2(n6941), .O(n7025) );
  NAND_GATE U7904 ( .I1(n7020), .I2(n7025), .O(n6943) );
  NAND3_GATE U7905 ( .I1(n7024), .I2(n7028), .I3(n6943), .O(n7009) );
  NAND_GATE U7906 ( .I1(n6952), .I2(n7009), .O(n7013) );
  INV_GATE U7907 ( .I1(n6951), .O(n6944) );
  NAND_GATE U7908 ( .I1(n6945), .I2(n6944), .O(n6948) );
  NAND_GATE U7909 ( .I1(n6946), .I2(n6951), .O(n6947) );
  NAND_GATE U7910 ( .I1(n6948), .I2(n6947), .O(n7005) );
  NAND_GATE U7911 ( .I1(n7006), .I2(n7005), .O(n6953) );
  NAND_GATE U7912 ( .I1(n6949), .I2(n6948), .O(n6955) );
  INV_GATE U7913 ( .I1(n6955), .O(n7004) );
  NAND3_GATE U7914 ( .I1(n6953), .I2(n7007), .I3(n6952), .O(n7017) );
  NAND_GATE U7915 ( .I1(n7006), .I2(n7005), .O(n6954) );
  NAND_GATE U7916 ( .I1(n6955), .I2(n6954), .O(n6956) );
  NAND_GATE U7917 ( .I1(n7003), .I2(n6956), .O(n7014) );
  NAND_GATE U7918 ( .I1(n7009), .I2(n7014), .O(n6957) );
  NAND3_GATE U7919 ( .I1(n7013), .I2(n7017), .I3(n6957), .O(n6997) );
  NAND_GATE U7920 ( .I1(n6966), .I2(n6997), .O(n6986) );
  NAND3_GATE U7921 ( .I1(n6960), .I2(n6961), .I3(n6959), .O(n6992) );
  NAND_GATE U7922 ( .I1(n6959), .I2(n6963), .O(n6991) );
  NAND_GATE U7923 ( .I1(n6961), .I2(n6960), .O(n6962) );
  NAND_GATE U7924 ( .I1(n6963), .I2(n6962), .O(n6993) );
  NAND_GATE U7925 ( .I1(n6994), .I2(n6993), .O(n6964) );
  NAND_GATE U7926 ( .I1(n6991), .I2(n6964), .O(n6965) );
  NAND_GATE U7927 ( .I1(n6992), .I2(n6965), .O(n6989) );
  NAND_GATE U7928 ( .I1(n6966), .I2(n6989), .O(n6985) );
  NAND_GATE U7929 ( .I1(n6997), .I2(n6989), .O(n6967) );
  NAND3_GATE U7930 ( .I1(n6986), .I2(n6985), .I3(n6967), .O(n15324) );
  INV_GATE U7931 ( .I1(n15324), .O(n6982) );
  INV_GATE U7932 ( .I1(n6968), .O(n6969) );
  NAND_GATE U7933 ( .I1(n6969), .I2(n6972), .O(n6981) );
  NAND_GATE U7934 ( .I1(n6971), .I2(n6975), .O(n6979) );
  NAND_GATE U7935 ( .I1(n6973), .I2(n6972), .O(n6974) );
  NAND_GATE U7936 ( .I1(n6975), .I2(n6974), .O(n6976) );
  NAND_GATE U7937 ( .I1(n6977), .I2(n6976), .O(n6978) );
  NAND_GATE U7938 ( .I1(n6979), .I2(n6978), .O(n6980) );
  NAND_GATE U7939 ( .I1(n6981), .I2(n6980), .O(n15323) );
  NAND_GATE U7940 ( .I1(n6982), .I2(n15323), .O(n6984) );
  NAND_GATE U7941 ( .I1(n6984), .I2(n6983), .O(\A1[48] ) );
  OR_GATE U7942 ( .I1(n6985), .I2(n6997), .O(n6988) );
  OR_GATE U7943 ( .I1(n6989), .I2(n6986), .O(n6987) );
  AND_GATE U7944 ( .I1(n6988), .I2(n6987), .O(n7002) );
  INV_GATE U7945 ( .I1(n6997), .O(n6990) );
  NAND_GATE U7946 ( .I1(n6990), .I2(n6989), .O(n7000) );
  NAND_GATE U7947 ( .I1(n6995), .I2(n6964), .O(n6996) );
  NAND_GATE U7948 ( .I1(n6997), .I2(n6996), .O(n6999) );
  NAND3_GATE U7949 ( .I1(n7000), .I2(n6999), .I3(n6998), .O(n7001) );
  INV_GATE U7950 ( .I1(n7009), .O(n7018) );
  NAND_GATE U7951 ( .I1(n7018), .I2(n7014), .O(n7012) );
  NAND_GATE U7952 ( .I1(n7004), .I2(n7003), .O(n7007) );
  NAND_GATE U7953 ( .I1(n7007), .I2(n6953), .O(n7008) );
  NAND_GATE U7954 ( .I1(n7009), .I2(n7008), .O(n7011) );
  NAND3_GATE U7955 ( .I1(n7012), .I2(n7011), .I3(n7010), .O(n7016) );
  OR_GATE U7956 ( .I1(n7014), .I2(n7013), .O(n7015) );
  NAND_GATE U7957 ( .I1(n7016), .I2(n7015), .O(n7019) );
  NAND_GATE U7958 ( .I1(n1382), .I2(A[31]), .O(n7877) );
  INV_GATE U7959 ( .I1(n7877), .O(n7872) );
  NAND_GATE U7960 ( .I1(n472), .I2(n7872), .O(n7870) );
  NAND_GATE U7961 ( .I1(n7019), .I2(n7877), .O(n7472) );
  NAND_GATE U7962 ( .I1(n278), .I2(n7877), .O(n7471) );
  NAND_GATE U7963 ( .I1(n221), .I2(n7025), .O(n7023) );
  NAND3_GATE U7964 ( .I1(n7023), .I2(n7022), .I3(n7021), .O(n7027) );
  OR_GATE U7965 ( .I1(n7025), .I2(n7024), .O(n7026) );
  NAND_GATE U7966 ( .I1(n7027), .I2(n7026), .O(n7030) );
  INV_GATE U7967 ( .I1(n7028), .O(n7029) );
  INV_GATE U7968 ( .I1(n7856), .O(n7859) );
  NAND_GATE U7969 ( .I1(n1382), .I2(A[30]), .O(n7863) );
  INV_GATE U7970 ( .I1(n7863), .O(n7857) );
  NAND_GATE U7971 ( .I1(n7859), .I2(n7857), .O(n7853) );
  NAND_GATE U7972 ( .I1(n7030), .I2(n7863), .O(n7469) );
  NAND_GATE U7973 ( .I1(n282), .I2(n7863), .O(n7468) );
  OR_GATE U7974 ( .I1(n7031), .I2(n7038), .O(n7034) );
  OR_GATE U7975 ( .I1(n7036), .I2(n7032), .O(n7033) );
  AND_GATE U7976 ( .I1(n7034), .I2(n7033), .O(n7043) );
  INV_GATE U7977 ( .I1(n7038), .O(n7035) );
  NAND_GATE U7978 ( .I1(n7035), .I2(n7036), .O(n7041) );
  INV_GATE U7979 ( .I1(n7036), .O(n7037) );
  NAND_GATE U7980 ( .I1(n7038), .I2(n7037), .O(n7040) );
  NAND3_GATE U7981 ( .I1(n7041), .I2(n7040), .I3(n7039), .O(n7042) );
  NAND_GATE U7982 ( .I1(n7043), .I2(n7042), .O(n7839) );
  INV_GATE U7983 ( .I1(n7839), .O(n7842) );
  NAND_GATE U7984 ( .I1(n1382), .I2(A[29]), .O(n7846) );
  INV_GATE U7985 ( .I1(n7846), .O(n7840) );
  NAND_GATE U7986 ( .I1(n7842), .I2(n7840), .O(n7837) );
  OR_GATE U7987 ( .I1(n7044), .I2(n7049), .O(n7047) );
  OR_GATE U7988 ( .I1(n7048), .I2(n7045), .O(n7046) );
  AND_GATE U7989 ( .I1(n7047), .I2(n7046), .O(n7054) );
  NAND_GATE U7990 ( .I1(n983), .I2(n7048), .O(n7052) );
  NAND3_GATE U7991 ( .I1(n7052), .I2(n7051), .I3(n7050), .O(n7053) );
  NAND_GATE U7992 ( .I1(n7054), .I2(n7053), .O(n7823) );
  INV_GATE U7993 ( .I1(n7823), .O(n7826) );
  NAND_GATE U7994 ( .I1(n1382), .I2(A[28]), .O(n7830) );
  INV_GATE U7995 ( .I1(n7830), .O(n7824) );
  NAND_GATE U7996 ( .I1(n7826), .I2(n7824), .O(n7820) );
  OR_GATE U7997 ( .I1(n7055), .I2(n7060), .O(n7058) );
  OR_GATE U7998 ( .I1(n7059), .I2(n7056), .O(n7057) );
  AND_GATE U7999 ( .I1(n7058), .I2(n7057), .O(n7065) );
  NAND_GATE U8000 ( .I1(n992), .I2(n7059), .O(n7063) );
  NAND3_GATE U8001 ( .I1(n7063), .I2(n7062), .I3(n7061), .O(n7064) );
  NAND_GATE U8002 ( .I1(n7065), .I2(n7064), .O(n7806) );
  NAND_GATE U8003 ( .I1(n1382), .I2(A[27]), .O(n7813) );
  INV_GATE U8004 ( .I1(n7813), .O(n7807) );
  NAND_GATE U8005 ( .I1(n7809), .I2(n7807), .O(n7804) );
  OR_GATE U8006 ( .I1(n7066), .I2(n7071), .O(n7069) );
  OR_GATE U8007 ( .I1(n7070), .I2(n7067), .O(n7068) );
  AND_GATE U8008 ( .I1(n7069), .I2(n7068), .O(n7076) );
  NAND_GATE U8009 ( .I1(n89), .I2(n7070), .O(n7074) );
  NAND3_GATE U8010 ( .I1(n7074), .I2(n7073), .I3(n7072), .O(n7075) );
  NAND_GATE U8011 ( .I1(n7076), .I2(n7075), .O(n7790) );
  NAND_GATE U8012 ( .I1(n1382), .I2(A[26]), .O(n7797) );
  INV_GATE U8013 ( .I1(n7797), .O(n7791) );
  NAND_GATE U8014 ( .I1(n7793), .I2(n7791), .O(n7788) );
  OR_GATE U8015 ( .I1(n7077), .I2(n7082), .O(n7080) );
  OR_GATE U8016 ( .I1(n7081), .I2(n7078), .O(n7079) );
  AND_GATE U8017 ( .I1(n7080), .I2(n7079), .O(n7087) );
  NAND_GATE U8018 ( .I1(n958), .I2(n7081), .O(n7085) );
  NAND3_GATE U8019 ( .I1(n7085), .I2(n7084), .I3(n7083), .O(n7086) );
  NAND_GATE U8020 ( .I1(n7087), .I2(n7086), .O(n7777) );
  NAND_GATE U8021 ( .I1(n1382), .I2(A[25]), .O(n7781) );
  INV_GATE U8022 ( .I1(n7781), .O(n7774) );
  NAND_GATE U8023 ( .I1(n7776), .I2(n7774), .O(n7772) );
  OR_GATE U8024 ( .I1(n7088), .I2(n7093), .O(n7091) );
  OR_GATE U8025 ( .I1(n7092), .I2(n7089), .O(n7090) );
  AND_GATE U8026 ( .I1(n7091), .I2(n7090), .O(n7098) );
  NAND_GATE U8027 ( .I1(n926), .I2(n7092), .O(n7096) );
  NAND3_GATE U8028 ( .I1(n7096), .I2(n7095), .I3(n7094), .O(n7097) );
  NAND_GATE U8029 ( .I1(n7098), .I2(n7097), .O(n7762) );
  NAND_GATE U8030 ( .I1(n1382), .I2(A[24]), .O(n7765) );
  INV_GATE U8031 ( .I1(n7765), .O(n7760) );
  NAND_GATE U8032 ( .I1(n832), .I2(n7760), .O(n7757) );
  OR_GATE U8033 ( .I1(n7099), .I2(n7104), .O(n7102) );
  OR_GATE U8034 ( .I1(n7103), .I2(n7100), .O(n7101) );
  AND_GATE U8035 ( .I1(n7102), .I2(n7101), .O(n7109) );
  NAND_GATE U8036 ( .I1(n925), .I2(n7103), .O(n7107) );
  NAND3_GATE U8037 ( .I1(n7107), .I2(n7106), .I3(n7105), .O(n7108) );
  NAND_GATE U8038 ( .I1(n1382), .I2(A[23]), .O(n7750) );
  INV_GATE U8039 ( .I1(n7750), .O(n7743) );
  NAND_GATE U8040 ( .I1(n7745), .I2(n7743), .O(n7740) );
  OR_GATE U8041 ( .I1(n7110), .I2(n7115), .O(n7113) );
  OR_GATE U8042 ( .I1(n7114), .I2(n7111), .O(n7112) );
  NAND_GATE U8043 ( .I1(n959), .I2(n7114), .O(n7118) );
  NAND3_GATE U8044 ( .I1(n7118), .I2(n7117), .I3(n7116), .O(n7119) );
  INV_GATE U8045 ( .I1(n7734), .O(n7731) );
  NAND_GATE U8046 ( .I1(n1382), .I2(A[22]), .O(n7732) );
  NAND_GATE U8047 ( .I1(n1382), .I2(A[21]), .O(n7991) );
  INV_GATE U8048 ( .I1(n7991), .O(n7722) );
  OR_GATE U8049 ( .I1(n7120), .I2(n7127), .O(n7123) );
  OR_GATE U8050 ( .I1(n7128), .I2(n7121), .O(n7122) );
  AND_GATE U8051 ( .I1(n7123), .I2(n7122), .O(n7134) );
  NAND_GATE U8052 ( .I1(n7125), .I2(n7124), .O(n7126) );
  NAND_GATE U8053 ( .I1(n7127), .I2(n7126), .O(n7131) );
  INV_GATE U8054 ( .I1(n7127), .O(n7129) );
  NAND_GATE U8055 ( .I1(n7129), .I2(n7128), .O(n7130) );
  NAND3_GATE U8056 ( .I1(n7132), .I2(n7131), .I3(n7130), .O(n7133) );
  NAND_GATE U8057 ( .I1(n7722), .I2(n858), .O(n7452) );
  NAND_GATE U8058 ( .I1(n1382), .I2(A[20]), .O(n8009) );
  INV_GATE U8059 ( .I1(n8009), .O(n7715) );
  INV_GATE U8060 ( .I1(n7135), .O(n7142) );
  NAND_GATE U8061 ( .I1(n7135), .I2(n631), .O(n7137) );
  NAND3_GATE U8062 ( .I1(n7138), .I2(n7137), .I3(n7136), .O(n7145) );
  OR_GATE U8063 ( .I1(n7141), .I2(n7139), .O(n7144) );
  NAND3_GATE U8064 ( .I1(n7142), .I2(n7141), .I3(n7140), .O(n7143) );
  NAND3_GATE U8065 ( .I1(n7145), .I2(n7144), .I3(n7143), .O(n7718) );
  INV_GATE U8066 ( .I1(n7718), .O(n7717) );
  NAND_GATE U8067 ( .I1(n7715), .I2(n7717), .O(n7449) );
  NAND_GATE U8068 ( .I1(n1382), .I2(A[19]), .O(n8022) );
  INV_GATE U8069 ( .I1(n8022), .O(n7481) );
  INV_GATE U8070 ( .I1(n7153), .O(n7157) );
  NAND_GATE U8071 ( .I1(n7149), .I2(n7148), .O(n7151) );
  NAND3_GATE U8072 ( .I1(n7150), .I2(n7157), .I3(n7151), .O(n7156) );
  NAND_GATE U8073 ( .I1(n7151), .I2(n7150), .O(n7152) );
  NAND_GATE U8074 ( .I1(n7153), .I2(n7152), .O(n7155) );
  NAND3_GATE U8075 ( .I1(n7156), .I2(n7155), .I3(n7154), .O(n7163) );
  NAND3_GATE U8076 ( .I1(n7158), .I2(n7157), .I3(n7160), .O(n7162) );
  OR_GATE U8077 ( .I1(n7160), .I2(n7159), .O(n7161) );
  NAND_GATE U8078 ( .I1(n7481), .I2(n733), .O(n7446) );
  NAND_GATE U8079 ( .I1(n1382), .I2(A[18]), .O(n8045) );
  INV_GATE U8080 ( .I1(n8045), .O(n7703) );
  NAND_GATE U8081 ( .I1(n1382), .I2(A[17]), .O(n7695) );
  INV_GATE U8082 ( .I1(n7695), .O(n7483) );
  NAND4_GATE U8083 ( .I1(n7165), .I2(n7164), .I3(n989), .I4(n184), .O(n7180)
         );
  NAND_GATE U8084 ( .I1(n7167), .I2(n7166), .O(n7170) );
  NAND3_GATE U8085 ( .I1(n7170), .I2(n7169), .I3(n7168), .O(n7171) );
  NAND_GATE U8086 ( .I1(n7172), .I2(n7171), .O(n7173) );
  OR_GATE U8087 ( .I1(n7173), .I2(n7431), .O(n7179) );
  NAND_GATE U8088 ( .I1(n184), .I2(n7173), .O(n7176) );
  NAND3_GATE U8089 ( .I1(n7177), .I2(n7176), .I3(n7175), .O(n7178) );
  NAND3_GATE U8090 ( .I1(n7180), .I2(n7179), .I3(n7178), .O(n7696) );
  INV_GATE U8091 ( .I1(n7696), .O(n7694) );
  NAND_GATE U8092 ( .I1(n7483), .I2(n7694), .O(n7414) );
  NAND_GATE U8093 ( .I1(n7181), .I2(n7183), .O(n7392) );
  INV_GATE U8094 ( .I1(n7392), .O(n7182) );
  NAND3_GATE U8095 ( .I1(n7387), .I2(n816), .I3(n7181), .O(n7394) );
  NAND_GATE U8096 ( .I1(n7182), .I2(n7394), .O(n7186) );
  NAND_GATE U8097 ( .I1(n7389), .I2(n1358), .O(n7183) );
  NAND_GATE U8098 ( .I1(n7391), .I2(n7183), .O(n7184) );
  NAND_GATE U8099 ( .I1(n7388), .I2(n7184), .O(n7185) );
  NAND_GATE U8100 ( .I1(n1382), .I2(A[15]), .O(n7499) );
  INV_GATE U8101 ( .I1(n7499), .O(n7386) );
  NAND3_GATE U8102 ( .I1(n7186), .I2(n7185), .I3(n7386), .O(n7502) );
  NAND3_GATE U8103 ( .I1(n7187), .I2(n7189), .I3(n7188), .O(n7197) );
  NAND3_GATE U8104 ( .I1(n7190), .I2(n1290), .I3(n7187), .O(n7196) );
  AND_GATE U8105 ( .I1(n7197), .I2(n7196), .O(n7192) );
  NAND3_GATE U8106 ( .I1(n7189), .I2(n7188), .I3(n7194), .O(n7199) );
  NAND_GATE U8107 ( .I1(n7190), .I2(n1290), .O(n7193) );
  NAND3_GATE U8108 ( .I1(n7199), .I2(n7193), .I3(n7194), .O(n7191) );
  NAND_GATE U8109 ( .I1(n1382), .I2(A[13]), .O(n7675) );
  INV_GATE U8110 ( .I1(n7675), .O(n7363) );
  NAND3_GATE U8111 ( .I1(n7192), .I2(n7191), .I3(n7363), .O(n7667) );
  NAND_GATE U8112 ( .I1(n7194), .I2(n7193), .O(n7195) );
  NAND3_GATE U8113 ( .I1(n7197), .I2(n7196), .I3(n7195), .O(n7198) );
  NAND_GATE U8114 ( .I1(n7199), .I2(n7198), .O(n7672) );
  NAND_GATE U8115 ( .I1(n1382), .I2(A[12]), .O(n7507) );
  INV_GATE U8116 ( .I1(n7507), .O(n7514) );
  INV_GATE U8117 ( .I1(n7213), .O(n7203) );
  NAND3_GATE U8118 ( .I1(n7203), .I2(n6714), .I3(n7206), .O(n7212) );
  NAND_GATE U8119 ( .I1(n7204), .I2(n7206), .O(n7209) );
  INV_GATE U8120 ( .I1(n7205), .O(n7207) );
  NAND_GATE U8121 ( .I1(n7207), .I2(n7206), .O(n7208) );
  NAND3_GATE U8122 ( .I1(n7213), .I2(n7209), .I3(n7208), .O(n7211) );
  NAND3_GATE U8123 ( .I1(n7212), .I2(n7211), .I3(n7210), .O(n7219) );
  OR_GATE U8124 ( .I1(n7214), .I2(n7213), .O(n7218) );
  OR_GATE U8125 ( .I1(n7216), .I2(n7215), .O(n7217) );
  NAND3_GATE U8126 ( .I1(n7219), .I2(n7218), .I3(n7217), .O(n7510) );
  NAND_GATE U8127 ( .I1(n7514), .I2(n766), .O(n7362) );
  NAND_GATE U8128 ( .I1(n1382), .I2(A[11]), .O(n7657) );
  INV_GATE U8129 ( .I1(n7657), .O(n7358) );
  OR_GATE U8130 ( .I1(n7224), .I2(n7220), .O(n7223) );
  OR_GATE U8131 ( .I1(n7221), .I2(n7226), .O(n7222) );
  AND_GATE U8132 ( .I1(n7223), .I2(n7222), .O(n7231) );
  NAND_GATE U8133 ( .I1(n575), .I2(n7224), .O(n7228) );
  INV_GATE U8134 ( .I1(n7224), .O(n7225) );
  NAND_GATE U8135 ( .I1(n7226), .I2(n7225), .O(n7227) );
  NAND3_GATE U8136 ( .I1(n7229), .I2(n7228), .I3(n7227), .O(n7230) );
  NAND_GATE U8137 ( .I1(n7231), .I2(n7230), .O(n7633) );
  NAND_GATE U8138 ( .I1(n1382), .I2(A[10]), .O(n7637) );
  INV_GATE U8139 ( .I1(n7637), .O(n7631) );
  NAND_GATE U8140 ( .I1(n1330), .I2(n7631), .O(n7640) );
  NAND_GATE U8141 ( .I1(n1382), .I2(A[9]), .O(n7520) );
  INV_GATE U8142 ( .I1(n7520), .O(n7346) );
  NAND_GATE U8143 ( .I1(n7236), .I2(n1359), .O(n7232) );
  NAND_GATE U8144 ( .I1(n7233), .I2(n7232), .O(n7239) );
  NAND_GATE U8145 ( .I1(n7234), .I2(n7241), .O(n7238) );
  NAND3_GATE U8146 ( .I1(n7236), .I2(n1359), .I3(n7235), .O(n7237) );
  NAND3_GATE U8147 ( .I1(n7239), .I2(n7238), .I3(n7237), .O(n7243) );
  NAND_GATE U8148 ( .I1(n7243), .I2(n7242), .O(n7523) );
  NAND_GATE U8149 ( .I1(n7346), .I2(n7523), .O(n7525) );
  NAND_GATE U8150 ( .I1(n1382), .I2(A[8]), .O(n7619) );
  INV_GATE U8151 ( .I1(n7246), .O(n7244) );
  NAND3_GATE U8152 ( .I1(n7253), .I2(n7244), .I3(n7245), .O(n7262) );
  INV_GATE U8153 ( .I1(n7253), .O(n7254) );
  NAND3_GATE U8154 ( .I1(n7246), .I2(n7254), .I3(n7245), .O(n7261) );
  NAND_GATE U8155 ( .I1(n7248), .I2(n7247), .O(n7256) );
  INV_GATE U8156 ( .I1(n7249), .O(n7250) );
  NAND_GATE U8157 ( .I1(n7251), .I2(n7250), .O(n7255) );
  NAND_GATE U8158 ( .I1(n7256), .I2(n7255), .O(n7252) );
  NAND_GATE U8159 ( .I1(n7253), .I2(n7252), .O(n7259) );
  NAND3_GATE U8160 ( .I1(n7256), .I2(n7255), .I3(n7254), .O(n7258) );
  NAND3_GATE U8161 ( .I1(n7259), .I2(n7258), .I3(n7257), .O(n7260) );
  NAND3_GATE U8162 ( .I1(n7262), .I2(n7261), .I3(n7260), .O(n7620) );
  NAND_GATE U8163 ( .I1(n1041), .I2(n7269), .O(n7265) );
  NAND3_GATE U8164 ( .I1(n7265), .I2(n7264), .I3(n7263), .O(n7272) );
  OR_GATE U8165 ( .I1(n7267), .I2(n7266), .O(n7271) );
  OR_GATE U8166 ( .I1(n7269), .I2(n7268), .O(n7270) );
  NAND3_GATE U8167 ( .I1(n7272), .I2(n7271), .I3(n7270), .O(n7608) );
  INV_GATE U8168 ( .I1(n7608), .O(n7610) );
  NAND_GATE U8169 ( .I1(n1382), .I2(A[6]), .O(n7611) );
  INV_GATE U8170 ( .I1(n7611), .O(n7607) );
  NAND_GATE U8171 ( .I1(n7610), .I2(n7607), .O(n7605) );
  NAND_GATE U8172 ( .I1(n1382), .I2(A[5]), .O(n7546) );
  INV_GATE U8173 ( .I1(n7546), .O(n7325) );
  OR_GATE U8174 ( .I1(n7278), .I2(n7274), .O(n7275) );
  AND_GATE U8175 ( .I1(n7276), .I2(n7275), .O(n7284) );
  INV_GATE U8176 ( .I1(n7279), .O(n7277) );
  NAND_GATE U8177 ( .I1(n7277), .I2(n7278), .O(n7282) );
  NAND_GATE U8178 ( .I1(n7279), .I2(n1288), .O(n7281) );
  NAND3_GATE U8179 ( .I1(n7282), .I2(n7281), .I3(n7280), .O(n7283) );
  NAND_GATE U8180 ( .I1(n7284), .I2(n7283), .O(n7589) );
  INV_GATE U8181 ( .I1(n7589), .O(n7592) );
  NAND_GATE U8182 ( .I1(n1382), .I2(A[4]), .O(n7596) );
  INV_GATE U8183 ( .I1(n7596), .O(n7590) );
  NAND_GATE U8184 ( .I1(n7592), .I2(n7590), .O(n7587) );
  NAND_GATE U8185 ( .I1(n1382), .I2(A[3]), .O(n7557) );
  INV_GATE U8186 ( .I1(n7557), .O(n7307) );
  NAND_GATE U8187 ( .I1(n1382), .I2(A[2]), .O(n7578) );
  INV_GATE U8188 ( .I1(n7578), .O(n7572) );
  NAND_GATE U8189 ( .I1(n1384), .I2(A[0]), .O(n7285) );
  NAND_GATE U8190 ( .I1(n14781), .I2(n7285), .O(n7286) );
  NAND_GATE U8191 ( .I1(B[19]), .I2(n7286), .O(n7290) );
  NAND_GATE U8192 ( .I1(n1385), .I2(A[1]), .O(n7287) );
  NAND_GATE U8193 ( .I1(n14784), .I2(n7287), .O(n7288) );
  NAND_GATE U8194 ( .I1(B[18]), .I2(n7288), .O(n7289) );
  NAND_GATE U8195 ( .I1(n7290), .I2(n7289), .O(n7574) );
  NAND_GATE U8196 ( .I1(n7572), .I2(n7574), .O(n7570) );
  NAND3_GATE U8197 ( .I1(n1382), .I2(B[18]), .I3(n1196), .O(n7571) );
  INV_GATE U8198 ( .I1(n7571), .O(n7573) );
  NAND_GATE U8199 ( .I1(n7578), .I2(n649), .O(n7291) );
  NAND_GATE U8200 ( .I1(n7573), .I2(n7291), .O(n7292) );
  NAND_GATE U8201 ( .I1(n7570), .I2(n7292), .O(n7556) );
  NAND_GATE U8202 ( .I1(n7307), .I2(n7556), .O(n7552) );
  OR_GATE U8203 ( .I1(n7294), .I2(n7293), .O(n7306) );
  NAND_GATE U8204 ( .I1(n7295), .I2(n7294), .O(n7300) );
  NAND_GATE U8205 ( .I1(n7296), .I2(n7300), .O(n7304) );
  NAND_GATE U8206 ( .I1(n7298), .I2(n7297), .O(n7299) );
  NAND_GATE U8207 ( .I1(n7300), .I2(n7299), .O(n7301) );
  NAND_GATE U8208 ( .I1(n7302), .I2(n7301), .O(n7303) );
  NAND_GATE U8209 ( .I1(n7304), .I2(n7303), .O(n7305) );
  NAND_GATE U8210 ( .I1(n7306), .I2(n7305), .O(n7555) );
  NAND_GATE U8211 ( .I1(n7556), .I2(n7555), .O(n7308) );
  NAND_GATE U8212 ( .I1(n7307), .I2(n7555), .O(n7551) );
  NAND3_GATE U8213 ( .I1(n7552), .I2(n7308), .I3(n7551), .O(n7591) );
  NAND_GATE U8214 ( .I1(n7589), .I2(n7596), .O(n7309) );
  NAND_GATE U8215 ( .I1(n7591), .I2(n7309), .O(n7310) );
  NAND_GATE U8216 ( .I1(n7587), .I2(n7310), .O(n7545) );
  NAND_GATE U8217 ( .I1(n7325), .I2(n7545), .O(n7541) );
  INV_GATE U8218 ( .I1(n7311), .O(n7312) );
  NAND_GATE U8219 ( .I1(n7312), .I2(n7316), .O(n7324) );
  INV_GATE U8220 ( .I1(n7316), .O(n7313) );
  NAND_GATE U8221 ( .I1(n7314), .I2(n7313), .O(n7318) );
  NAND_GATE U8222 ( .I1(n7315), .I2(n7318), .O(n7322) );
  NAND_GATE U8223 ( .I1(n553), .I2(n7316), .O(n7317) );
  NAND_GATE U8224 ( .I1(n7318), .I2(n7317), .O(n7319) );
  NAND_GATE U8225 ( .I1(n7320), .I2(n7319), .O(n7321) );
  NAND_GATE U8226 ( .I1(n7322), .I2(n7321), .O(n7323) );
  NAND_GATE U8227 ( .I1(n7324), .I2(n7323), .O(n7544) );
  NAND_GATE U8228 ( .I1(n7545), .I2(n7544), .O(n7326) );
  NAND_GATE U8229 ( .I1(n7325), .I2(n7544), .O(n7540) );
  NAND3_GATE U8230 ( .I1(n7541), .I2(n7326), .I3(n7540), .O(n7609) );
  NAND_GATE U8231 ( .I1(n7608), .I2(n7611), .O(n7327) );
  NAND_GATE U8232 ( .I1(n7609), .I2(n7327), .O(n7328) );
  NAND_GATE U8233 ( .I1(n7605), .I2(n7328), .O(n7533) );
  INV_GATE U8234 ( .I1(n7340), .O(n7334) );
  NAND3_GATE U8235 ( .I1(n7331), .I2(n7330), .I3(n7329), .O(n7335) );
  NAND_GATE U8236 ( .I1(n7334), .I2(n7335), .O(n7332) );
  NAND_GATE U8237 ( .I1(n7339), .I2(n7332), .O(n7338) );
  NAND3_GATE U8238 ( .I1(n7334), .I2(n7335), .I3(n7333), .O(n7337) );
  NAND_GATE U8239 ( .I1(n7340), .I2(n1229), .O(n7336) );
  NAND3_GATE U8240 ( .I1(n7338), .I2(n7337), .I3(n7336), .O(n7342) );
  NAND3_GATE U8241 ( .I1(n7340), .I2(n1229), .I3(n7339), .O(n7341) );
  NAND_GATE U8242 ( .I1(n7342), .I2(n7341), .O(n7536) );
  NAND_GATE U8243 ( .I1(n7533), .I2(n7536), .O(n7344) );
  NAND_GATE U8244 ( .I1(n1382), .I2(A[7]), .O(n7532) );
  INV_GATE U8245 ( .I1(n7532), .O(n7343) );
  NAND_GATE U8246 ( .I1(n7343), .I2(n7536), .O(n7534) );
  NAND_GATE U8247 ( .I1(n7343), .I2(n7533), .O(n7535) );
  NAND_GATE U8248 ( .I1(n7619), .I2(n7620), .O(n7345) );
  NAND_GATE U8249 ( .I1(n7523), .I2(n7526), .O(n7347) );
  NAND_GATE U8250 ( .I1(n7346), .I2(n7526), .O(n7524) );
  NAND3_GATE U8251 ( .I1(n7525), .I2(n7347), .I3(n7524), .O(n7641) );
  NAND_GATE U8252 ( .I1(n7633), .I2(n7637), .O(n7348) );
  NAND_GATE U8253 ( .I1(n7641), .I2(n7348), .O(n7349) );
  NAND_GATE U8254 ( .I1(n7640), .I2(n7349), .O(n7652) );
  NAND_GATE U8255 ( .I1(n7358), .I2(n7652), .O(n7658) );
  NAND3_GATE U8256 ( .I1(n7354), .I2(n7350), .I3(n7353), .O(n7648) );
  INV_GATE U8257 ( .I1(n7354), .O(n7352) );
  NAND_GATE U8258 ( .I1(n7350), .I2(n7356), .O(n7647) );
  NAND_GATE U8259 ( .I1(n7352), .I2(n7351), .O(n7356) );
  NAND_GATE U8260 ( .I1(n7354), .I2(n7353), .O(n7355) );
  NAND_GATE U8261 ( .I1(n7356), .I2(n7355), .O(n7649) );
  NAND_GATE U8262 ( .I1(n7647), .I2(n7653), .O(n7357) );
  NAND_GATE U8263 ( .I1(n7648), .I2(n7357), .O(n7659) );
  NAND_GATE U8264 ( .I1(n7652), .I2(n7659), .O(n7359) );
  NAND_GATE U8265 ( .I1(n7358), .I2(n7659), .O(n7660) );
  NAND3_GATE U8266 ( .I1(n7658), .I2(n7359), .I3(n7660), .O(n7508) );
  NAND_GATE U8267 ( .I1(n7507), .I2(n7510), .O(n7360) );
  NAND_GATE U8268 ( .I1(n7508), .I2(n7360), .O(n7361) );
  NAND_GATE U8269 ( .I1(n7362), .I2(n7361), .O(n7671) );
  NAND_GATE U8270 ( .I1(n7672), .I2(n7671), .O(n7364) );
  NAND_GATE U8271 ( .I1(n7363), .I2(n7671), .O(n7668) );
  NAND_GATE U8272 ( .I1(n1382), .I2(A[14]), .O(n8254) );
  NAND_GATE U8273 ( .I1(n7365), .I2(n208), .O(n7368) );
  NAND_GATE U8274 ( .I1(n7366), .I2(n1302), .O(n7367) );
  NAND3_GATE U8275 ( .I1(n7369), .I2(n7368), .I3(n7367), .O(n7370) );
  NAND_GATE U8276 ( .I1(n7371), .I2(n7370), .O(n7379) );
  NAND_GATE U8277 ( .I1(n255), .I2(n7379), .O(n7374) );
  NAND_GATE U8278 ( .I1(n7372), .I2(n207), .O(n7373) );
  NAND3_GATE U8279 ( .I1(n7375), .I2(n7374), .I3(n7373), .O(n7382) );
  NAND3_GATE U8280 ( .I1(n7377), .I2(n7376), .I3(n255), .O(n7381) );
  OR_GATE U8281 ( .I1(n7379), .I2(n7378), .O(n7380) );
  NAND3_GATE U8282 ( .I1(n7382), .I2(n7381), .I3(n7380), .O(n7685) );
  NAND_GATE U8283 ( .I1(n8254), .I2(n7685), .O(n7383) );
  NAND_GATE U8284 ( .I1(n7684), .I2(n7383), .O(n7385) );
  INV_GATE U8285 ( .I1(n8254), .O(n7682) );
  INV_GATE U8286 ( .I1(n7685), .O(n7683) );
  NAND_GATE U8287 ( .I1(n7682), .I2(n7683), .O(n7384) );
  NAND_GATE U8288 ( .I1(n7385), .I2(n7384), .O(n7503) );
  NAND_GATE U8289 ( .I1(n7386), .I2(n7503), .O(n7500) );
  NAND_GATE U8290 ( .I1(n816), .I2(n7387), .O(n7391) );
  NAND3_GATE U8291 ( .I1(n7389), .I2(n1358), .I3(n7388), .O(n7390) );
  NAND3_GATE U8292 ( .I1(n7392), .I2(n7391), .I3(n7390), .O(n7393) );
  NAND_GATE U8293 ( .I1(n7503), .I2(n7501), .O(n7395) );
  NAND_GATE U8294 ( .I1(n1382), .I2(A[16]), .O(n7691) );
  INV_GATE U8295 ( .I1(n7401), .O(n7403) );
  NAND3_GATE U8296 ( .I1(n7397), .I2(n7396), .I3(n7403), .O(n7400) );
  OR_GATE U8297 ( .I1(n7402), .I2(n7398), .O(n7399) );
  AND_GATE U8298 ( .I1(n7400), .I2(n7399), .O(n7408) );
  NAND_GATE U8299 ( .I1(n7403), .I2(n7402), .O(n7404) );
  NAND3_GATE U8300 ( .I1(n7406), .I2(n7405), .I3(n7404), .O(n7407) );
  NAND_GATE U8301 ( .I1(n7408), .I2(n7407), .O(n7491) );
  NAND_GATE U8302 ( .I1(n7691), .I2(n7491), .O(n7409) );
  NAND_GATE U8303 ( .I1(n7495), .I2(n7409), .O(n7411) );
  INV_GATE U8304 ( .I1(n7691), .O(n7494) );
  INV_GATE U8305 ( .I1(n7491), .O(n7493) );
  NAND_GATE U8306 ( .I1(n7494), .I2(n7493), .O(n7410) );
  NAND_GATE U8307 ( .I1(n7695), .I2(n7696), .O(n7412) );
  NAND_GATE U8308 ( .I1(n7693), .I2(n7412), .O(n7413) );
  NAND_GATE U8309 ( .I1(n7414), .I2(n7413), .O(n7706) );
  OR_GATE U8310 ( .I1(n7415), .I2(n7436), .O(n7419) );
  OR_GATE U8311 ( .I1(n7417), .I2(n7416), .O(n7418) );
  AND_GATE U8312 ( .I1(n7419), .I2(n7418), .O(n7441) );
  INV_GATE U8313 ( .I1(n7420), .O(n7421) );
  NAND_GATE U8314 ( .I1(n7422), .I2(n7421), .O(n7434) );
  NAND_GATE U8315 ( .I1(n7424), .I2(n7423), .O(n7427) );
  NAND_GATE U8316 ( .I1(n7425), .I2(n827), .O(n7426) );
  NAND_GATE U8317 ( .I1(n7427), .I2(n7426), .O(n7428) );
  NAND_GATE U8318 ( .I1(n7429), .I2(n7428), .O(n7433) );
  NAND5_GATE U8319 ( .I1(n7434), .I2(n7433), .I3(n7432), .I4(n7431), .I5(n7430), .O(n7439) );
  NAND_GATE U8320 ( .I1(n7434), .I2(n7433), .O(n7435) );
  NAND_GATE U8321 ( .I1(n7436), .I2(n7435), .O(n7438) );
  NAND3_GATE U8322 ( .I1(n7439), .I2(n7438), .I3(n7437), .O(n7440) );
  NAND_GATE U8323 ( .I1(n7441), .I2(n7440), .O(n7707) );
  NAND_GATE U8324 ( .I1(n8045), .I2(n596), .O(n7442) );
  NAND_GATE U8325 ( .I1(n7705), .I2(n7442), .O(n7443) );
  NAND_GATE U8326 ( .I1(n7704), .I2(n7443), .O(n7480) );
  NAND_GATE U8327 ( .I1(n8022), .I2(n711), .O(n7444) );
  NAND_GATE U8328 ( .I1(n7480), .I2(n7444), .O(n7445) );
  NAND_GATE U8329 ( .I1(n7446), .I2(n7445), .O(n7716) );
  NAND_GATE U8330 ( .I1(n8009), .I2(n7718), .O(n7447) );
  NAND_GATE U8331 ( .I1(n7716), .I2(n7447), .O(n7448) );
  NAND_GATE U8332 ( .I1(n7449), .I2(n7448), .O(n7723) );
  NAND_GATE U8333 ( .I1(n7723), .I2(n7450), .O(n7451) );
  NAND_GATE U8334 ( .I1(n7452), .I2(n7451), .O(n7730) );
  NAND_GATE U8335 ( .I1(n7734), .I2(n7732), .O(n7453) );
  NAND_GATE U8336 ( .I1(n7747), .I2(n7750), .O(n7454) );
  NAND_GATE U8337 ( .I1(n7744), .I2(n7454), .O(n7455) );
  NAND_GATE U8338 ( .I1(n7740), .I2(n7455), .O(n7761) );
  NAND_GATE U8339 ( .I1(n7762), .I2(n7765), .O(n7456) );
  NAND_GATE U8340 ( .I1(n7761), .I2(n7456), .O(n7457) );
  NAND_GATE U8341 ( .I1(n7757), .I2(n7457), .O(n7775) );
  NAND_GATE U8342 ( .I1(n7777), .I2(n7781), .O(n7458) );
  NAND_GATE U8343 ( .I1(n7775), .I2(n7458), .O(n7459) );
  NAND_GATE U8344 ( .I1(n7772), .I2(n7459), .O(n7792) );
  NAND_GATE U8345 ( .I1(n7790), .I2(n7797), .O(n7460) );
  NAND_GATE U8346 ( .I1(n7792), .I2(n7460), .O(n7461) );
  NAND_GATE U8347 ( .I1(n7788), .I2(n7461), .O(n7808) );
  NAND_GATE U8348 ( .I1(n7806), .I2(n7813), .O(n7462) );
  NAND_GATE U8349 ( .I1(n7808), .I2(n7462), .O(n7463) );
  NAND_GATE U8350 ( .I1(n7804), .I2(n7463), .O(n7825) );
  NAND_GATE U8351 ( .I1(n7823), .I2(n7830), .O(n7464) );
  NAND_GATE U8352 ( .I1(n7825), .I2(n7464), .O(n7465) );
  NAND_GATE U8353 ( .I1(n7820), .I2(n7465), .O(n7841) );
  NAND_GATE U8354 ( .I1(n7839), .I2(n7846), .O(n7466) );
  NAND_GATE U8355 ( .I1(n7841), .I2(n7466), .O(n7467) );
  NAND_GATE U8356 ( .I1(n7837), .I2(n7467), .O(n7858) );
  NAND3_GATE U8357 ( .I1(n7469), .I2(n7468), .I3(n7858), .O(n7470) );
  NAND_GATE U8358 ( .I1(n7853), .I2(n7470), .O(n7873) );
  NAND3_GATE U8359 ( .I1(n7472), .I2(n7471), .I3(n7873), .O(n7473) );
  NAND_GATE U8360 ( .I1(n7870), .I2(n7473), .O(n7474) );
  NAND_GATE U8361 ( .I1(n471), .I2(n7474), .O(n15325) );
  AND_GATE U8362 ( .I1(n15325), .I2(n7475), .O(\A1[47] ) );
  NAND_GATE U8363 ( .I1(B[16]), .I2(A[31]), .O(n7892) );
  INV_GATE U8364 ( .I1(n7892), .O(n7868) );
  NAND_GATE U8365 ( .I1(B[16]), .I2(A[30]), .O(n7903) );
  INV_GATE U8366 ( .I1(n7903), .O(n7851) );
  NAND_GATE U8367 ( .I1(B[16]), .I2(A[29]), .O(n7914) );
  INV_GATE U8368 ( .I1(n7914), .O(n7835) );
  NAND_GATE U8369 ( .I1(B[16]), .I2(A[28]), .O(n7925) );
  INV_GATE U8370 ( .I1(n7925), .O(n7818) );
  NAND_GATE U8371 ( .I1(B[16]), .I2(A[27]), .O(n7935) );
  INV_GATE U8372 ( .I1(n7935), .O(n7802) );
  NAND_GATE U8373 ( .I1(B[16]), .I2(A[26]), .O(n7945) );
  INV_GATE U8374 ( .I1(n7945), .O(n7786) );
  NAND_GATE U8375 ( .I1(B[16]), .I2(A[25]), .O(n7956) );
  INV_GATE U8376 ( .I1(n7956), .O(n7770) );
  NAND_GATE U8377 ( .I1(B[16]), .I2(A[24]), .O(n7967) );
  INV_GATE U8378 ( .I1(n7967), .O(n7755) );
  NAND_GATE U8379 ( .I1(B[16]), .I2(A[23]), .O(n7980) );
  INV_GATE U8380 ( .I1(n7980), .O(n7738) );
  NAND_GATE U8381 ( .I1(B[16]), .I2(A[22]), .O(n7998) );
  INV_GATE U8382 ( .I1(n7998), .O(n7728) );
  NAND_GATE U8383 ( .I1(B[16]), .I2(A[21]), .O(n8005) );
  INV_GATE U8384 ( .I1(n8005), .O(n8014) );
  NAND_GATE U8385 ( .I1(B[16]), .I2(A[20]), .O(n8030) );
  INV_GATE U8386 ( .I1(n8030), .O(n7712) );
  NAND_GATE U8387 ( .I1(n733), .I2(n7480), .O(n7477) );
  NAND_GATE U8388 ( .I1(n7477), .I2(n7476), .O(n8021) );
  NAND_GATE U8389 ( .I1(n8022), .I2(n8021), .O(n7479) );
  NAND_GATE U8390 ( .I1(n711), .I2(n597), .O(n7478) );
  NAND_GATE U8391 ( .I1(n7481), .I2(n7478), .O(n8023) );
  NAND_GATE U8392 ( .I1(n7479), .I2(n8023), .O(n7482) );
  NAND3_GATE U8393 ( .I1(n7481), .I2(n7480), .I3(n733), .O(n8024) );
  NAND_GATE U8394 ( .I1(n7482), .I2(n8024), .O(n8033) );
  NAND_GATE U8395 ( .I1(B[16]), .I2(A[19]), .O(n8048) );
  INV_GATE U8396 ( .I1(n8048), .O(n7710) );
  NAND_GATE U8397 ( .I1(n7483), .I2(n7486), .O(n7698) );
  INV_GATE U8398 ( .I1(n7698), .O(n7484) );
  NAND3_GATE U8399 ( .I1(n7693), .I2(n7694), .I3(n7483), .O(n7700) );
  NAND_GATE U8400 ( .I1(n7484), .I2(n7700), .O(n7489) );
  NAND_GATE U8401 ( .I1(n7696), .I2(n1344), .O(n7486) );
  NAND_GATE U8402 ( .I1(n7694), .I2(n7693), .O(n7485) );
  NAND_GATE U8403 ( .I1(n7486), .I2(n7485), .O(n7487) );
  NAND_GATE U8404 ( .I1(n7695), .I2(n7487), .O(n7488) );
  NAND_GATE U8405 ( .I1(B[16]), .I2(A[18]), .O(n8060) );
  INV_GATE U8406 ( .I1(n8060), .O(n8051) );
  NAND3_GATE U8407 ( .I1(n7489), .I2(n7488), .I3(n8051), .O(n8052) );
  NAND_GATE U8408 ( .I1(B[16]), .I2(A[17]), .O(n8295) );
  INV_GATE U8409 ( .I1(n8295), .O(n7496) );
  NAND_GATE U8410 ( .I1(n7490), .I2(n7492), .O(n7690) );
  NAND_GATE U8411 ( .I1(n260), .I2(n7491), .O(n7492) );
  NAND3_GATE U8412 ( .I1(n7495), .I2(n7494), .I3(n7493), .O(n8285) );
  NAND_GATE U8413 ( .I1(n1214), .I2(n8285), .O(n8292) );
  NAND3_GATE U8414 ( .I1(n7496), .I2(n8282), .I3(n8292), .O(n8287) );
  NAND_GATE U8415 ( .I1(B[16]), .I2(A[16]), .O(n8271) );
  INV_GATE U8416 ( .I1(n8271), .O(n8274) );
  NAND_GATE U8417 ( .I1(n7503), .I2(n679), .O(n7497) );
  NAND3_GATE U8418 ( .I1(n7499), .I2(n7498), .I3(n7497), .O(n7506) );
  OR_GATE U8419 ( .I1(n7501), .I2(n7500), .O(n7505) );
  OR_GATE U8420 ( .I1(n7503), .I2(n7502), .O(n7504) );
  NAND3_GATE U8421 ( .I1(n7506), .I2(n7505), .I3(n7504), .O(n8272) );
  NAND_GATE U8422 ( .I1(n8274), .I2(n1240), .O(n8291) );
  NAND_GATE U8423 ( .I1(B[16]), .I2(A[15]), .O(n8265) );
  INV_GATE U8424 ( .I1(n8265), .O(n7687) );
  NAND3_GATE U8425 ( .I1(n7507), .I2(n7508), .I3(n766), .O(n7517) );
  NAND3_GATE U8426 ( .I1(n7510), .I2(n7509), .I3(n7507), .O(n7516) );
  AND_GATE U8427 ( .I1(n7517), .I2(n7516), .O(n7512) );
  NAND3_GATE U8428 ( .I1(n7508), .I2(n766), .I3(n7514), .O(n7519) );
  NAND_GATE U8429 ( .I1(n7510), .I2(n7509), .O(n7513) );
  NAND3_GATE U8430 ( .I1(n7519), .I2(n7513), .I3(n7514), .O(n7511) );
  NAND_GATE U8431 ( .I1(B[16]), .I2(A[13]), .O(n8071) );
  INV_GATE U8432 ( .I1(n8071), .O(n7665) );
  NAND3_GATE U8433 ( .I1(n7512), .I2(n7511), .I3(n7665), .O(n8072) );
  NAND_GATE U8434 ( .I1(n7514), .I2(n7513), .O(n7515) );
  NAND3_GATE U8435 ( .I1(n7517), .I2(n7516), .I3(n7515), .O(n7518) );
  NAND_GATE U8436 ( .I1(n7519), .I2(n7518), .O(n8074) );
  NAND_GATE U8437 ( .I1(B[16]), .I2(A[11]), .O(n8088) );
  INV_GATE U8438 ( .I1(n8088), .O(n7645) );
  NAND_GATE U8439 ( .I1(B[16]), .I2(A[10]), .O(n8216) );
  INV_GATE U8440 ( .I1(n8216), .O(n8212) );
  NAND_GATE U8441 ( .I1(n7523), .I2(n524), .O(n7522) );
  NAND_GATE U8442 ( .I1(n1207), .I2(n7526), .O(n7521) );
  NAND3_GATE U8443 ( .I1(n7522), .I2(n7521), .I3(n7520), .O(n7529) );
  OR_GATE U8444 ( .I1(n7524), .I2(n7523), .O(n7528) );
  OR_GATE U8445 ( .I1(n7526), .I2(n7525), .O(n7527) );
  NAND3_GATE U8446 ( .I1(n7529), .I2(n7528), .I3(n7527), .O(n8213) );
  NAND_GATE U8447 ( .I1(n8212), .I2(n1205), .O(n8219) );
  NAND_GATE U8448 ( .I1(B[16]), .I2(A[9]), .O(n8099) );
  INV_GATE U8449 ( .I1(n8099), .O(n7627) );
  NAND_GATE U8450 ( .I1(B[16]), .I2(A[8]), .O(n8435) );
  INV_GATE U8451 ( .I1(n8435), .O(n8200) );
  NAND_GATE U8452 ( .I1(n939), .I2(n7536), .O(n7531) );
  NAND3_GATE U8453 ( .I1(n7532), .I2(n7531), .I3(n7530), .O(n7539) );
  OR_GATE U8454 ( .I1(n7534), .I2(n7533), .O(n7538) );
  OR_GATE U8455 ( .I1(n7536), .I2(n7535), .O(n7537) );
  NAND3_GATE U8456 ( .I1(n7539), .I2(n7538), .I3(n7537), .O(n8204) );
  INV_GATE U8457 ( .I1(n8204), .O(n8202) );
  NAND_GATE U8458 ( .I1(n8200), .I2(n8202), .O(n7618) );
  NAND_GATE U8459 ( .I1(B[16]), .I2(A[7]), .O(n8105) );
  INV_GATE U8460 ( .I1(n8105), .O(n7614) );
  OR_GATE U8461 ( .I1(n7544), .I2(n7541), .O(n7542) );
  AND_GATE U8462 ( .I1(n7543), .I2(n7542), .O(n7550) );
  NAND_GATE U8463 ( .I1(n1066), .I2(n7544), .O(n7548) );
  NAND3_GATE U8464 ( .I1(n7548), .I2(n7547), .I3(n7546), .O(n7549) );
  NAND_GATE U8465 ( .I1(n7550), .I2(n7549), .O(n8184) );
  INV_GATE U8466 ( .I1(n8184), .O(n8187) );
  NAND_GATE U8467 ( .I1(B[16]), .I2(A[6]), .O(n8191) );
  INV_GATE U8468 ( .I1(n8191), .O(n8185) );
  NAND_GATE U8469 ( .I1(n8187), .I2(n8185), .O(n8182) );
  NAND_GATE U8470 ( .I1(B[16]), .I2(A[5]), .O(n8122) );
  INV_GATE U8471 ( .I1(n8122), .O(n7601) );
  OR_GATE U8472 ( .I1(n7551), .I2(n7556), .O(n7554) );
  OR_GATE U8473 ( .I1(n7555), .I2(n7552), .O(n7553) );
  AND_GATE U8474 ( .I1(n7554), .I2(n7553), .O(n7561) );
  NAND_GATE U8475 ( .I1(n1149), .I2(n7555), .O(n7559) );
  NAND3_GATE U8476 ( .I1(n7559), .I2(n7558), .I3(n7557), .O(n7560) );
  NAND_GATE U8477 ( .I1(n7561), .I2(n7560), .O(n8167) );
  NAND_GATE U8478 ( .I1(B[16]), .I2(A[4]), .O(n8173) );
  INV_GATE U8479 ( .I1(n8173), .O(n8168) );
  NAND_GATE U8480 ( .I1(n607), .I2(n8168), .O(n8164) );
  NAND_GATE U8481 ( .I1(B[16]), .I2(A[3]), .O(n8133) );
  INV_GATE U8482 ( .I1(n8133), .O(n7583) );
  NAND_GATE U8483 ( .I1(B[16]), .I2(A[2]), .O(n8155) );
  INV_GATE U8484 ( .I1(n8155), .O(n8149) );
  NAND_GATE U8485 ( .I1(n1383), .I2(A[0]), .O(n7562) );
  NAND_GATE U8486 ( .I1(n14781), .I2(n7562), .O(n7563) );
  NAND_GATE U8487 ( .I1(B[18]), .I2(n7563), .O(n7567) );
  NAND_GATE U8488 ( .I1(n1384), .I2(A[1]), .O(n7564) );
  NAND_GATE U8489 ( .I1(n14784), .I2(n7564), .O(n7565) );
  NAND_GATE U8490 ( .I1(n1382), .I2(n7565), .O(n7566) );
  NAND_GATE U8491 ( .I1(n7567), .I2(n7566), .O(n8151) );
  NAND_GATE U8492 ( .I1(n8149), .I2(n8151), .O(n8146) );
  NAND3_GATE U8493 ( .I1(B[16]), .I2(n1382), .I3(n1196), .O(n8147) );
  INV_GATE U8494 ( .I1(n8147), .O(n8150) );
  INV_GATE U8495 ( .I1(n8151), .O(n8148) );
  NAND_GATE U8496 ( .I1(n8155), .I2(n8148), .O(n7568) );
  NAND_GATE U8497 ( .I1(n8150), .I2(n7568), .O(n7569) );
  NAND_GATE U8498 ( .I1(n8146), .I2(n7569), .O(n8132) );
  NAND_GATE U8499 ( .I1(n7583), .I2(n8132), .O(n8128) );
  OR_GATE U8500 ( .I1(n7571), .I2(n7570), .O(n7582) );
  NAND_GATE U8501 ( .I1(n7572), .I2(n7576), .O(n7580) );
  NAND_GATE U8502 ( .I1(n7574), .I2(n7573), .O(n7575) );
  NAND_GATE U8503 ( .I1(n7576), .I2(n7575), .O(n7577) );
  NAND_GATE U8504 ( .I1(n7578), .I2(n7577), .O(n7579) );
  NAND_GATE U8505 ( .I1(n7580), .I2(n7579), .O(n7581) );
  NAND_GATE U8506 ( .I1(n7582), .I2(n7581), .O(n8131) );
  NAND_GATE U8507 ( .I1(n8132), .I2(n8131), .O(n7584) );
  NAND_GATE U8508 ( .I1(n7583), .I2(n8131), .O(n8127) );
  NAND3_GATE U8509 ( .I1(n8128), .I2(n7584), .I3(n8127), .O(n8169) );
  NAND_GATE U8510 ( .I1(n8167), .I2(n8173), .O(n7585) );
  NAND_GATE U8511 ( .I1(n8169), .I2(n7585), .O(n7586) );
  NAND_GATE U8512 ( .I1(n8164), .I2(n7586), .O(n8121) );
  NAND_GATE U8513 ( .I1(n7601), .I2(n8121), .O(n8116) );
  INV_GATE U8514 ( .I1(n7591), .O(n7588) );
  NAND_GATE U8515 ( .I1(n7589), .I2(n7588), .O(n7594) );
  NAND_GATE U8516 ( .I1(n7590), .I2(n7594), .O(n7598) );
  NAND_GATE U8517 ( .I1(n7592), .I2(n7591), .O(n7593) );
  NAND_GATE U8518 ( .I1(n7594), .I2(n7593), .O(n7595) );
  NAND_GATE U8519 ( .I1(n7596), .I2(n7595), .O(n7597) );
  NAND_GATE U8520 ( .I1(n7598), .I2(n7597), .O(n7599) );
  NAND_GATE U8521 ( .I1(n7600), .I2(n7599), .O(n8120) );
  NAND_GATE U8522 ( .I1(n8121), .I2(n8120), .O(n7602) );
  NAND_GATE U8523 ( .I1(n7601), .I2(n8120), .O(n8115) );
  NAND3_GATE U8524 ( .I1(n8116), .I2(n7602), .I3(n8115), .O(n8186) );
  NAND_GATE U8525 ( .I1(n8184), .I2(n8191), .O(n7603) );
  NAND_GATE U8526 ( .I1(n8186), .I2(n7603), .O(n7604) );
  NAND_GATE U8527 ( .I1(n8182), .I2(n7604), .O(n8108) );
  NAND_GATE U8528 ( .I1(n7614), .I2(n8108), .O(n8110) );
  NAND_GATE U8529 ( .I1(n7608), .I2(n917), .O(n7606) );
  NAND_GATE U8530 ( .I1(n7607), .I2(n7606), .O(n7613) );
  NAND_GATE U8531 ( .I1(n7613), .I2(n7612), .O(n8103) );
  NAND_GATE U8532 ( .I1(n8104), .I2(n8103), .O(n8111) );
  NAND_GATE U8533 ( .I1(n8108), .I2(n8111), .O(n7615) );
  NAND_GATE U8534 ( .I1(n7614), .I2(n8111), .O(n8109) );
  NAND3_GATE U8535 ( .I1(n8110), .I2(n7615), .I3(n8109), .O(n8201) );
  NAND_GATE U8536 ( .I1(n8435), .I2(n8204), .O(n7616) );
  NAND_GATE U8537 ( .I1(n8201), .I2(n7616), .O(n7617) );
  NAND_GATE U8538 ( .I1(n7618), .I2(n7617), .O(n8095) );
  NAND_GATE U8539 ( .I1(n7627), .I2(n8095), .O(n8092) );
  NAND3_GATE U8540 ( .I1(n7620), .I2(n189), .I3(n7619), .O(n7621) );
  NAND3_GATE U8541 ( .I1(n7623), .I2(n7622), .I3(n7621), .O(n7626) );
  NAND_GATE U8542 ( .I1(n1355), .I2(n7624), .O(n7625) );
  NAND_GATE U8543 ( .I1(n7626), .I2(n7625), .O(n8096) );
  NAND_GATE U8544 ( .I1(n8095), .I2(n8096), .O(n7628) );
  NAND_GATE U8545 ( .I1(n7627), .I2(n8096), .O(n8091) );
  NAND3_GATE U8546 ( .I1(n8092), .I2(n7628), .I3(n8091), .O(n8220) );
  NAND_GATE U8547 ( .I1(n8216), .I2(n8213), .O(n7629) );
  NAND_GATE U8548 ( .I1(n8220), .I2(n7629), .O(n7630) );
  NAND_GATE U8549 ( .I1(n8219), .I2(n7630), .O(n8085) );
  NAND_GATE U8550 ( .I1(n7645), .I2(n8085), .O(n8080) );
  INV_GATE U8551 ( .I1(n7641), .O(n7632) );
  NAND_GATE U8552 ( .I1(n7631), .I2(n7635), .O(n7639) );
  NAND_GATE U8553 ( .I1(n7633), .I2(n7632), .O(n7635) );
  NAND_GATE U8554 ( .I1(n1330), .I2(n7641), .O(n7634) );
  NAND_GATE U8555 ( .I1(n7635), .I2(n7634), .O(n7636) );
  NAND_GATE U8556 ( .I1(n7637), .I2(n7636), .O(n7638) );
  NAND_GATE U8557 ( .I1(n7639), .I2(n7638), .O(n7644) );
  INV_GATE U8558 ( .I1(n7640), .O(n7642) );
  NAND_GATE U8559 ( .I1(n7642), .I2(n7641), .O(n7643) );
  NAND_GATE U8560 ( .I1(n7644), .I2(n7643), .O(n8084) );
  NAND_GATE U8561 ( .I1(n8085), .I2(n8084), .O(n7646) );
  NAND_GATE U8562 ( .I1(n7645), .I2(n8084), .O(n8079) );
  NAND3_GATE U8563 ( .I1(n8080), .I2(n7646), .I3(n8079), .O(n8231) );
  NAND_GATE U8564 ( .I1(B[16]), .I2(A[12]), .O(n8230) );
  NAND_GATE U8565 ( .I1(n7650), .I2(n7649), .O(n7653) );
  NAND_GATE U8566 ( .I1(n7654), .I2(n7653), .O(n7651) );
  NAND_GATE U8567 ( .I1(n7652), .I2(n7651), .O(n7656) );
  INV_GATE U8568 ( .I1(n7652), .O(n7661) );
  NAND3_GATE U8569 ( .I1(n7661), .I2(n7654), .I3(n7653), .O(n7655) );
  NAND3_GATE U8570 ( .I1(n7657), .I2(n7656), .I3(n7655), .O(n8234) );
  NAND3_GATE U8571 ( .I1(n8234), .I2(n8233), .I3(n8232), .O(n8241) );
  NAND_GATE U8572 ( .I1(n8230), .I2(n8241), .O(n7662) );
  NAND_GATE U8573 ( .I1(n8231), .I2(n7662), .O(n7664) );
  INV_GATE U8574 ( .I1(n8230), .O(n8245) );
  INV_GATE U8575 ( .I1(n8241), .O(n8229) );
  NAND_GATE U8576 ( .I1(n8245), .I2(n8229), .O(n7663) );
  NAND_GATE U8577 ( .I1(n7664), .I2(n7663), .O(n8073) );
  NAND_GATE U8578 ( .I1(n8074), .I2(n8073), .O(n7666) );
  NAND_GATE U8579 ( .I1(n7665), .I2(n8073), .O(n8075) );
  NAND3_GATE U8580 ( .I1(n8072), .I2(n7666), .I3(n8075), .O(n8066) );
  NAND_GATE U8581 ( .I1(B[16]), .I2(A[14]), .O(n8375) );
  OR_GATE U8582 ( .I1(n7671), .I2(n7667), .O(n7670) );
  OR_GATE U8583 ( .I1(n7668), .I2(n7672), .O(n7669) );
  AND_GATE U8584 ( .I1(n7670), .I2(n7669), .O(n7677) );
  NAND_GATE U8585 ( .I1(n7672), .I2(n937), .O(n7673) );
  NAND3_GATE U8586 ( .I1(n7675), .I2(n7674), .I3(n7673), .O(n7676) );
  NAND_GATE U8587 ( .I1(n7677), .I2(n7676), .O(n8062) );
  NAND_GATE U8588 ( .I1(n8375), .I2(n8062), .O(n7678) );
  NAND_GATE U8589 ( .I1(n8066), .I2(n7678), .O(n7680) );
  INV_GATE U8590 ( .I1(n8375), .O(n8064) );
  NAND_GATE U8591 ( .I1(n8064), .I2(n8065), .O(n7679) );
  NAND_GATE U8592 ( .I1(n7680), .I2(n7679), .O(n8260) );
  NAND_GATE U8593 ( .I1(n7687), .I2(n8260), .O(n8255) );
  NAND_GATE U8594 ( .I1(n1256), .I2(n7685), .O(n7681) );
  NAND_GATE U8595 ( .I1(n1255), .I2(n8258), .O(n8262) );
  NAND_GATE U8596 ( .I1(n7686), .I2(n7681), .O(n8253) );
  NAND_GATE U8597 ( .I1(n8254), .I2(n8253), .O(n8261) );
  NAND3_GATE U8598 ( .I1(n8260), .I2(n8262), .I3(n8261), .O(n7689) );
  NAND_GATE U8599 ( .I1(n8261), .I2(n952), .O(n7688) );
  NAND_GATE U8600 ( .I1(n8291), .I2(n8290), .O(n8294) );
  NAND_GATE U8601 ( .I1(n7691), .I2(n7690), .O(n8282) );
  NAND3_GATE U8602 ( .I1(n8292), .I2(n8294), .I3(n8282), .O(n7692) );
  NAND3_GATE U8603 ( .I1(n8287), .I2(n7692), .I3(n8284), .O(n8057) );
  NAND3_GATE U8604 ( .I1(n7696), .I2(n1344), .I3(n7695), .O(n7697) );
  NAND3_GATE U8605 ( .I1(n7698), .I2(n7485), .I3(n7697), .O(n7699) );
  NAND_GATE U8606 ( .I1(n7700), .I2(n7699), .O(n8055) );
  NAND_GATE U8607 ( .I1(n8057), .I2(n8055), .O(n7702) );
  NAND_GATE U8608 ( .I1(n8051), .I2(n8057), .O(n7701) );
  NAND3_GATE U8609 ( .I1(n8052), .I2(n7702), .I3(n7701), .O(n8306) );
  NAND_GATE U8610 ( .I1(n7710), .I2(n8306), .O(n8038) );
  NAND_GATE U8611 ( .I1(n7703), .I2(n7708), .O(n8040) );
  NAND_GATE U8612 ( .I1(n276), .I2(n7705), .O(n8042) );
  NAND_GATE U8613 ( .I1(n7706), .I2(n7705), .O(n7709) );
  NAND_GATE U8614 ( .I1(n596), .I2(n7707), .O(n7708) );
  NAND_GATE U8615 ( .I1(n7709), .I2(n7708), .O(n8044) );
  NAND_GATE U8616 ( .I1(n8045), .I2(n8044), .O(n8039) );
  NAND3_GATE U8617 ( .I1(n8306), .I2(n8046), .I3(n8039), .O(n7711) );
  NAND3_GATE U8618 ( .I1(n7710), .I2(n8046), .I3(n8039), .O(n8307) );
  NAND3_GATE U8619 ( .I1(n8038), .I2(n7711), .I3(n8307), .O(n8032) );
  NAND_GATE U8620 ( .I1(n8033), .I2(n8032), .O(n7713) );
  NAND_GATE U8621 ( .I1(n7712), .I2(n8032), .O(n8034) );
  NAND3_GATE U8622 ( .I1(n8031), .I2(n7713), .I3(n8034), .O(n8004) );
  NAND_GATE U8623 ( .I1(n8014), .I2(n8004), .O(n8016) );
  NAND_GATE U8624 ( .I1(n7718), .I2(n707), .O(n7714) );
  NAND_GATE U8625 ( .I1(n7715), .I2(n7714), .O(n8011) );
  NAND3_GATE U8626 ( .I1(n7715), .I2(n7716), .I3(n7717), .O(n8013) );
  NAND_GATE U8627 ( .I1(n7717), .I2(n7716), .O(n7719) );
  NAND_GATE U8628 ( .I1(n7719), .I2(n7714), .O(n8008) );
  NAND3_GATE U8629 ( .I1(n8014), .I2(n8002), .I3(n8010), .O(n7721) );
  NAND3_GATE U8630 ( .I1(n8004), .I2(n8002), .I3(n8010), .O(n7720) );
  NAND3_GATE U8631 ( .I1(n8016), .I2(n7721), .I3(n7720), .O(n7997) );
  NAND_GATE U8632 ( .I1(n7728), .I2(n7997), .O(n7986) );
  NAND3_GATE U8633 ( .I1(n7722), .I2(n7723), .I3(n858), .O(n7993) );
  NAND_GATE U8634 ( .I1(n7722), .I2(n7724), .O(n7992) );
  NAND_GATE U8635 ( .I1(n858), .I2(n7723), .O(n7725) );
  NAND_GATE U8636 ( .I1(n7725), .I2(n7724), .O(n7990) );
  NAND_GATE U8637 ( .I1(n7991), .I2(n7990), .O(n7726) );
  NAND_GATE U8638 ( .I1(n7992), .I2(n7726), .O(n7727) );
  NAND_GATE U8639 ( .I1(n7993), .I2(n7727), .O(n7987) );
  NAND_GATE U8640 ( .I1(n7728), .I2(n7987), .O(n7985) );
  NAND_GATE U8641 ( .I1(n7997), .I2(n7987), .O(n7729) );
  NAND3_GATE U8642 ( .I1(n7986), .I2(n7985), .I3(n7729), .O(n7978) );
  NAND_GATE U8643 ( .I1(n7738), .I2(n7978), .O(n7973) );
  NAND_GATE U8644 ( .I1(n1250), .I2(n7730), .O(n7979) );
  INV_GATE U8645 ( .I1(n7730), .O(n7733) );
  NAND_GATE U8646 ( .I1(n7731), .I2(n7730), .O(n7736) );
  NAND3_GATE U8647 ( .I1(n7734), .I2(n7733), .I3(n7732), .O(n7735) );
  NAND3_GATE U8648 ( .I1(n7737), .I2(n7736), .I3(n7735), .O(n7977) );
  NAND_GATE U8649 ( .I1(n7979), .I2(n7977), .O(n7976) );
  NAND_GATE U8650 ( .I1(n7738), .I2(n7976), .O(n7972) );
  NAND_GATE U8651 ( .I1(n7978), .I2(n7976), .O(n7739) );
  NAND3_GATE U8652 ( .I1(n7973), .I2(n7972), .I3(n7739), .O(n7966) );
  NAND_GATE U8653 ( .I1(n7755), .I2(n7966), .O(n7962) );
  INV_GATE U8654 ( .I1(n7740), .O(n7741) );
  NAND_GATE U8655 ( .I1(n7741), .I2(n7744), .O(n7754) );
  INV_GATE U8656 ( .I1(n7744), .O(n7746) );
  NAND_GATE U8657 ( .I1(n7747), .I2(n7746), .O(n7742) );
  NAND_GATE U8658 ( .I1(n7743), .I2(n7742), .O(n7752) );
  NAND_GATE U8659 ( .I1(n7745), .I2(n7744), .O(n7748) );
  NAND_GATE U8660 ( .I1(n7748), .I2(n7742), .O(n7749) );
  NAND_GATE U8661 ( .I1(n7750), .I2(n7749), .O(n7751) );
  NAND_GATE U8662 ( .I1(n7752), .I2(n7751), .O(n7753) );
  NAND_GATE U8663 ( .I1(n7754), .I2(n7753), .O(n7965) );
  NAND_GATE U8664 ( .I1(n7755), .I2(n7965), .O(n7961) );
  NAND_GATE U8665 ( .I1(n7966), .I2(n7965), .O(n7756) );
  NAND3_GATE U8666 ( .I1(n7962), .I2(n7961), .I3(n7756), .O(n7955) );
  NAND_GATE U8667 ( .I1(n7770), .I2(n7955), .O(n7951) );
  INV_GATE U8668 ( .I1(n7757), .O(n7758) );
  NAND_GATE U8669 ( .I1(n7758), .I2(n7761), .O(n7769) );
  NAND_GATE U8670 ( .I1(n7762), .I2(n272), .O(n7759) );
  NAND_GATE U8671 ( .I1(n7760), .I2(n7759), .O(n7767) );
  NAND_GATE U8672 ( .I1(n832), .I2(n7761), .O(n7763) );
  NAND_GATE U8673 ( .I1(n7763), .I2(n7759), .O(n7764) );
  NAND_GATE U8674 ( .I1(n7765), .I2(n7764), .O(n7766) );
  NAND_GATE U8675 ( .I1(n7767), .I2(n7766), .O(n7768) );
  NAND_GATE U8676 ( .I1(n7769), .I2(n7768), .O(n7954) );
  NAND_GATE U8677 ( .I1(n7955), .I2(n7954), .O(n7771) );
  NAND3_GATE U8678 ( .I1(n7951), .I2(n7950), .I3(n7771), .O(n7944) );
  NAND_GATE U8679 ( .I1(n7786), .I2(n7944), .O(n7940) );
  INV_GATE U8680 ( .I1(n7772), .O(n7773) );
  NAND_GATE U8681 ( .I1(n7773), .I2(n7775), .O(n7785) );
  NAND_GATE U8682 ( .I1(n7774), .I2(n7778), .O(n7783) );
  NAND_GATE U8683 ( .I1(n7776), .I2(n7775), .O(n7779) );
  NAND_GATE U8684 ( .I1(n7777), .I2(n90), .O(n7778) );
  NAND_GATE U8685 ( .I1(n7779), .I2(n7778), .O(n7780) );
  NAND_GATE U8686 ( .I1(n7781), .I2(n7780), .O(n7782) );
  NAND_GATE U8687 ( .I1(n7783), .I2(n7782), .O(n7784) );
  NAND_GATE U8688 ( .I1(n7785), .I2(n7784), .O(n7943) );
  NAND_GATE U8689 ( .I1(n7944), .I2(n7943), .O(n7787) );
  NAND3_GATE U8690 ( .I1(n7940), .I2(n7939), .I3(n7787), .O(n7934) );
  NAND_GATE U8691 ( .I1(n7802), .I2(n7934), .O(n7930) );
  INV_GATE U8692 ( .I1(n7788), .O(n7789) );
  NAND_GATE U8693 ( .I1(n7789), .I2(n7792), .O(n7801) );
  NAND_GATE U8694 ( .I1(n7791), .I2(n7795), .O(n7799) );
  NAND_GATE U8695 ( .I1(n7793), .I2(n7792), .O(n7794) );
  NAND_GATE U8696 ( .I1(n7795), .I2(n7794), .O(n7796) );
  NAND_GATE U8697 ( .I1(n7797), .I2(n7796), .O(n7798) );
  NAND_GATE U8698 ( .I1(n7799), .I2(n7798), .O(n7800) );
  NAND_GATE U8699 ( .I1(n7801), .I2(n7800), .O(n7933) );
  NAND_GATE U8700 ( .I1(n7802), .I2(n7933), .O(n7929) );
  NAND_GATE U8701 ( .I1(n7934), .I2(n7933), .O(n7803) );
  NAND3_GATE U8702 ( .I1(n7930), .I2(n7929), .I3(n7803), .O(n7924) );
  NAND_GATE U8703 ( .I1(n7818), .I2(n7924), .O(n7920) );
  INV_GATE U8704 ( .I1(n7804), .O(n7805) );
  NAND_GATE U8705 ( .I1(n7805), .I2(n7808), .O(n7817) );
  NAND_GATE U8706 ( .I1(n7807), .I2(n7811), .O(n7815) );
  NAND_GATE U8707 ( .I1(n7809), .I2(n7808), .O(n7810) );
  NAND_GATE U8708 ( .I1(n7811), .I2(n7810), .O(n7812) );
  NAND_GATE U8709 ( .I1(n7813), .I2(n7812), .O(n7814) );
  NAND_GATE U8710 ( .I1(n7815), .I2(n7814), .O(n7816) );
  NAND_GATE U8711 ( .I1(n7817), .I2(n7816), .O(n7923) );
  NAND_GATE U8712 ( .I1(n7818), .I2(n7923), .O(n7919) );
  NAND_GATE U8713 ( .I1(n7924), .I2(n7923), .O(n7819) );
  NAND3_GATE U8714 ( .I1(n7920), .I2(n7919), .I3(n7819), .O(n7913) );
  NAND_GATE U8715 ( .I1(n7835), .I2(n7913), .O(n7909) );
  INV_GATE U8716 ( .I1(n7820), .O(n7821) );
  NAND_GATE U8717 ( .I1(n7821), .I2(n7825), .O(n7834) );
  INV_GATE U8718 ( .I1(n7825), .O(n7822) );
  NAND_GATE U8719 ( .I1(n7823), .I2(n7822), .O(n7828) );
  NAND_GATE U8720 ( .I1(n7824), .I2(n7828), .O(n7832) );
  NAND_GATE U8721 ( .I1(n7826), .I2(n7825), .O(n7827) );
  NAND_GATE U8722 ( .I1(n7828), .I2(n7827), .O(n7829) );
  NAND_GATE U8723 ( .I1(n7830), .I2(n7829), .O(n7831) );
  NAND_GATE U8724 ( .I1(n7832), .I2(n7831), .O(n7833) );
  NAND_GATE U8725 ( .I1(n7834), .I2(n7833), .O(n7912) );
  NAND_GATE U8726 ( .I1(n7835), .I2(n7912), .O(n7908) );
  NAND_GATE U8727 ( .I1(n7913), .I2(n7912), .O(n7836) );
  NAND3_GATE U8728 ( .I1(n7909), .I2(n7908), .I3(n7836), .O(n7902) );
  NAND_GATE U8729 ( .I1(n7851), .I2(n7902), .O(n7898) );
  INV_GATE U8730 ( .I1(n7837), .O(n7838) );
  NAND_GATE U8731 ( .I1(n7838), .I2(n7841), .O(n7850) );
  NAND_GATE U8732 ( .I1(n7840), .I2(n7844), .O(n7848) );
  NAND_GATE U8733 ( .I1(n7842), .I2(n7841), .O(n7843) );
  NAND_GATE U8734 ( .I1(n7844), .I2(n7843), .O(n7845) );
  NAND_GATE U8735 ( .I1(n7846), .I2(n7845), .O(n7847) );
  NAND_GATE U8736 ( .I1(n7848), .I2(n7847), .O(n7849) );
  NAND_GATE U8737 ( .I1(n7850), .I2(n7849), .O(n7901) );
  NAND_GATE U8738 ( .I1(n7851), .I2(n7901), .O(n7897) );
  NAND_GATE U8739 ( .I1(n7902), .I2(n7901), .O(n7852) );
  NAND3_GATE U8740 ( .I1(n7898), .I2(n7897), .I3(n7852), .O(n7891) );
  NAND_GATE U8741 ( .I1(n7868), .I2(n7891), .O(n7887) );
  INV_GATE U8742 ( .I1(n7853), .O(n7854) );
  NAND_GATE U8743 ( .I1(n7854), .I2(n7858), .O(n7867) );
  INV_GATE U8744 ( .I1(n7858), .O(n7855) );
  NAND_GATE U8745 ( .I1(n7856), .I2(n7855), .O(n7861) );
  NAND_GATE U8746 ( .I1(n7857), .I2(n7861), .O(n7865) );
  NAND_GATE U8747 ( .I1(n7859), .I2(n7858), .O(n7860) );
  NAND_GATE U8748 ( .I1(n7861), .I2(n7860), .O(n7862) );
  NAND_GATE U8749 ( .I1(n7863), .I2(n7862), .O(n7864) );
  NAND_GATE U8750 ( .I1(n7865), .I2(n7864), .O(n7866) );
  NAND_GATE U8751 ( .I1(n7867), .I2(n7866), .O(n7890) );
  NAND_GATE U8752 ( .I1(n7868), .I2(n7890), .O(n7886) );
  NAND_GATE U8753 ( .I1(n7891), .I2(n7890), .O(n7869) );
  NAND3_GATE U8754 ( .I1(n7887), .I2(n7886), .I3(n7869), .O(n15327) );
  INV_GATE U8755 ( .I1(n15327), .O(n7882) );
  INV_GATE U8756 ( .I1(n7870), .O(n7871) );
  NAND_GATE U8757 ( .I1(n7871), .I2(n7873), .O(n7881) );
  NAND_GATE U8758 ( .I1(n7872), .I2(n7875), .O(n7879) );
  NAND_GATE U8759 ( .I1(n472), .I2(n7873), .O(n7874) );
  NAND_GATE U8760 ( .I1(n7875), .I2(n7874), .O(n7876) );
  NAND_GATE U8761 ( .I1(n7877), .I2(n7876), .O(n7878) );
  NAND_GATE U8762 ( .I1(n7879), .I2(n7878), .O(n7880) );
  NAND_GATE U8763 ( .I1(n7881), .I2(n7880), .O(n15326) );
  NAND_GATE U8764 ( .I1(n7882), .I2(n15326), .O(n7885) );
  INV_GATE U8765 ( .I1(n15326), .O(n7883) );
  NAND_GATE U8766 ( .I1(n15327), .I2(n7883), .O(n7884) );
  NAND_GATE U8767 ( .I1(n7885), .I2(n7884), .O(\A1[46] ) );
  OR_GATE U8768 ( .I1(n7886), .I2(n7891), .O(n7889) );
  OR_GATE U8769 ( .I1(n7890), .I2(n7887), .O(n7888) );
  AND_GATE U8770 ( .I1(n7889), .I2(n7888), .O(n7896) );
  NAND_GATE U8771 ( .I1(n914), .I2(n7890), .O(n7894) );
  NAND3_GATE U8772 ( .I1(n7894), .I2(n7893), .I3(n7892), .O(n7895) );
  NAND_GATE U8773 ( .I1(n7896), .I2(n7895), .O(n8337) );
  OR_GATE U8774 ( .I1(n7897), .I2(n7902), .O(n7900) );
  OR_GATE U8775 ( .I1(n7901), .I2(n7898), .O(n7899) );
  AND_GATE U8776 ( .I1(n7900), .I2(n7899), .O(n7907) );
  NAND_GATE U8777 ( .I1(n913), .I2(n7901), .O(n7905) );
  NAND3_GATE U8778 ( .I1(n7905), .I2(n7904), .I3(n7903), .O(n7906) );
  NAND_GATE U8779 ( .I1(n7907), .I2(n7906), .O(n8767) );
  INV_GATE U8780 ( .I1(n8767), .O(n8770) );
  NAND_GATE U8781 ( .I1(n1379), .I2(A[31]), .O(n8774) );
  INV_GATE U8782 ( .I1(n8774), .O(n8768) );
  NAND_GATE U8783 ( .I1(n8770), .I2(n8768), .O(n8765) );
  OR_GATE U8784 ( .I1(n7908), .I2(n7913), .O(n7911) );
  OR_GATE U8785 ( .I1(n7912), .I2(n7909), .O(n7910) );
  AND_GATE U8786 ( .I1(n7911), .I2(n7910), .O(n7918) );
  NAND_GATE U8787 ( .I1(n911), .I2(n7912), .O(n7916) );
  NAND3_GATE U8788 ( .I1(n7916), .I2(n7915), .I3(n7914), .O(n7917) );
  NAND_GATE U8789 ( .I1(n7918), .I2(n7917), .O(n8751) );
  INV_GATE U8790 ( .I1(n8751), .O(n8754) );
  NAND_GATE U8791 ( .I1(n1379), .I2(A[30]), .O(n8758) );
  INV_GATE U8792 ( .I1(n8758), .O(n8752) );
  NAND_GATE U8793 ( .I1(n8754), .I2(n8752), .O(n8748) );
  OR_GATE U8794 ( .I1(n7919), .I2(n7924), .O(n7922) );
  OR_GATE U8795 ( .I1(n7923), .I2(n7920), .O(n7921) );
  NAND_GATE U8796 ( .I1(n905), .I2(n7923), .O(n7927) );
  NAND3_GATE U8797 ( .I1(n7927), .I2(n7926), .I3(n7925), .O(n7928) );
  NAND_GATE U8798 ( .I1(n1379), .I2(A[29]), .O(n8741) );
  INV_GATE U8799 ( .I1(n8741), .O(n8735) );
  NAND_GATE U8800 ( .I1(n8737), .I2(n8735), .O(n8732) );
  OR_GATE U8801 ( .I1(n7929), .I2(n7934), .O(n7932) );
  OR_GATE U8802 ( .I1(n7933), .I2(n7930), .O(n7931) );
  NAND_GATE U8803 ( .I1(n904), .I2(n7933), .O(n7937) );
  NAND3_GATE U8804 ( .I1(n7937), .I2(n7936), .I3(n7935), .O(n7938) );
  NAND_GATE U8805 ( .I1(n1379), .I2(A[28]), .O(n8725) );
  INV_GATE U8806 ( .I1(n8725), .O(n8719) );
  NAND_GATE U8807 ( .I1(n8721), .I2(n8719), .O(n8716) );
  OR_GATE U8808 ( .I1(n7943), .I2(n7940), .O(n7941) );
  AND_GATE U8809 ( .I1(n7942), .I2(n7941), .O(n7949) );
  NAND_GATE U8810 ( .I1(n887), .I2(n7943), .O(n7947) );
  NAND3_GATE U8811 ( .I1(n7947), .I2(n7946), .I3(n7945), .O(n7948) );
  NAND_GATE U8812 ( .I1(n7949), .I2(n7948), .O(n8707) );
  NAND_GATE U8813 ( .I1(n1379), .I2(A[27]), .O(n8709) );
  INV_GATE U8814 ( .I1(n8709), .O(n8703) );
  NAND_GATE U8815 ( .I1(n8705), .I2(n8703), .O(n8700) );
  OR_GATE U8816 ( .I1(n7950), .I2(n7955), .O(n7953) );
  OR_GATE U8817 ( .I1(n7954), .I2(n7951), .O(n7952) );
  AND_GATE U8818 ( .I1(n7953), .I2(n7952), .O(n7960) );
  NAND_GATE U8819 ( .I1(n886), .I2(n7954), .O(n7958) );
  NAND3_GATE U8820 ( .I1(n7958), .I2(n7957), .I3(n7956), .O(n7959) );
  NAND_GATE U8821 ( .I1(n7960), .I2(n7959), .O(n8689) );
  NAND_GATE U8822 ( .I1(n1379), .I2(A[26]), .O(n8693) );
  INV_GATE U8823 ( .I1(n8693), .O(n8686) );
  NAND_GATE U8824 ( .I1(n831), .I2(n8686), .O(n8684) );
  OR_GATE U8825 ( .I1(n7965), .I2(n7962), .O(n7963) );
  AND_GATE U8826 ( .I1(n7964), .I2(n7963), .O(n7971) );
  NAND_GATE U8827 ( .I1(n885), .I2(n7965), .O(n7969) );
  NAND3_GATE U8828 ( .I1(n7969), .I2(n7968), .I3(n7967), .O(n7970) );
  NAND_GATE U8829 ( .I1(n7971), .I2(n7970), .O(n8674) );
  NAND_GATE U8830 ( .I1(n1379), .I2(A[25]), .O(n8677) );
  INV_GATE U8831 ( .I1(n8677), .O(n8670) );
  NAND_GATE U8832 ( .I1(n8672), .I2(n8670), .O(n8667) );
  OR_GATE U8833 ( .I1(n7976), .I2(n7973), .O(n7974) );
  AND_GATE U8834 ( .I1(n7975), .I2(n7974), .O(n7984) );
  NAND_GATE U8835 ( .I1(n18), .I2(n7976), .O(n7982) );
  NAND3_GATE U8836 ( .I1(n7979), .I2(n7978), .I3(n7977), .O(n7981) );
  NAND3_GATE U8837 ( .I1(n7982), .I2(n7981), .I3(n7980), .O(n7983) );
  NAND_GATE U8838 ( .I1(n7984), .I2(n7983), .O(n8659) );
  INV_GATE U8839 ( .I1(n8659), .O(n8658) );
  NAND_GATE U8840 ( .I1(n1379), .I2(A[24]), .O(n8662) );
  INV_GATE U8841 ( .I1(n8662), .O(n8657) );
  NAND_GATE U8842 ( .I1(n8658), .I2(n8657), .O(n8655) );
  NAND_GATE U8843 ( .I1(n1379), .I2(A[23]), .O(n8643) );
  INV_GATE U8844 ( .I1(n8643), .O(n8647) );
  OR_GATE U8845 ( .I1(n7985), .I2(n7997), .O(n7989) );
  OR_GATE U8846 ( .I1(n7987), .I2(n7986), .O(n7988) );
  INV_GATE U8847 ( .I1(n7997), .O(n7994) );
  NAND3_GATE U8848 ( .I1(n7726), .I2(n7994), .I3(n7995), .O(n8000) );
  NAND_GATE U8849 ( .I1(n7995), .I2(n7726), .O(n7996) );
  NAND_GATE U8850 ( .I1(n7997), .I2(n7996), .O(n7999) );
  NAND3_GATE U8851 ( .I1(n8000), .I2(n7999), .I3(n7998), .O(n8001) );
  INV_GATE U8852 ( .I1(n8642), .O(n8645) );
  NAND_GATE U8853 ( .I1(n8647), .I2(n8645), .O(n8321) );
  NAND_GATE U8854 ( .I1(n1379), .I2(A[22]), .O(n8882) );
  INV_GATE U8855 ( .I1(n8882), .O(n8633) );
  NAND3_GATE U8856 ( .I1(n8002), .I2(n8010), .I3(n8015), .O(n8007) );
  NAND_GATE U8857 ( .I1(n8002), .I2(n8010), .O(n8003) );
  NAND_GATE U8858 ( .I1(n8004), .I2(n8003), .O(n8006) );
  NAND3_GATE U8859 ( .I1(n8007), .I2(n8006), .I3(n8005), .O(n8020) );
  NAND_GATE U8860 ( .I1(n8009), .I2(n8008), .O(n8010) );
  NAND_GATE U8861 ( .I1(n8011), .I2(n8010), .O(n8012) );
  NAND_GATE U8862 ( .I1(n8013), .I2(n8012), .O(n8017) );
  NAND3_GATE U8863 ( .I1(n8015), .I2(n8017), .I3(n8014), .O(n8019) );
  OR_GATE U8864 ( .I1(n8017), .I2(n8016), .O(n8018) );
  NAND3_GATE U8865 ( .I1(n8020), .I2(n8019), .I3(n8018), .O(n8637) );
  NAND_GATE U8866 ( .I1(n8633), .I2(n8635), .O(n8318) );
  NAND_GATE U8867 ( .I1(n1379), .I2(A[21]), .O(n8892) );
  INV_GATE U8868 ( .I1(n8892), .O(n8340) );
  NAND_GATE U8869 ( .I1(n7479), .I2(n8027), .O(n8025) );
  NAND_GATE U8870 ( .I1(n8032), .I2(n8025), .O(n8029) );
  INV_GATE U8871 ( .I1(n8032), .O(n8026) );
  NAND3_GATE U8872 ( .I1(n8027), .I2(n8026), .I3(n7479), .O(n8028) );
  NAND3_GATE U8873 ( .I1(n8030), .I2(n8029), .I3(n8028), .O(n8037) );
  OR_GATE U8874 ( .I1(n8032), .I2(n8031), .O(n8036) );
  OR_GATE U8875 ( .I1(n8034), .I2(n8033), .O(n8035) );
  NAND3_GATE U8876 ( .I1(n8037), .I2(n8036), .I3(n8035), .O(n8344) );
  INV_GATE U8877 ( .I1(n8344), .O(n8342) );
  NAND_GATE U8878 ( .I1(n8340), .I2(n8342), .O(n8315) );
  INV_GATE U8879 ( .I1(n8038), .O(n8043) );
  NAND_GATE U8880 ( .I1(n8040), .I2(n8039), .O(n8041) );
  NAND3_GATE U8881 ( .I1(n8043), .I2(n8042), .I3(n8041), .O(n8310) );
  NAND_GATE U8882 ( .I1(n8046), .I2(n8039), .O(n8047) );
  NAND_GATE U8883 ( .I1(n8306), .I2(n8047), .O(n8050) );
  OR_GATE U8884 ( .I1(n8047), .I2(n8306), .O(n8049) );
  NAND3_GATE U8885 ( .I1(n8050), .I2(n8049), .I3(n8048), .O(n8308) );
  NAND_GATE U8886 ( .I1(n1379), .I2(A[19]), .O(n8919) );
  INV_GATE U8887 ( .I1(n8919), .O(n8607) );
  NAND3_GATE U8888 ( .I1(n551), .I2(n8051), .I3(n8057), .O(n8054) );
  OR_GATE U8889 ( .I1(n8057), .I2(n8052), .O(n8053) );
  INV_GATE U8890 ( .I1(n8057), .O(n8056) );
  NAND_GATE U8891 ( .I1(n8056), .I2(n8055), .O(n8059) );
  NAND_GATE U8892 ( .I1(n8057), .I2(n551), .O(n8058) );
  NAND3_GATE U8893 ( .I1(n8060), .I2(n8059), .I3(n8058), .O(n8061) );
  INV_GATE U8894 ( .I1(n8608), .O(n8609) );
  NAND_GATE U8895 ( .I1(n8607), .I2(n8609), .O(n8305) );
  NAND_GATE U8896 ( .I1(n1379), .I2(A[17]), .O(n8354) );
  INV_GATE U8897 ( .I1(n8354), .O(n8347) );
  NAND_GATE U8898 ( .I1(n1379), .I2(A[16]), .O(n8359) );
  INV_GATE U8899 ( .I1(n8359), .O(n8363) );
  NAND_GATE U8900 ( .I1(n1379), .I2(A[15]), .O(n8387) );
  INV_GATE U8901 ( .I1(n8387), .O(n8251) );
  INV_GATE U8902 ( .I1(n8066), .O(n8063) );
  NAND_GATE U8903 ( .I1(n8063), .I2(n8062), .O(n8068) );
  NAND_GATE U8904 ( .I1(n8064), .I2(n8068), .O(n8376) );
  NAND3_GATE U8905 ( .I1(n8066), .I2(n8064), .I3(n8065), .O(n8378) );
  NAND_GATE U8906 ( .I1(n8066), .I2(n8065), .O(n8067) );
  NAND_GATE U8907 ( .I1(n8068), .I2(n8067), .O(n8374) );
  NAND_GATE U8908 ( .I1(n8375), .I2(n8374), .O(n8385) );
  NAND3_GATE U8909 ( .I1(n8251), .I2(n8384), .I3(n8385), .O(n8381) );
  NAND_GATE U8910 ( .I1(n8074), .I2(n1258), .O(n8069) );
  NAND3_GATE U8911 ( .I1(n8071), .I2(n8070), .I3(n8069), .O(n8078) );
  OR_GATE U8912 ( .I1(n8073), .I2(n8072), .O(n8077) );
  OR_GATE U8913 ( .I1(n8075), .I2(n8074), .O(n8076) );
  NAND3_GATE U8914 ( .I1(n8078), .I2(n8077), .I3(n8076), .O(n8397) );
  NAND_GATE U8915 ( .I1(n1379), .I2(A[14]), .O(n8584) );
  INV_GATE U8916 ( .I1(n8584), .O(n8394) );
  NAND_GATE U8917 ( .I1(n673), .I2(n8394), .O(n8395) );
  NAND_GATE U8918 ( .I1(n1379), .I2(A[13]), .O(n8399) );
  INV_GATE U8919 ( .I1(n8399), .O(n8238) );
  NAND_GATE U8920 ( .I1(n1379), .I2(A[12]), .O(n8415) );
  INV_GATE U8921 ( .I1(n8415), .O(n8409) );
  OR_GATE U8922 ( .I1(n8079), .I2(n8085), .O(n8082) );
  OR_GATE U8923 ( .I1(n8084), .I2(n8080), .O(n8081) );
  AND_GATE U8924 ( .I1(n8082), .I2(n8081), .O(n8090) );
  INV_GATE U8925 ( .I1(n8085), .O(n8083) );
  NAND_GATE U8926 ( .I1(n8083), .I2(n8084), .O(n8087) );
  NAND_GATE U8927 ( .I1(n8085), .I2(n526), .O(n8086) );
  NAND3_GATE U8928 ( .I1(n8088), .I2(n8087), .I3(n8086), .O(n8089) );
  NAND_GATE U8929 ( .I1(n8409), .I2(n1329), .O(n8418) );
  NAND_GATE U8930 ( .I1(n1379), .I2(A[11]), .O(n8431) );
  INV_GATE U8931 ( .I1(n8431), .O(n8224) );
  NAND_GATE U8932 ( .I1(n1379), .I2(A[10]), .O(n8567) );
  INV_GATE U8933 ( .I1(n8567), .O(n8563) );
  OR_GATE U8934 ( .I1(n8096), .I2(n8092), .O(n8093) );
  AND_GATE U8935 ( .I1(n8094), .I2(n8093), .O(n8101) );
  NAND_GATE U8936 ( .I1(n173), .I2(n8096), .O(n8097) );
  NAND3_GATE U8937 ( .I1(n8099), .I2(n8098), .I3(n8097), .O(n8100) );
  NAND_GATE U8938 ( .I1(n8101), .I2(n8100), .O(n8566) );
  INV_GATE U8939 ( .I1(n8566), .O(n8564) );
  NAND_GATE U8940 ( .I1(n8563), .I2(n8564), .O(n8570) );
  NAND_GATE U8941 ( .I1(n1379), .I2(A[9]), .O(n8447) );
  INV_GATE U8942 ( .I1(n8447), .O(n8207) );
  INV_GATE U8943 ( .I1(n8108), .O(n8102) );
  NAND_GATE U8944 ( .I1(n8102), .I2(n8111), .O(n8107) );
  NAND3_GATE U8945 ( .I1(n8104), .I2(n8108), .I3(n8103), .O(n8106) );
  NAND3_GATE U8946 ( .I1(n8107), .I2(n8106), .I3(n8105), .O(n8114) );
  OR_GATE U8947 ( .I1(n8109), .I2(n8108), .O(n8113) );
  OR_GATE U8948 ( .I1(n8111), .I2(n8110), .O(n8112) );
  NAND_GATE U8949 ( .I1(n1379), .I2(A[8]), .O(n8553) );
  NAND_GATE U8950 ( .I1(n874), .I2(n731), .O(n8548) );
  NAND_GATE U8951 ( .I1(n1379), .I2(A[7]), .O(n8459) );
  INV_GATE U8952 ( .I1(n8459), .O(n8196) );
  OR_GATE U8953 ( .I1(n8120), .I2(n8116), .O(n8117) );
  AND_GATE U8954 ( .I1(n8118), .I2(n8117), .O(n8126) );
  INV_GATE U8955 ( .I1(n8121), .O(n8119) );
  NAND_GATE U8956 ( .I1(n8119), .I2(n8120), .O(n8124) );
  NAND_GATE U8957 ( .I1(n8121), .I2(n1287), .O(n8123) );
  NAND3_GATE U8958 ( .I1(n8124), .I2(n8123), .I3(n8122), .O(n8125) );
  NAND_GATE U8959 ( .I1(n8126), .I2(n8125), .O(n8533) );
  INV_GATE U8960 ( .I1(n8533), .O(n8536) );
  NAND_GATE U8961 ( .I1(n1379), .I2(A[6]), .O(n8540) );
  INV_GATE U8962 ( .I1(n8540), .O(n8534) );
  NAND_GATE U8963 ( .I1(n8536), .I2(n8534), .O(n8530) );
  NAND_GATE U8964 ( .I1(n1379), .I2(A[5]), .O(n8469) );
  INV_GATE U8965 ( .I1(n8469), .O(n8178) );
  OR_GATE U8966 ( .I1(n8131), .I2(n8128), .O(n8129) );
  AND_GATE U8967 ( .I1(n8130), .I2(n8129), .O(n8137) );
  NAND_GATE U8968 ( .I1(n1160), .I2(n8131), .O(n8135) );
  NAND3_GATE U8969 ( .I1(n8135), .I2(n8134), .I3(n8133), .O(n8136) );
  NAND_GATE U8970 ( .I1(n8137), .I2(n8136), .O(n8514) );
  INV_GATE U8971 ( .I1(n8514), .O(n8517) );
  NAND_GATE U8972 ( .I1(n1379), .I2(A[4]), .O(n8521) );
  INV_GATE U8973 ( .I1(n8521), .O(n8515) );
  NAND_GATE U8974 ( .I1(n8517), .I2(n8515), .O(n8511) );
  NAND_GATE U8975 ( .I1(n1379), .I2(A[3]), .O(n8480) );
  INV_GATE U8976 ( .I1(n8480), .O(n8160) );
  NAND_GATE U8977 ( .I1(n1379), .I2(A[2]), .O(n8502) );
  INV_GATE U8978 ( .I1(n8502), .O(n8496) );
  NAND_GATE U8979 ( .I1(n1381), .I2(A[0]), .O(n8138) );
  NAND_GATE U8980 ( .I1(n14781), .I2(n8138), .O(n8139) );
  NAND_GATE U8981 ( .I1(n1382), .I2(n8139), .O(n8143) );
  NAND_GATE U8982 ( .I1(n1383), .I2(A[1]), .O(n8140) );
  NAND_GATE U8983 ( .I1(n14784), .I2(n8140), .O(n8141) );
  NAND_GATE U8984 ( .I1(B[16]), .I2(n8141), .O(n8142) );
  NAND_GATE U8985 ( .I1(n8143), .I2(n8142), .O(n8498) );
  NAND_GATE U8986 ( .I1(n8496), .I2(n8498), .O(n8493) );
  NAND3_GATE U8987 ( .I1(n1379), .I2(B[16]), .I3(n1196), .O(n8494) );
  INV_GATE U8988 ( .I1(n8494), .O(n8497) );
  INV_GATE U8989 ( .I1(n8498), .O(n8495) );
  NAND_GATE U8990 ( .I1(n8502), .I2(n8495), .O(n8144) );
  NAND_GATE U8991 ( .I1(n8497), .I2(n8144), .O(n8145) );
  NAND_GATE U8992 ( .I1(n8493), .I2(n8145), .O(n8479) );
  NAND_GATE U8993 ( .I1(n8160), .I2(n8479), .O(n8475) );
  OR_GATE U8994 ( .I1(n8147), .I2(n8146), .O(n8159) );
  NAND_GATE U8995 ( .I1(n8148), .I2(n8147), .O(n8153) );
  NAND_GATE U8996 ( .I1(n8149), .I2(n8153), .O(n8157) );
  NAND_GATE U8997 ( .I1(n8151), .I2(n8150), .O(n8152) );
  NAND_GATE U8998 ( .I1(n8153), .I2(n8152), .O(n8154) );
  NAND_GATE U8999 ( .I1(n8155), .I2(n8154), .O(n8156) );
  NAND_GATE U9000 ( .I1(n8157), .I2(n8156), .O(n8158) );
  NAND_GATE U9001 ( .I1(n8159), .I2(n8158), .O(n8478) );
  NAND_GATE U9002 ( .I1(n8479), .I2(n8478), .O(n8161) );
  NAND_GATE U9003 ( .I1(n8160), .I2(n8478), .O(n8474) );
  NAND3_GATE U9004 ( .I1(n8475), .I2(n8161), .I3(n8474), .O(n8516) );
  NAND_GATE U9005 ( .I1(n8514), .I2(n8521), .O(n8162) );
  NAND_GATE U9006 ( .I1(n8516), .I2(n8162), .O(n8163) );
  NAND_GATE U9007 ( .I1(n8511), .I2(n8163), .O(n8468) );
  NAND_GATE U9008 ( .I1(n8178), .I2(n8468), .O(n8464) );
  INV_GATE U9009 ( .I1(n8164), .O(n8165) );
  NAND_GATE U9010 ( .I1(n8165), .I2(n8169), .O(n8177) );
  INV_GATE U9011 ( .I1(n8169), .O(n8166) );
  NAND_GATE U9012 ( .I1(n8167), .I2(n8166), .O(n8171) );
  NAND_GATE U9013 ( .I1(n8168), .I2(n8171), .O(n8175) );
  NAND_GATE U9014 ( .I1(n607), .I2(n8169), .O(n8170) );
  NAND_GATE U9015 ( .I1(n8171), .I2(n8170), .O(n8172) );
  NAND_GATE U9016 ( .I1(n8173), .I2(n8172), .O(n8174) );
  NAND_GATE U9017 ( .I1(n8175), .I2(n8174), .O(n8176) );
  NAND_GATE U9018 ( .I1(n8177), .I2(n8176), .O(n8467) );
  NAND_GATE U9019 ( .I1(n8468), .I2(n8467), .O(n8179) );
  NAND_GATE U9020 ( .I1(n8178), .I2(n8467), .O(n8463) );
  NAND3_GATE U9021 ( .I1(n8464), .I2(n8179), .I3(n8463), .O(n8535) );
  NAND_GATE U9022 ( .I1(n8533), .I2(n8540), .O(n8180) );
  NAND_GATE U9023 ( .I1(n8535), .I2(n8180), .O(n8181) );
  NAND_GATE U9024 ( .I1(n8530), .I2(n8181), .O(n8458) );
  NAND_GATE U9025 ( .I1(n8196), .I2(n8458), .O(n8454) );
  INV_GATE U9026 ( .I1(n8182), .O(n8183) );
  NAND_GATE U9027 ( .I1(n8183), .I2(n8186), .O(n8195) );
  NAND_GATE U9028 ( .I1(n8184), .I2(n859), .O(n8189) );
  NAND_GATE U9029 ( .I1(n8185), .I2(n8189), .O(n8193) );
  NAND_GATE U9030 ( .I1(n8189), .I2(n8188), .O(n8190) );
  NAND_GATE U9031 ( .I1(n8191), .I2(n8190), .O(n8192) );
  NAND_GATE U9032 ( .I1(n8193), .I2(n8192), .O(n8194) );
  NAND_GATE U9033 ( .I1(n8195), .I2(n8194), .O(n8457) );
  NAND_GATE U9034 ( .I1(n8458), .I2(n8457), .O(n8197) );
  NAND_GATE U9035 ( .I1(n8196), .I2(n8457), .O(n8453) );
  NAND3_GATE U9036 ( .I1(n8454), .I2(n8197), .I3(n8453), .O(n8550) );
  NAND_GATE U9037 ( .I1(n158), .I2(n8553), .O(n8198) );
  NAND_GATE U9038 ( .I1(n8550), .I2(n8198), .O(n8199) );
  NAND_GATE U9039 ( .I1(n8548), .I2(n8199), .O(n8446) );
  NAND_GATE U9040 ( .I1(n8207), .I2(n8446), .O(n8438) );
  INV_GATE U9041 ( .I1(n8201), .O(n8203) );
  NAND3_GATE U9042 ( .I1(n8201), .I2(n8202), .I3(n8200), .O(n8441) );
  NAND_GATE U9043 ( .I1(n1261), .I2(n8441), .O(n8444) );
  NAND_GATE U9044 ( .I1(n8202), .I2(n8201), .O(n8206) );
  NAND_GATE U9045 ( .I1(n8204), .I2(n8203), .O(n8205) );
  NAND_GATE U9046 ( .I1(n8206), .I2(n8205), .O(n8434) );
  NAND3_GATE U9047 ( .I1(n8446), .I2(n8444), .I3(n8436), .O(n8208) );
  NAND3_GATE U9048 ( .I1(n8207), .I2(n8444), .I3(n8436), .O(n8442) );
  NAND3_GATE U9049 ( .I1(n8438), .I2(n8208), .I3(n8442), .O(n8571) );
  NAND_GATE U9050 ( .I1(n8567), .I2(n8566), .O(n8209) );
  NAND_GATE U9051 ( .I1(n8571), .I2(n8209), .O(n8210) );
  NAND_GATE U9052 ( .I1(n8570), .I2(n8210), .O(n8428) );
  NAND_GATE U9053 ( .I1(n8224), .I2(n8428), .O(n8423) );
  NAND_GATE U9054 ( .I1(n8213), .I2(n165), .O(n8211) );
  NAND_GATE U9055 ( .I1(n8212), .I2(n8211), .O(n8218) );
  NAND_GATE U9056 ( .I1(n1205), .I2(n8220), .O(n8214) );
  NAND_GATE U9057 ( .I1(n8214), .I2(n8211), .O(n8215) );
  NAND_GATE U9058 ( .I1(n8216), .I2(n8215), .O(n8217) );
  NAND_GATE U9059 ( .I1(n8218), .I2(n8217), .O(n8223) );
  INV_GATE U9060 ( .I1(n8219), .O(n8221) );
  NAND_GATE U9061 ( .I1(n8221), .I2(n8220), .O(n8222) );
  NAND_GATE U9062 ( .I1(n8223), .I2(n8222), .O(n8427) );
  NAND_GATE U9063 ( .I1(n8428), .I2(n8427), .O(n8225) );
  NAND_GATE U9064 ( .I1(n8224), .I2(n8427), .O(n8422) );
  NAND3_GATE U9065 ( .I1(n8423), .I2(n8225), .I3(n8422), .O(n8419) );
  NAND_GATE U9066 ( .I1(n8415), .I2(n8411), .O(n8226) );
  NAND_GATE U9067 ( .I1(n8419), .I2(n8226), .O(n8227) );
  NAND_GATE U9068 ( .I1(n8231), .I2(n8245), .O(n8236) );
  INV_GATE U9069 ( .I1(n8236), .O(n8228) );
  NAND_GATE U9070 ( .I1(n8229), .I2(n8228), .O(n8243) );
  INV_GATE U9071 ( .I1(n8231), .O(n8242) );
  NAND3_GATE U9072 ( .I1(n8242), .I2(n8230), .I3(n8241), .O(n8240) );
  NAND3_GATE U9073 ( .I1(n8231), .I2(n8230), .I3(n8229), .O(n8239) );
  NAND4_GATE U9074 ( .I1(n8234), .I2(n8233), .I3(n8245), .I4(n8232), .O(n8235)
         );
  NAND4_GATE U9075 ( .I1(n8236), .I2(n8240), .I3(n8239), .I4(n8235), .O(n8237)
         );
  NAND_GATE U9076 ( .I1(n8243), .I2(n8237), .O(n8405) );
  NAND_GATE U9077 ( .I1(n8402), .I2(n8405), .O(n8248) );
  AND3_GATE U9078 ( .I1(n8240), .I2(n8239), .I3(n8238), .O(n8247) );
  NAND_GATE U9079 ( .I1(n8242), .I2(n8241), .O(n8244) );
  NAND3_GATE U9080 ( .I1(n8245), .I2(n8244), .I3(n8243), .O(n8246) );
  NAND_GATE U9081 ( .I1(n8247), .I2(n8246), .O(n8403) );
  NAND_GATE U9082 ( .I1(n8397), .I2(n8584), .O(n8249) );
  NAND_GATE U9083 ( .I1(n8396), .I2(n8249), .O(n8250) );
  NAND_GATE U9084 ( .I1(n8395), .I2(n8250), .O(n8383) );
  NAND3_GATE U9085 ( .I1(n8384), .I2(n8383), .I3(n8385), .O(n8252) );
  NAND_GATE U9086 ( .I1(n8251), .I2(n8383), .O(n8377) );
  NAND3_GATE U9087 ( .I1(n8381), .I2(n8252), .I3(n8377), .O(n8358) );
  NAND_GATE U9088 ( .I1(n8363), .I2(n8358), .O(n8364) );
  INV_GATE U9089 ( .I1(n8255), .O(n8256) );
  NAND3_GATE U9090 ( .I1(n8258), .I2(n8257), .I3(n8256), .O(n8268) );
  NAND3_GATE U9091 ( .I1(n245), .I2(n952), .I3(n8261), .O(n8267) );
  NAND_GATE U9092 ( .I1(n8262), .I2(n8261), .O(n8259) );
  NAND_GATE U9093 ( .I1(n8260), .I2(n8259), .O(n8264) );
  NAND3_GATE U9094 ( .I1(n245), .I2(n8262), .I3(n8261), .O(n8263) );
  NAND3_GATE U9095 ( .I1(n8265), .I2(n8264), .I3(n8263), .O(n8266) );
  NAND3_GATE U9096 ( .I1(n8268), .I2(n8267), .I3(n8266), .O(n8360) );
  INV_GATE U9097 ( .I1(n8358), .O(n8361) );
  NAND_GATE U9098 ( .I1(n8359), .I2(n8361), .O(n8269) );
  NAND_GATE U9099 ( .I1(n8365), .I2(n8269), .O(n8270) );
  NAND_GATE U9100 ( .I1(n8364), .I2(n8270), .O(n8351) );
  NAND_GATE U9101 ( .I1(n8347), .I2(n8351), .O(n8348) );
  NAND3_GATE U9102 ( .I1(n8272), .I2(n1360), .I3(n8271), .O(n8275) );
  NAND_GATE U9103 ( .I1(n8272), .I2(n1360), .O(n8273) );
  NAND3_GATE U9104 ( .I1(n8274), .I2(n8273), .I3(n8279), .O(n8346) );
  NAND3_GATE U9105 ( .I1(n990), .I2(n8346), .I3(n8347), .O(n8281) );
  NAND_GATE U9106 ( .I1(n8274), .I2(n8273), .O(n8276) );
  NAND3_GATE U9107 ( .I1(n8277), .I2(n8276), .I3(n8275), .O(n8278) );
  NAND_GATE U9108 ( .I1(n8279), .I2(n8278), .O(n8350) );
  NAND_GATE U9109 ( .I1(n8351), .I2(n8350), .O(n8280) );
  NAND_GATE U9110 ( .I1(n1379), .I2(A[18]), .O(n9179) );
  NAND_GATE U9111 ( .I1(n8283), .I2(n8282), .O(n8286) );
  NAND3_GATE U9112 ( .I1(n8286), .I2(n202), .I3(n8285), .O(n8289) );
  OR_GATE U9113 ( .I1(n8294), .I2(n8287), .O(n8288) );
  AND_GATE U9114 ( .I1(n8289), .I2(n8288), .O(n8299) );
  NAND4_GATE U9115 ( .I1(n8291), .I2(n8290), .I3(n8282), .I4(n8292), .O(n8297)
         );
  NAND_GATE U9116 ( .I1(n8282), .I2(n8292), .O(n8293) );
  NAND_GATE U9117 ( .I1(n8294), .I2(n8293), .O(n8296) );
  NAND3_GATE U9118 ( .I1(n8297), .I2(n8296), .I3(n8295), .O(n8298) );
  NAND_GATE U9119 ( .I1(n8299), .I2(n8298), .O(n8601) );
  NAND_GATE U9120 ( .I1(n9179), .I2(n8601), .O(n8300) );
  NAND_GATE U9121 ( .I1(n8603), .I2(n8300), .O(n8302) );
  INV_GATE U9122 ( .I1(n9179), .O(n8602) );
  NAND_GATE U9123 ( .I1(n8602), .I2(n807), .O(n8301) );
  NAND_GATE U9124 ( .I1(n8919), .I2(n8608), .O(n8303) );
  NAND_GATE U9125 ( .I1(n252), .I2(n8303), .O(n8304) );
  NAND_GATE U9126 ( .I1(n8305), .I2(n8304), .O(n8617) );
  NAND4_GATE U9127 ( .I1(n8310), .I2(n8308), .I3(n8617), .I4(n8309), .O(n8312)
         );
  NAND_GATE U9128 ( .I1(n1379), .I2(A[20]), .O(n8914) );
  INV_GATE U9129 ( .I1(n8914), .O(n8615) );
  NAND_GATE U9130 ( .I1(n8615), .I2(n8617), .O(n8311) );
  NAND3_GATE U9131 ( .I1(n8310), .I2(n8309), .I3(n8308), .O(n8619) );
  INV_GATE U9132 ( .I1(n8619), .O(n8618) );
  NAND_GATE U9133 ( .I1(n8615), .I2(n8618), .O(n8616) );
  NAND3_GATE U9134 ( .I1(n8312), .I2(n8311), .I3(n8616), .O(n8341) );
  NAND_GATE U9135 ( .I1(n8892), .I2(n8344), .O(n8313) );
  NAND_GATE U9136 ( .I1(n8341), .I2(n8313), .O(n8314) );
  NAND_GATE U9137 ( .I1(n8315), .I2(n8314), .O(n8634) );
  NAND_GATE U9138 ( .I1(n8882), .I2(n8637), .O(n8316) );
  NAND_GATE U9139 ( .I1(n8634), .I2(n8316), .O(n8317) );
  NAND_GATE U9140 ( .I1(n8643), .I2(n8642), .O(n8319) );
  NAND_GATE U9141 ( .I1(n8644), .I2(n8319), .O(n8320) );
  NAND_GATE U9142 ( .I1(n8655), .I2(n8322), .O(n8671) );
  NAND_GATE U9143 ( .I1(n8674), .I2(n8677), .O(n8323) );
  NAND_GATE U9144 ( .I1(n8671), .I2(n8323), .O(n8324) );
  NAND_GATE U9145 ( .I1(n8667), .I2(n8324), .O(n8687) );
  NAND_GATE U9146 ( .I1(n8689), .I2(n8693), .O(n8325) );
  NAND_GATE U9147 ( .I1(n8687), .I2(n8325), .O(n8326) );
  NAND_GATE U9148 ( .I1(n8684), .I2(n8326), .O(n8704) );
  NAND_GATE U9149 ( .I1(n8707), .I2(n8709), .O(n8327) );
  NAND_GATE U9150 ( .I1(n8704), .I2(n8327), .O(n8328) );
  NAND_GATE U9151 ( .I1(n8700), .I2(n8328), .O(n8720) );
  NAND_GATE U9152 ( .I1(n8718), .I2(n8725), .O(n8329) );
  NAND_GATE U9153 ( .I1(n8720), .I2(n8329), .O(n8330) );
  NAND_GATE U9154 ( .I1(n8716), .I2(n8330), .O(n8736) );
  NAND_GATE U9155 ( .I1(n8734), .I2(n8741), .O(n8331) );
  NAND_GATE U9156 ( .I1(n8736), .I2(n8331), .O(n8332) );
  NAND_GATE U9157 ( .I1(n8732), .I2(n8332), .O(n8753) );
  NAND_GATE U9158 ( .I1(n8751), .I2(n8758), .O(n8333) );
  NAND_GATE U9159 ( .I1(n8753), .I2(n8333), .O(n8334) );
  NAND_GATE U9160 ( .I1(n8748), .I2(n8334), .O(n8769) );
  NAND_GATE U9161 ( .I1(n8767), .I2(n8774), .O(n8335) );
  NAND_GATE U9162 ( .I1(n8769), .I2(n8335), .O(n8336) );
  NAND_GATE U9163 ( .I1(n8337), .I2(n285), .O(n8338) );
  AND_GATE U9164 ( .I1(n15328), .I2(n8338), .O(\A1[45] ) );
  NAND_GATE U9165 ( .I1(B[14]), .I2(A[31]), .O(n8789) );
  INV_GATE U9166 ( .I1(n8789), .O(n8763) );
  NAND_GATE U9167 ( .I1(B[14]), .I2(A[30]), .O(n8800) );
  INV_GATE U9168 ( .I1(n8800), .O(n8746) );
  NAND_GATE U9169 ( .I1(B[14]), .I2(A[29]), .O(n8811) );
  INV_GATE U9170 ( .I1(n8811), .O(n8730) );
  NAND_GATE U9171 ( .I1(B[14]), .I2(A[28]), .O(n8822) );
  INV_GATE U9172 ( .I1(n8822), .O(n8714) );
  NAND_GATE U9173 ( .I1(B[14]), .I2(A[27]), .O(n8833) );
  INV_GATE U9174 ( .I1(n8833), .O(n8698) );
  NAND_GATE U9175 ( .I1(B[14]), .I2(A[26]), .O(n8844) );
  INV_GATE U9176 ( .I1(n8844), .O(n8682) );
  NAND_GATE U9177 ( .I1(B[14]), .I2(A[25]), .O(n8858) );
  INV_GATE U9178 ( .I1(n8858), .O(n8665) );
  NAND_GATE U9179 ( .I1(B[14]), .I2(A[24]), .O(n8863) );
  INV_GATE U9180 ( .I1(n8863), .O(n8868) );
  NAND_GATE U9181 ( .I1(B[14]), .I2(A[23]), .O(n8887) );
  INV_GATE U9182 ( .I1(n8887), .O(n8640) );
  NAND_GATE U9183 ( .I1(B[14]), .I2(A[22]), .O(n8895) );
  INV_GATE U9184 ( .I1(n8895), .O(n8629) );
  NAND_GATE U9185 ( .I1(n8344), .I2(n8343), .O(n8339) );
  NAND_GATE U9186 ( .I1(n8340), .I2(n8339), .O(n8626) );
  NAND3_GATE U9187 ( .I1(n8340), .I2(n8341), .I3(n8342), .O(n8628) );
  NAND_GATE U9188 ( .I1(n8342), .I2(n8341), .O(n8345) );
  NAND_GATE U9189 ( .I1(n8345), .I2(n8339), .O(n8891) );
  NAND_GATE U9190 ( .I1(n919), .I2(n8625), .O(n8631) );
  NAND_GATE U9191 ( .I1(B[14]), .I2(A[21]), .O(n8912) );
  INV_GATE U9192 ( .I1(n8912), .O(n8622) );
  NAND_GATE U9193 ( .I1(B[14]), .I2(A[20]), .O(n8928) );
  INV_GATE U9194 ( .I1(n8928), .O(n8613) );
  NAND_GATE U9195 ( .I1(B[14]), .I2(A[18]), .O(n9235) );
  INV_GATE U9196 ( .I1(n9235), .O(n9169) );
  INV_GATE U9197 ( .I1(n8351), .O(n8349) );
  NAND4_GATE U9198 ( .I1(n8347), .I2(n8349), .I3(n990), .I4(n8346), .O(n8357)
         );
  OR_GATE U9199 ( .I1(n8350), .I2(n8348), .O(n8356) );
  NAND_GATE U9200 ( .I1(n8349), .I2(n8350), .O(n8353) );
  NAND3_GATE U9201 ( .I1(n8354), .I2(n8353), .I3(n8352), .O(n8355) );
  NAND3_GATE U9202 ( .I1(n8357), .I2(n8356), .I3(n8355), .O(n9170) );
  NAND_GATE U9203 ( .I1(n9169), .I2(n9172), .O(n8598) );
  NAND3_GATE U9204 ( .I1(n8359), .I2(n8358), .I3(n8365), .O(n8371) );
  NAND3_GATE U9205 ( .I1(n8361), .I2(n8360), .I3(n8359), .O(n8370) );
  NAND_GATE U9206 ( .I1(B[14]), .I2(A[17]), .O(n8938) );
  INV_GATE U9207 ( .I1(n8938), .O(n8594) );
  AND3_GATE U9208 ( .I1(n8371), .I2(n8370), .I3(n8594), .O(n8368) );
  NAND_GATE U9209 ( .I1(n8361), .I2(n8360), .O(n8362) );
  NAND_GATE U9210 ( .I1(n8363), .I2(n8362), .O(n8369) );
  INV_GATE U9211 ( .I1(n8364), .O(n8366) );
  NAND_GATE U9212 ( .I1(n8366), .I2(n8365), .O(n8373) );
  NAND_GATE U9213 ( .I1(n8368), .I2(n8367), .O(n8941) );
  NAND3_GATE U9214 ( .I1(n8371), .I2(n8370), .I3(n8369), .O(n8372) );
  NAND_GATE U9215 ( .I1(n8373), .I2(n8372), .O(n8939) );
  NAND_GATE U9216 ( .I1(B[14]), .I2(A[16]), .O(n9258) );
  INV_GATE U9217 ( .I1(n9258), .O(n9158) );
  NAND_GATE U9218 ( .I1(n8376), .I2(n8385), .O(n8380) );
  INV_GATE U9219 ( .I1(n8377), .O(n8379) );
  NAND3_GATE U9220 ( .I1(n8380), .I2(n8379), .I3(n8378), .O(n8392) );
  OR_GATE U9221 ( .I1(n8383), .I2(n8381), .O(n8391) );
  NAND_GATE U9222 ( .I1(n8384), .I2(n8385), .O(n8382) );
  NAND_GATE U9223 ( .I1(n8383), .I2(n8382), .O(n8389) );
  INV_GATE U9224 ( .I1(n8383), .O(n8386) );
  NAND3_GATE U9225 ( .I1(n8386), .I2(n8385), .I3(n8384), .O(n8388) );
  NAND3_GATE U9226 ( .I1(n8389), .I2(n8388), .I3(n8387), .O(n8390) );
  NAND3_GATE U9227 ( .I1(n8392), .I2(n8391), .I3(n8390), .O(n9159) );
  NAND_GATE U9228 ( .I1(n9158), .I2(n9161), .O(n8593) );
  NAND_GATE U9229 ( .I1(n8397), .I2(n770), .O(n8393) );
  NAND_GATE U9230 ( .I1(n8394), .I2(n8393), .O(n8586) );
  NAND_GATE U9231 ( .I1(n673), .I2(n8396), .O(n8398) );
  NAND_GATE U9232 ( .I1(n8398), .I2(n8393), .O(n8583) );
  NAND_GATE U9233 ( .I1(B[14]), .I2(A[15]), .O(n8950) );
  INV_GATE U9234 ( .I1(n8950), .O(n8589) );
  NAND3_GATE U9235 ( .I1(n8952), .I2(n8585), .I3(n8589), .O(n8953) );
  NAND_GATE U9236 ( .I1(B[14]), .I2(A[14]), .O(n9142) );
  INV_GATE U9237 ( .I1(n9142), .O(n9145) );
  NAND_GATE U9238 ( .I1(n772), .I2(n8405), .O(n8401) );
  NAND3_GATE U9239 ( .I1(n8401), .I2(n8400), .I3(n8399), .O(n8408) );
  OR_GATE U9240 ( .I1(n8403), .I2(n8402), .O(n8407) );
  OR_GATE U9241 ( .I1(n8405), .I2(n8404), .O(n8406) );
  NAND3_GATE U9242 ( .I1(n8408), .I2(n8407), .I3(n8406), .O(n9143) );
  NAND_GATE U9243 ( .I1(n9145), .I2(n9139), .O(n9148) );
  NAND_GATE U9244 ( .I1(B[14]), .I2(A[13]), .O(n9131) );
  INV_GATE U9245 ( .I1(n9131), .O(n8579) );
  INV_GATE U9246 ( .I1(n8419), .O(n8410) );
  NAND_GATE U9247 ( .I1(n8409), .I2(n8412), .O(n8417) );
  NAND_GATE U9248 ( .I1(n1329), .I2(n8419), .O(n8413) );
  NAND_GATE U9249 ( .I1(n8411), .I2(n8410), .O(n8412) );
  NAND_GATE U9250 ( .I1(n8413), .I2(n8412), .O(n8414) );
  NAND_GATE U9251 ( .I1(n8415), .I2(n8414), .O(n8416) );
  NAND_GATE U9252 ( .I1(n8417), .I2(n8416), .O(n8421) );
  NAND_GATE U9253 ( .I1(n8421), .I2(n8420), .O(n9128) );
  NAND_GATE U9254 ( .I1(n8579), .I2(n9128), .O(n9132) );
  NAND_GATE U9255 ( .I1(B[14]), .I2(A[12]), .O(n9116) );
  INV_GATE U9256 ( .I1(n9116), .O(n9112) );
  OR_GATE U9257 ( .I1(n8422), .I2(n8428), .O(n8425) );
  OR_GATE U9258 ( .I1(n8427), .I2(n8423), .O(n8424) );
  AND_GATE U9259 ( .I1(n8425), .I2(n8424), .O(n8433) );
  INV_GATE U9260 ( .I1(n8428), .O(n8426) );
  NAND_GATE U9261 ( .I1(n8426), .I2(n8427), .O(n8430) );
  NAND_GATE U9262 ( .I1(n8428), .I2(n166), .O(n8429) );
  NAND3_GATE U9263 ( .I1(n8431), .I2(n8430), .I3(n8429), .O(n8432) );
  NAND_GATE U9264 ( .I1(n8433), .I2(n8432), .O(n9113) );
  NAND_GATE U9265 ( .I1(n9112), .I2(n1204), .O(n9119) );
  NAND_GATE U9266 ( .I1(B[14]), .I2(A[11]), .O(n8969) );
  INV_GATE U9267 ( .I1(n8969), .O(n8575) );
  NAND_GATE U9268 ( .I1(n8435), .I2(n8434), .O(n8436) );
  NAND_GATE U9269 ( .I1(n8437), .I2(n8436), .O(n8440) );
  INV_GATE U9270 ( .I1(n8438), .O(n8439) );
  NAND3_GATE U9271 ( .I1(n8441), .I2(n8440), .I3(n8439), .O(n8452) );
  OR_GATE U9272 ( .I1(n8442), .I2(n8446), .O(n8451) );
  INV_GATE U9273 ( .I1(n8446), .O(n8443) );
  NAND3_GATE U9274 ( .I1(n8444), .I2(n8436), .I3(n8443), .O(n8449) );
  NAND_GATE U9275 ( .I1(n8444), .I2(n8436), .O(n8445) );
  NAND_GATE U9276 ( .I1(n8446), .I2(n8445), .O(n8448) );
  NAND3_GATE U9277 ( .I1(n8449), .I2(n8448), .I3(n8447), .O(n8450) );
  NAND_GATE U9278 ( .I1(B[14]), .I2(A[10]), .O(n8979) );
  INV_GATE U9279 ( .I1(n8979), .O(n8974) );
  NAND_GATE U9280 ( .I1(n746), .I2(n8974), .O(n8972) );
  NAND_GATE U9281 ( .I1(B[14]), .I2(A[9]), .O(n8990) );
  INV_GATE U9282 ( .I1(n8990), .O(n8558) );
  OR_GATE U9283 ( .I1(n8453), .I2(n8458), .O(n8456) );
  OR_GATE U9284 ( .I1(n8457), .I2(n8454), .O(n8455) );
  NAND_GATE U9285 ( .I1(n970), .I2(n8457), .O(n8461) );
  NAND3_GATE U9286 ( .I1(n8461), .I2(n8460), .I3(n8459), .O(n8462) );
  NAND_GATE U9287 ( .I1(B[14]), .I2(A[8]), .O(n9098) );
  INV_GATE U9288 ( .I1(n9098), .O(n9094) );
  NAND_GATE U9289 ( .I1(B[14]), .I2(A[7]), .O(n9000) );
  INV_GATE U9290 ( .I1(n9000), .O(n8545) );
  OR_GATE U9291 ( .I1(n8463), .I2(n8468), .O(n8466) );
  OR_GATE U9292 ( .I1(n8467), .I2(n8464), .O(n8465) );
  AND_GATE U9293 ( .I1(n8466), .I2(n8465), .O(n8473) );
  NAND_GATE U9294 ( .I1(n1043), .I2(n8467), .O(n8471) );
  NAND3_GATE U9295 ( .I1(n8471), .I2(n8470), .I3(n8469), .O(n8472) );
  NAND_GATE U9296 ( .I1(n8473), .I2(n8472), .O(n9075) );
  INV_GATE U9297 ( .I1(n9075), .O(n9078) );
  NAND_GATE U9298 ( .I1(B[14]), .I2(A[6]), .O(n9082) );
  INV_GATE U9299 ( .I1(n9082), .O(n9076) );
  NAND_GATE U9300 ( .I1(n9078), .I2(n9076), .O(n9072) );
  NAND_GATE U9301 ( .I1(B[14]), .I2(A[5]), .O(n9011) );
  INV_GATE U9302 ( .I1(n9011), .O(n8526) );
  OR_GATE U9303 ( .I1(n8474), .I2(n8479), .O(n8477) );
  OR_GATE U9304 ( .I1(n8478), .I2(n8475), .O(n8476) );
  AND_GATE U9305 ( .I1(n8477), .I2(n8476), .O(n8484) );
  NAND_GATE U9306 ( .I1(n1166), .I2(n8478), .O(n8482) );
  NAND3_GATE U9307 ( .I1(n8482), .I2(n8481), .I3(n8480), .O(n8483) );
  NAND_GATE U9308 ( .I1(n8484), .I2(n8483), .O(n9056) );
  INV_GATE U9309 ( .I1(n9056), .O(n9059) );
  NAND_GATE U9310 ( .I1(B[14]), .I2(A[4]), .O(n9063) );
  INV_GATE U9311 ( .I1(n9063), .O(n9057) );
  NAND_GATE U9312 ( .I1(n9059), .I2(n9057), .O(n9053) );
  NAND_GATE U9313 ( .I1(B[14]), .I2(A[3]), .O(n9022) );
  INV_GATE U9314 ( .I1(n9022), .O(n8507) );
  NAND_GATE U9315 ( .I1(B[14]), .I2(A[2]), .O(n9036) );
  INV_GATE U9316 ( .I1(n9036), .O(n9030) );
  NAND_GATE U9317 ( .I1(n1380), .I2(A[0]), .O(n8485) );
  NAND_GATE U9318 ( .I1(n14781), .I2(n8485), .O(n8486) );
  NAND_GATE U9319 ( .I1(B[16]), .I2(n8486), .O(n8490) );
  NAND_GATE U9320 ( .I1(n1381), .I2(A[1]), .O(n8487) );
  NAND_GATE U9321 ( .I1(n14784), .I2(n8487), .O(n8488) );
  NAND_GATE U9322 ( .I1(n1379), .I2(n8488), .O(n8489) );
  NAND_GATE U9323 ( .I1(n8490), .I2(n8489), .O(n9032) );
  NAND_GATE U9324 ( .I1(n9030), .I2(n9032), .O(n9027) );
  NAND3_GATE U9325 ( .I1(B[14]), .I2(n1379), .I3(n1196), .O(n9028) );
  INV_GATE U9326 ( .I1(n9028), .O(n9031) );
  INV_GATE U9327 ( .I1(n9032), .O(n9029) );
  NAND_GATE U9328 ( .I1(n9036), .I2(n9029), .O(n8491) );
  NAND_GATE U9329 ( .I1(n9031), .I2(n8491), .O(n8492) );
  NAND_GATE U9330 ( .I1(n9027), .I2(n8492), .O(n9021) );
  NAND_GATE U9331 ( .I1(n8507), .I2(n9021), .O(n9017) );
  OR_GATE U9332 ( .I1(n8494), .I2(n8493), .O(n8506) );
  NAND_GATE U9333 ( .I1(n8495), .I2(n8494), .O(n8500) );
  NAND_GATE U9334 ( .I1(n8496), .I2(n8500), .O(n8504) );
  NAND_GATE U9335 ( .I1(n8498), .I2(n8497), .O(n8499) );
  NAND_GATE U9336 ( .I1(n8500), .I2(n8499), .O(n8501) );
  NAND_GATE U9337 ( .I1(n8502), .I2(n8501), .O(n8503) );
  NAND_GATE U9338 ( .I1(n8504), .I2(n8503), .O(n8505) );
  NAND_GATE U9339 ( .I1(n8506), .I2(n8505), .O(n9020) );
  NAND_GATE U9340 ( .I1(n9021), .I2(n9020), .O(n8508) );
  NAND_GATE U9341 ( .I1(n8507), .I2(n9020), .O(n9016) );
  NAND3_GATE U9342 ( .I1(n9017), .I2(n8508), .I3(n9016), .O(n9058) );
  NAND_GATE U9343 ( .I1(n9056), .I2(n9063), .O(n8509) );
  NAND_GATE U9344 ( .I1(n9058), .I2(n8509), .O(n8510) );
  NAND_GATE U9345 ( .I1(n9053), .I2(n8510), .O(n9010) );
  NAND_GATE U9346 ( .I1(n8526), .I2(n9010), .O(n9006) );
  INV_GATE U9347 ( .I1(n8511), .O(n8512) );
  NAND_GATE U9348 ( .I1(n8512), .I2(n8516), .O(n8525) );
  INV_GATE U9349 ( .I1(n8516), .O(n8513) );
  NAND_GATE U9350 ( .I1(n8514), .I2(n8513), .O(n8519) );
  NAND_GATE U9351 ( .I1(n8515), .I2(n8519), .O(n8523) );
  NAND_GATE U9352 ( .I1(n8517), .I2(n8516), .O(n8518) );
  NAND_GATE U9353 ( .I1(n8519), .I2(n8518), .O(n8520) );
  NAND_GATE U9354 ( .I1(n8521), .I2(n8520), .O(n8522) );
  NAND_GATE U9355 ( .I1(n8523), .I2(n8522), .O(n8524) );
  NAND_GATE U9356 ( .I1(n8525), .I2(n8524), .O(n9009) );
  NAND_GATE U9357 ( .I1(n9010), .I2(n9009), .O(n8527) );
  NAND_GATE U9358 ( .I1(n8526), .I2(n9009), .O(n9005) );
  NAND3_GATE U9359 ( .I1(n9006), .I2(n8527), .I3(n9005), .O(n9077) );
  NAND_GATE U9360 ( .I1(n9075), .I2(n9082), .O(n8528) );
  NAND_GATE U9361 ( .I1(n9077), .I2(n8528), .O(n8529) );
  NAND_GATE U9362 ( .I1(n9072), .I2(n8529), .O(n8999) );
  NAND_GATE U9363 ( .I1(n8545), .I2(n8999), .O(n8995) );
  INV_GATE U9364 ( .I1(n8530), .O(n8531) );
  NAND_GATE U9365 ( .I1(n8531), .I2(n8535), .O(n8544) );
  INV_GATE U9366 ( .I1(n8535), .O(n8532) );
  NAND_GATE U9367 ( .I1(n8533), .I2(n8532), .O(n8538) );
  NAND_GATE U9368 ( .I1(n8534), .I2(n8538), .O(n8542) );
  NAND_GATE U9369 ( .I1(n8536), .I2(n8535), .O(n8537) );
  NAND_GATE U9370 ( .I1(n8538), .I2(n8537), .O(n8539) );
  NAND_GATE U9371 ( .I1(n8540), .I2(n8539), .O(n8541) );
  NAND_GATE U9372 ( .I1(n8542), .I2(n8541), .O(n8543) );
  NAND_GATE U9373 ( .I1(n8544), .I2(n8543), .O(n8998) );
  NAND_GATE U9374 ( .I1(n8545), .I2(n8998), .O(n8994) );
  NAND_GATE U9375 ( .I1(n9093), .I2(n9098), .O(n8546) );
  NAND_GATE U9376 ( .I1(n9095), .I2(n8546), .O(n8547) );
  NAND_GATE U9377 ( .I1(n9091), .I2(n8547), .O(n8989) );
  NAND_GATE U9378 ( .I1(n8558), .I2(n8989), .O(n8985) );
  INV_GATE U9379 ( .I1(n8548), .O(n8549) );
  NAND_GATE U9380 ( .I1(n8549), .I2(n8550), .O(n8557) );
  NAND_GATE U9381 ( .I1(n731), .I2(n8552), .O(n8555) );
  NAND_GATE U9382 ( .I1(n874), .I2(n8550), .O(n8551) );
  NAND_GATE U9383 ( .I1(n8555), .I2(n8554), .O(n8556) );
  NAND_GATE U9384 ( .I1(n8557), .I2(n8556), .O(n8988) );
  NAND_GATE U9385 ( .I1(n8989), .I2(n8988), .O(n8559) );
  NAND_GATE U9386 ( .I1(n8558), .I2(n8988), .O(n8984) );
  NAND3_GATE U9387 ( .I1(n8985), .I2(n8559), .I3(n8984), .O(n8975) );
  NAND_GATE U9388 ( .I1(n8975), .I2(n8560), .O(n8561) );
  NAND_GATE U9389 ( .I1(n8972), .I2(n8561), .O(n8966) );
  NAND_GATE U9390 ( .I1(n8575), .I2(n8966), .O(n8962) );
  INV_GATE U9391 ( .I1(n8571), .O(n8565) );
  NAND_GATE U9392 ( .I1(n8566), .I2(n8565), .O(n8562) );
  NAND_GATE U9393 ( .I1(n8563), .I2(n8562), .O(n8569) );
  NAND_GATE U9394 ( .I1(n8569), .I2(n8568), .O(n8574) );
  INV_GATE U9395 ( .I1(n8570), .O(n8572) );
  NAND_GATE U9396 ( .I1(n8572), .I2(n8571), .O(n8573) );
  NAND_GATE U9397 ( .I1(n8574), .I2(n8573), .O(n8965) );
  NAND_GATE U9398 ( .I1(n8966), .I2(n8965), .O(n8576) );
  NAND_GATE U9399 ( .I1(n8575), .I2(n8965), .O(n8961) );
  NAND3_GATE U9400 ( .I1(n8962), .I2(n8576), .I3(n8961), .O(n9120) );
  NAND_GATE U9401 ( .I1(n9116), .I2(n9113), .O(n8577) );
  NAND_GATE U9402 ( .I1(n9120), .I2(n8577), .O(n8578) );
  NAND_GATE U9403 ( .I1(n9119), .I2(n8578), .O(n9133) );
  NAND_GATE U9404 ( .I1(n9128), .I2(n9133), .O(n8580) );
  NAND_GATE U9405 ( .I1(n8579), .I2(n9133), .O(n9126) );
  NAND3_GATE U9406 ( .I1(n9132), .I2(n8580), .I3(n9126), .O(n9149) );
  NAND_GATE U9407 ( .I1(n9142), .I2(n9143), .O(n8581) );
  NAND_GATE U9408 ( .I1(n9149), .I2(n8581), .O(n8582) );
  NAND_GATE U9409 ( .I1(n9148), .I2(n8582), .O(n8951) );
  NAND_GATE U9410 ( .I1(n8584), .I2(n8583), .O(n8585) );
  NAND_GATE U9411 ( .I1(n8586), .I2(n8585), .O(n8587) );
  NAND_GATE U9412 ( .I1(n8588), .I2(n8587), .O(n8946) );
  NAND_GATE U9413 ( .I1(n8951), .I2(n8946), .O(n8590) );
  NAND_GATE U9414 ( .I1(n8589), .I2(n8951), .O(n8947) );
  NAND_GATE U9415 ( .I1(n9258), .I2(n9159), .O(n8591) );
  NAND_GATE U9416 ( .I1(n9160), .I2(n8591), .O(n8592) );
  NAND_GATE U9417 ( .I1(n8593), .I2(n8592), .O(n8942) );
  NAND_GATE U9418 ( .I1(n8939), .I2(n8942), .O(n8595) );
  NAND_GATE U9419 ( .I1(n8594), .I2(n8942), .O(n8940) );
  NAND_GATE U9420 ( .I1(n9235), .I2(n9170), .O(n8596) );
  NAND_GATE U9421 ( .I1(n9171), .I2(n8596), .O(n8597) );
  NAND_GATE U9422 ( .I1(n8598), .I2(n8597), .O(n9185) );
  NAND_GATE U9423 ( .I1(n8603), .I2(n807), .O(n8600) );
  NAND_GATE U9424 ( .I1(n257), .I2(n8601), .O(n8599) );
  NAND_GATE U9425 ( .I1(n8600), .I2(n8599), .O(n9178) );
  NAND_GATE U9426 ( .I1(n9182), .I2(n9180), .O(n8604) );
  NAND3_GATE U9427 ( .I1(n8603), .I2(n8602), .I3(n807), .O(n9181) );
  NAND_GATE U9428 ( .I1(n8604), .I2(n9181), .O(n9192) );
  NAND_GATE U9429 ( .I1(n9185), .I2(n9192), .O(n8606) );
  NAND_GATE U9430 ( .I1(B[14]), .I2(A[19]), .O(n9186) );
  INV_GATE U9431 ( .I1(n9186), .O(n9189) );
  NAND_GATE U9432 ( .I1(n9189), .I2(n9192), .O(n8605) );
  NAND_GATE U9433 ( .I1(n9189), .I2(n9185), .O(n9191) );
  NAND3_GATE U9434 ( .I1(n8606), .I2(n8605), .I3(n9191), .O(n8929) );
  NAND_GATE U9435 ( .I1(n8613), .I2(n8929), .O(n8931) );
  NAND3_GATE U9436 ( .I1(n8607), .I2(n252), .I3(n8609), .O(n8922) );
  NAND_GATE U9437 ( .I1(n8607), .I2(n8611), .O(n8920) );
  NAND_GATE U9438 ( .I1(n8608), .I2(n261), .O(n8611) );
  NAND_GATE U9439 ( .I1(n8609), .I2(n252), .O(n8610) );
  NAND_GATE U9440 ( .I1(n8611), .I2(n8610), .O(n8918) );
  NAND_GATE U9441 ( .I1(n8920), .I2(n8925), .O(n8612) );
  NAND_GATE U9442 ( .I1(n8922), .I2(n8612), .O(n8932) );
  NAND_GATE U9443 ( .I1(n8929), .I2(n8932), .O(n8614) );
  NAND3_GATE U9444 ( .I1(n8931), .I2(n8930), .I3(n8614), .O(n8909) );
  NAND_GATE U9445 ( .I1(n8622), .I2(n8909), .O(n8916) );
  NAND_GATE U9446 ( .I1(n8615), .I2(n8620), .O(n8915) );
  INV_GATE U9447 ( .I1(n8915), .O(n8906) );
  NAND_GATE U9448 ( .I1(n8906), .I2(n8917), .O(n8623) );
  NAND_GATE U9449 ( .I1(n8618), .I2(n8617), .O(n8621) );
  NAND_GATE U9450 ( .I1(n8619), .I2(n590), .O(n8620) );
  NAND_GATE U9451 ( .I1(n8621), .I2(n8620), .O(n8913) );
  NAND3_GATE U9452 ( .I1(n8622), .I2(n8623), .I3(n8907), .O(n8905) );
  NAND3_GATE U9453 ( .I1(n8909), .I2(n8623), .I3(n8907), .O(n8624) );
  NAND3_GATE U9454 ( .I1(n8916), .I2(n8905), .I3(n8624), .O(n8898) );
  NAND_GATE U9455 ( .I1(n8892), .I2(n8891), .O(n8625) );
  NAND_GATE U9456 ( .I1(n8626), .I2(n8625), .O(n8627) );
  NAND_GATE U9457 ( .I1(n8628), .I2(n8627), .O(n8900) );
  NAND_GATE U9458 ( .I1(n8898), .I2(n8900), .O(n8630) );
  NAND_GATE U9459 ( .I1(n8629), .I2(n8898), .O(n8901) );
  NAND3_GATE U9460 ( .I1(n8631), .I2(n8630), .I3(n8901), .O(n8886) );
  NAND_GATE U9461 ( .I1(n8640), .I2(n8886), .O(n8875) );
  NAND3_GATE U9462 ( .I1(n8633), .I2(n8634), .I3(n8635), .O(n8880) );
  INV_GATE U9463 ( .I1(n8634), .O(n8636) );
  NAND_GATE U9464 ( .I1(n8637), .I2(n8636), .O(n8632) );
  NAND_GATE U9465 ( .I1(n8633), .I2(n8632), .O(n8879) );
  NAND_GATE U9466 ( .I1(n8635), .I2(n8634), .O(n8638) );
  NAND_GATE U9467 ( .I1(n8638), .I2(n8632), .O(n8881) );
  NAND_GATE U9468 ( .I1(n8879), .I2(n8883), .O(n8639) );
  NAND_GATE U9469 ( .I1(n8880), .I2(n8639), .O(n8876) );
  NAND_GATE U9470 ( .I1(n8640), .I2(n8876), .O(n8874) );
  NAND_GATE U9471 ( .I1(n8886), .I2(n8876), .O(n8641) );
  NAND3_GATE U9472 ( .I1(n8875), .I2(n8874), .I3(n8641), .O(n8862) );
  NAND_GATE U9473 ( .I1(n8868), .I2(n8862), .O(n8869) );
  NAND3_GATE U9474 ( .I1(n8647), .I2(n8644), .I3(n8645), .O(n8652) );
  NAND_GATE U9475 ( .I1(n8642), .I2(n175), .O(n8646) );
  NAND3_GATE U9476 ( .I1(n8647), .I2(n8652), .I3(n8646), .O(n8867) );
  NAND3_GATE U9477 ( .I1(n8642), .I2(n175), .I3(n8643), .O(n8648) );
  NAND3_GATE U9478 ( .I1(n8645), .I2(n8644), .I3(n8643), .O(n8650) );
  NAND3_GATE U9479 ( .I1(n8868), .I2(n8867), .I3(n1000), .O(n8654) );
  NAND_GATE U9480 ( .I1(n8647), .I2(n8646), .O(n8649) );
  NAND3_GATE U9481 ( .I1(n8650), .I2(n8649), .I3(n8648), .O(n8651) );
  NAND_GATE U9482 ( .I1(n8652), .I2(n8651), .O(n8870) );
  NAND_GATE U9483 ( .I1(n8862), .I2(n8870), .O(n8653) );
  NAND3_GATE U9484 ( .I1(n8869), .I2(n8654), .I3(n8653), .O(n8856) );
  NAND_GATE U9485 ( .I1(n8665), .I2(n8856), .O(n8850) );
  NAND_GATE U9486 ( .I1(n8659), .I2(n791), .O(n8656) );
  NAND_GATE U9487 ( .I1(n8657), .I2(n8656), .O(n8664) );
  NAND_GATE U9488 ( .I1(n8660), .I2(n8656), .O(n8661) );
  NAND_GATE U9489 ( .I1(n8662), .I2(n8661), .O(n8663) );
  NAND_GATE U9490 ( .I1(n8664), .I2(n8663), .O(n8855) );
  NAND_GATE U9491 ( .I1(n8857), .I2(n8855), .O(n8853) );
  NAND_GATE U9492 ( .I1(n8665), .I2(n8853), .O(n8849) );
  NAND_GATE U9493 ( .I1(n8856), .I2(n8853), .O(n8666) );
  NAND3_GATE U9494 ( .I1(n8850), .I2(n8849), .I3(n8666), .O(n8843) );
  NAND_GATE U9495 ( .I1(n8682), .I2(n8843), .O(n8839) );
  INV_GATE U9496 ( .I1(n8667), .O(n8668) );
  NAND_GATE U9497 ( .I1(n8668), .I2(n8671), .O(n8681) );
  INV_GATE U9498 ( .I1(n8671), .O(n8673) );
  NAND_GATE U9499 ( .I1(n8674), .I2(n8673), .O(n8669) );
  NAND_GATE U9500 ( .I1(n8670), .I2(n8669), .O(n8679) );
  NAND_GATE U9501 ( .I1(n8672), .I2(n8671), .O(n8675) );
  NAND_GATE U9502 ( .I1(n8675), .I2(n8669), .O(n8676) );
  NAND_GATE U9503 ( .I1(n8677), .I2(n8676), .O(n8678) );
  NAND_GATE U9504 ( .I1(n8679), .I2(n8678), .O(n8680) );
  NAND_GATE U9505 ( .I1(n8681), .I2(n8680), .O(n8842) );
  NAND_GATE U9506 ( .I1(n8843), .I2(n8842), .O(n8683) );
  NAND3_GATE U9507 ( .I1(n8839), .I2(n8838), .I3(n8683), .O(n8832) );
  NAND_GATE U9508 ( .I1(n8698), .I2(n8832), .O(n8828) );
  INV_GATE U9509 ( .I1(n8684), .O(n8685) );
  NAND_GATE U9510 ( .I1(n8685), .I2(n8687), .O(n8697) );
  NAND_GATE U9511 ( .I1(n8686), .I2(n8690), .O(n8695) );
  NAND_GATE U9512 ( .I1(n831), .I2(n8687), .O(n8691) );
  NAND_GATE U9513 ( .I1(n8689), .I2(n8688), .O(n8690) );
  NAND_GATE U9514 ( .I1(n8691), .I2(n8690), .O(n8692) );
  NAND_GATE U9515 ( .I1(n8693), .I2(n8692), .O(n8694) );
  NAND_GATE U9516 ( .I1(n8695), .I2(n8694), .O(n8696) );
  NAND_GATE U9517 ( .I1(n8697), .I2(n8696), .O(n8831) );
  NAND_GATE U9518 ( .I1(n8832), .I2(n8831), .O(n8699) );
  NAND3_GATE U9519 ( .I1(n8828), .I2(n8827), .I3(n8699), .O(n8821) );
  NAND_GATE U9520 ( .I1(n8714), .I2(n8821), .O(n8817) );
  INV_GATE U9521 ( .I1(n8700), .O(n8701) );
  NAND_GATE U9522 ( .I1(n8701), .I2(n8704), .O(n8713) );
  INV_GATE U9523 ( .I1(n8704), .O(n8706) );
  NAND_GATE U9524 ( .I1(n8707), .I2(n8706), .O(n8702) );
  NAND_GATE U9525 ( .I1(n8703), .I2(n8702), .O(n8711) );
  NAND_GATE U9526 ( .I1(n8705), .I2(n8704), .O(n8708) );
  NAND_GATE U9527 ( .I1(n8711), .I2(n8710), .O(n8712) );
  NAND_GATE U9528 ( .I1(n8713), .I2(n8712), .O(n8820) );
  NAND_GATE U9529 ( .I1(n8821), .I2(n8820), .O(n8715) );
  NAND3_GATE U9530 ( .I1(n8817), .I2(n8816), .I3(n8715), .O(n8810) );
  NAND_GATE U9531 ( .I1(n8730), .I2(n8810), .O(n8806) );
  INV_GATE U9532 ( .I1(n8716), .O(n8717) );
  NAND_GATE U9533 ( .I1(n8717), .I2(n8720), .O(n8729) );
  NAND_GATE U9534 ( .I1(n8719), .I2(n8723), .O(n8727) );
  NAND_GATE U9535 ( .I1(n8721), .I2(n8720), .O(n8722) );
  NAND_GATE U9536 ( .I1(n8723), .I2(n8722), .O(n8724) );
  NAND_GATE U9537 ( .I1(n8725), .I2(n8724), .O(n8726) );
  NAND_GATE U9538 ( .I1(n8727), .I2(n8726), .O(n8728) );
  NAND_GATE U9539 ( .I1(n8729), .I2(n8728), .O(n8809) );
  NAND_GATE U9540 ( .I1(n8810), .I2(n8809), .O(n8731) );
  NAND3_GATE U9541 ( .I1(n8806), .I2(n8805), .I3(n8731), .O(n8799) );
  NAND_GATE U9542 ( .I1(n8746), .I2(n8799), .O(n8795) );
  INV_GATE U9543 ( .I1(n8732), .O(n8733) );
  NAND_GATE U9544 ( .I1(n8733), .I2(n8736), .O(n8745) );
  NAND_GATE U9545 ( .I1(n8735), .I2(n8739), .O(n8743) );
  NAND_GATE U9546 ( .I1(n8737), .I2(n8736), .O(n8738) );
  NAND_GATE U9547 ( .I1(n8739), .I2(n8738), .O(n8740) );
  NAND_GATE U9548 ( .I1(n8741), .I2(n8740), .O(n8742) );
  NAND_GATE U9549 ( .I1(n8743), .I2(n8742), .O(n8744) );
  NAND_GATE U9550 ( .I1(n8745), .I2(n8744), .O(n8798) );
  NAND_GATE U9551 ( .I1(n8799), .I2(n8798), .O(n8747) );
  NAND3_GATE U9552 ( .I1(n8795), .I2(n8794), .I3(n8747), .O(n8788) );
  NAND_GATE U9553 ( .I1(n8763), .I2(n8788), .O(n8784) );
  INV_GATE U9554 ( .I1(n8748), .O(n8749) );
  NAND_GATE U9555 ( .I1(n8749), .I2(n8753), .O(n8762) );
  INV_GATE U9556 ( .I1(n8753), .O(n8750) );
  NAND_GATE U9557 ( .I1(n8751), .I2(n8750), .O(n8756) );
  NAND_GATE U9558 ( .I1(n8752), .I2(n8756), .O(n8760) );
  NAND_GATE U9559 ( .I1(n8754), .I2(n8753), .O(n8755) );
  NAND_GATE U9560 ( .I1(n8756), .I2(n8755), .O(n8757) );
  NAND_GATE U9561 ( .I1(n8758), .I2(n8757), .O(n8759) );
  NAND_GATE U9562 ( .I1(n8760), .I2(n8759), .O(n8761) );
  NAND_GATE U9563 ( .I1(n8762), .I2(n8761), .O(n8787) );
  NAND_GATE U9564 ( .I1(n8763), .I2(n8787), .O(n8783) );
  NAND_GATE U9565 ( .I1(n8788), .I2(n8787), .O(n8764) );
  NAND3_GATE U9566 ( .I1(n8784), .I2(n8783), .I3(n8764), .O(n15330) );
  INV_GATE U9567 ( .I1(n15330), .O(n8779) );
  INV_GATE U9568 ( .I1(n8765), .O(n8766) );
  NAND_GATE U9569 ( .I1(n8766), .I2(n8769), .O(n8778) );
  NAND_GATE U9570 ( .I1(n8768), .I2(n8772), .O(n8776) );
  NAND_GATE U9571 ( .I1(n8770), .I2(n8769), .O(n8771) );
  NAND_GATE U9572 ( .I1(n8772), .I2(n8771), .O(n8773) );
  NAND_GATE U9573 ( .I1(n8774), .I2(n8773), .O(n8775) );
  NAND_GATE U9574 ( .I1(n8776), .I2(n8775), .O(n8777) );
  NAND_GATE U9575 ( .I1(n8778), .I2(n8777), .O(n15329) );
  NAND_GATE U9576 ( .I1(n8779), .I2(n15329), .O(n8782) );
  INV_GATE U9577 ( .I1(n15329), .O(n8780) );
  NAND_GATE U9578 ( .I1(n15330), .I2(n8780), .O(n8781) );
  NAND_GATE U9579 ( .I1(n8782), .I2(n8781), .O(\A1[44] ) );
  OR_GATE U9580 ( .I1(n8783), .I2(n8788), .O(n8786) );
  OR_GATE U9581 ( .I1(n8787), .I2(n8784), .O(n8785) );
  AND_GATE U9582 ( .I1(n8786), .I2(n8785), .O(n8793) );
  NAND_GATE U9583 ( .I1(n912), .I2(n8787), .O(n8791) );
  NAND3_GATE U9584 ( .I1(n8791), .I2(n8790), .I3(n8789), .O(n8792) );
  NAND_GATE U9585 ( .I1(n8793), .I2(n8792), .O(n9224) );
  OR_GATE U9586 ( .I1(n8794), .I2(n8799), .O(n8797) );
  OR_GATE U9587 ( .I1(n8798), .I2(n8795), .O(n8796) );
  AND_GATE U9588 ( .I1(n8797), .I2(n8796), .O(n8804) );
  NAND_GATE U9589 ( .I1(n95), .I2(n8798), .O(n8802) );
  NAND3_GATE U9590 ( .I1(n8802), .I2(n8801), .I3(n8800), .O(n8803) );
  NAND_GATE U9591 ( .I1(n8804), .I2(n8803), .O(n9635) );
  NAND_GATE U9592 ( .I1(B[13]), .I2(A[31]), .O(n9642) );
  INV_GATE U9593 ( .I1(n9642), .O(n9636) );
  NAND_GATE U9594 ( .I1(n9638), .I2(n9636), .O(n9633) );
  OR_GATE U9595 ( .I1(n8805), .I2(n8810), .O(n8808) );
  OR_GATE U9596 ( .I1(n8809), .I2(n8806), .O(n8807) );
  AND_GATE U9597 ( .I1(n8808), .I2(n8807), .O(n8815) );
  NAND_GATE U9598 ( .I1(n80), .I2(n8809), .O(n8813) );
  NAND3_GATE U9599 ( .I1(n8813), .I2(n8812), .I3(n8811), .O(n8814) );
  NAND_GATE U9600 ( .I1(n8815), .I2(n8814), .O(n9619) );
  NAND_GATE U9601 ( .I1(B[13]), .I2(A[30]), .O(n9626) );
  INV_GATE U9602 ( .I1(n9626), .O(n9620) );
  NAND_GATE U9603 ( .I1(n9622), .I2(n9620), .O(n9617) );
  OR_GATE U9604 ( .I1(n8820), .I2(n8817), .O(n8818) );
  AND_GATE U9605 ( .I1(n8819), .I2(n8818), .O(n8826) );
  NAND_GATE U9606 ( .I1(n888), .I2(n8820), .O(n8824) );
  NAND3_GATE U9607 ( .I1(n8824), .I2(n8823), .I3(n8822), .O(n8825) );
  NAND_GATE U9608 ( .I1(n8826), .I2(n8825), .O(n9607) );
  NAND_GATE U9609 ( .I1(B[13]), .I2(A[29]), .O(n9610) );
  INV_GATE U9610 ( .I1(n9610), .O(n9604) );
  NAND_GATE U9611 ( .I1(n617), .I2(n9604), .O(n9601) );
  OR_GATE U9612 ( .I1(n8827), .I2(n8832), .O(n8830) );
  OR_GATE U9613 ( .I1(n8831), .I2(n8828), .O(n8829) );
  AND_GATE U9614 ( .I1(n8830), .I2(n8829), .O(n8837) );
  NAND_GATE U9615 ( .I1(n9), .I2(n8831), .O(n8835) );
  NAND3_GATE U9616 ( .I1(n8835), .I2(n8834), .I3(n8833), .O(n8836) );
  NAND_GATE U9617 ( .I1(n8837), .I2(n8836), .O(n9591) );
  NAND_GATE U9618 ( .I1(B[13]), .I2(A[28]), .O(n9594) );
  INV_GATE U9619 ( .I1(n9594), .O(n9589) );
  NAND_GATE U9620 ( .I1(n830), .I2(n9589), .O(n9586) );
  OR_GATE U9621 ( .I1(n8842), .I2(n8839), .O(n8840) );
  AND_GATE U9622 ( .I1(n8841), .I2(n8840), .O(n8848) );
  NAND_GATE U9623 ( .I1(n884), .I2(n8842), .O(n8846) );
  NAND3_GATE U9624 ( .I1(n8846), .I2(n8845), .I3(n8844), .O(n8847) );
  NAND_GATE U9625 ( .I1(n8848), .I2(n8847), .O(n9578) );
  INV_GATE U9626 ( .I1(n9578), .O(n9576) );
  NAND_GATE U9627 ( .I1(B[13]), .I2(A[27]), .O(n9580) );
  INV_GATE U9628 ( .I1(n9580), .O(n9574) );
  NAND_GATE U9629 ( .I1(n9576), .I2(n9574), .O(n9572) );
  OR_GATE U9630 ( .I1(n8849), .I2(n8856), .O(n8852) );
  OR_GATE U9631 ( .I1(n8853), .I2(n8850), .O(n8851) );
  INV_GATE U9632 ( .I1(n8856), .O(n8854) );
  NAND_GATE U9633 ( .I1(n8854), .I2(n8853), .O(n8860) );
  NAND3_GATE U9634 ( .I1(n8857), .I2(n8856), .I3(n8855), .O(n8859) );
  NAND3_GATE U9635 ( .I1(n8860), .I2(n8859), .I3(n8858), .O(n8861) );
  NAND_GATE U9636 ( .I1(B[13]), .I2(A[26]), .O(n9567) );
  INV_GATE U9637 ( .I1(n9567), .O(n9562) );
  NAND_GATE U9638 ( .I1(n630), .I2(n9562), .O(n9560) );
  INV_GATE U9639 ( .I1(n8862), .O(n8866) );
  NAND_GATE U9640 ( .I1(n8866), .I2(n8870), .O(n8865) );
  NAND_GATE U9641 ( .I1(n8862), .I2(n130), .O(n8864) );
  NAND3_GATE U9642 ( .I1(n8865), .I2(n8864), .I3(n8863), .O(n8873) );
  NAND4_GATE U9643 ( .I1(n8868), .I2(n8867), .I3(n1000), .I4(n8866), .O(n8872)
         );
  OR_GATE U9644 ( .I1(n8870), .I2(n8869), .O(n8871) );
  NAND3_GATE U9645 ( .I1(n8873), .I2(n8872), .I3(n8871), .O(n9552) );
  INV_GATE U9646 ( .I1(n9552), .O(n9549) );
  NAND_GATE U9647 ( .I1(B[13]), .I2(A[25]), .O(n9550) );
  INV_GATE U9648 ( .I1(n9550), .O(n9547) );
  NAND_GATE U9649 ( .I1(B[13]), .I2(A[24]), .O(n9720) );
  INV_GATE U9650 ( .I1(n9720), .O(n9535) );
  OR_GATE U9651 ( .I1(n8876), .I2(n8875), .O(n8877) );
  NAND_GATE U9652 ( .I1(n8882), .I2(n8881), .O(n8883) );
  NAND_GATE U9653 ( .I1(n8884), .I2(n8883), .O(n8885) );
  NAND_GATE U9654 ( .I1(n8886), .I2(n8885), .O(n8888) );
  NAND3_GATE U9655 ( .I1(n8889), .I2(n8888), .I3(n8887), .O(n8890) );
  INV_GATE U9656 ( .I1(n9538), .O(n9537) );
  NAND_GATE U9657 ( .I1(n9535), .I2(n9537), .O(n9209) );
  NAND_GATE U9658 ( .I1(B[13]), .I2(A[23]), .O(n9522) );
  INV_GATE U9659 ( .I1(n9522), .O(n9521) );
  NAND_GATE U9660 ( .I1(n8893), .I2(n8625), .O(n8894) );
  OR_GATE U9661 ( .I1(n8894), .I2(n8898), .O(n8897) );
  NAND_GATE U9662 ( .I1(n8898), .I2(n8894), .O(n8896) );
  NAND3_GATE U9663 ( .I1(n8897), .I2(n8896), .I3(n8895), .O(n8904) );
  INV_GATE U9664 ( .I1(n8898), .O(n8899) );
  NAND3_GATE U9665 ( .I1(n8899), .I2(n8625), .I3(n919), .O(n8903) );
  OR_GATE U9666 ( .I1(n8901), .I2(n8900), .O(n8902) );
  NAND3_GATE U9667 ( .I1(n8904), .I2(n8903), .I3(n8902), .O(n9524) );
  NAND_GATE U9668 ( .I1(n9521), .I2(n4), .O(n9528) );
  NAND_GATE U9669 ( .I1(n8914), .I2(n8913), .O(n8907) );
  NAND3_GATE U9670 ( .I1(n737), .I2(n8623), .I3(n8907), .O(n8911) );
  NAND_GATE U9671 ( .I1(n8623), .I2(n8907), .O(n8908) );
  NAND_GATE U9672 ( .I1(n8909), .I2(n8908), .O(n8910) );
  NAND3_GATE U9673 ( .I1(n8912), .I2(n8911), .I3(n8910), .O(n9200) );
  NAND_GATE U9674 ( .I1(B[13]), .I2(A[21]), .O(n9764) );
  NAND_GATE U9675 ( .I1(n8919), .I2(n8918), .O(n8925) );
  INV_GATE U9676 ( .I1(n8920), .O(n8921) );
  NAND_GATE U9677 ( .I1(n8922), .I2(n8921), .O(n8924) );
  NAND_GATE U9678 ( .I1(n8925), .I2(n8924), .O(n8923) );
  NAND_GATE U9679 ( .I1(n8929), .I2(n8923), .O(n8927) );
  NAND3_GATE U9680 ( .I1(n8925), .I2(n8924), .I3(n815), .O(n8926) );
  NAND3_GATE U9681 ( .I1(n8928), .I2(n8927), .I3(n8926), .O(n8935) );
  OR_GATE U9682 ( .I1(n8930), .I2(n8929), .O(n8934) );
  OR_GATE U9683 ( .I1(n8932), .I2(n8931), .O(n8933) );
  NAND3_GATE U9684 ( .I1(n8935), .I2(n8934), .I3(n8933), .O(n9232) );
  NAND_GATE U9685 ( .I1(B[13]), .I2(A[19]), .O(n9244) );
  INV_GATE U9686 ( .I1(n9244), .O(n9176) );
  NAND_GATE U9687 ( .I1(n8939), .I2(n931), .O(n8936) );
  NAND3_GATE U9688 ( .I1(n8938), .I2(n8937), .I3(n8936), .O(n8945) );
  OR_GATE U9689 ( .I1(n8940), .I2(n8939), .O(n8944) );
  OR_GATE U9690 ( .I1(n8942), .I2(n8941), .O(n8943) );
  NAND3_GATE U9691 ( .I1(n8945), .I2(n8944), .I3(n8943), .O(n9484) );
  NAND_GATE U9692 ( .I1(B[13]), .I2(A[18]), .O(n9498) );
  INV_GATE U9693 ( .I1(n9498), .O(n9485) );
  NAND_GATE U9694 ( .I1(n9494), .I2(n9485), .O(n9482) );
  NAND_GATE U9695 ( .I1(B[13]), .I2(A[17]), .O(n9265) );
  INV_GATE U9696 ( .I1(n9265), .O(n9164) );
  NAND_GATE U9697 ( .I1(n8952), .I2(n8585), .O(n8948) );
  NAND_GATE U9698 ( .I1(n8951), .I2(n8948), .O(n8949) );
  AND_GATE U9699 ( .I1(n8950), .I2(n8949), .O(n8956) );
  INV_GATE U9700 ( .I1(n8951), .O(n8954) );
  NAND3_GATE U9701 ( .I1(n8952), .I2(n8954), .I3(n8585), .O(n8957) );
  NAND_GATE U9702 ( .I1(n8956), .I2(n8957), .O(n8955) );
  NAND3_GATE U9703 ( .I1(n8959), .I2(n8955), .I3(n8958), .O(n9271) );
  NAND_GATE U9704 ( .I1(B[13]), .I2(A[16]), .O(n9817) );
  NAND3_GATE U9705 ( .I1(n8957), .I2(n9817), .I3(n8956), .O(n9156) );
  NAND_GATE U9706 ( .I1(n8959), .I2(n8958), .O(n8960) );
  NAND_GATE U9707 ( .I1(n9817), .I2(n8960), .O(n9155) );
  NAND_GATE U9708 ( .I1(B[13]), .I2(A[15]), .O(n9277) );
  INV_GATE U9709 ( .I1(n9277), .O(n9153) );
  NAND_GATE U9710 ( .I1(B[13]), .I2(A[14]), .O(n9834) );
  INV_GATE U9711 ( .I1(n9834), .O(n9468) );
  NAND_GATE U9712 ( .I1(B[13]), .I2(A[13]), .O(n9295) );
  INV_GATE U9713 ( .I1(n9295), .O(n9124) );
  OR_GATE U9714 ( .I1(n8961), .I2(n8966), .O(n8964) );
  OR_GATE U9715 ( .I1(n8965), .I2(n8962), .O(n8963) );
  AND_GATE U9716 ( .I1(n8964), .I2(n8963), .O(n8971) );
  NAND_GATE U9717 ( .I1(n1306), .I2(n8965), .O(n8968) );
  NAND3_GATE U9718 ( .I1(n8969), .I2(n8968), .I3(n8967), .O(n8970) );
  NAND_GATE U9719 ( .I1(n8971), .I2(n8970), .O(n9299) );
  NAND_GATE U9720 ( .I1(B[13]), .I2(A[12]), .O(n9459) );
  INV_GATE U9721 ( .I1(n9459), .O(n9301) );
  NAND_GATE U9722 ( .I1(B[13]), .I2(A[11]), .O(n9309) );
  INV_GATE U9723 ( .I1(n9309), .O(n9107) );
  INV_GATE U9724 ( .I1(n8972), .O(n8973) );
  NAND_GATE U9725 ( .I1(n8973), .I2(n8975), .O(n8983) );
  NAND_GATE U9726 ( .I1(n8974), .I2(n8976), .O(n8981) );
  NAND_GATE U9727 ( .I1(n746), .I2(n8975), .O(n8977) );
  NAND_GATE U9728 ( .I1(n8977), .I2(n8976), .O(n8978) );
  NAND_GATE U9729 ( .I1(n8979), .I2(n8978), .O(n8980) );
  NAND_GATE U9730 ( .I1(n8981), .I2(n8980), .O(n8982) );
  NAND_GATE U9731 ( .I1(n8983), .I2(n8982), .O(n9308) );
  NAND_GATE U9732 ( .I1(n9107), .I2(n9308), .O(n9312) );
  OR_GATE U9733 ( .I1(n8984), .I2(n8989), .O(n8987) );
  OR_GATE U9734 ( .I1(n8988), .I2(n8985), .O(n8986) );
  NAND_GATE U9735 ( .I1(n942), .I2(n8988), .O(n8992) );
  NAND3_GATE U9736 ( .I1(n8992), .I2(n8991), .I3(n8990), .O(n8993) );
  INV_GATE U9737 ( .I1(n9445), .O(n9448) );
  NAND_GATE U9738 ( .I1(B[13]), .I2(A[10]), .O(n9450) );
  INV_GATE U9739 ( .I1(n9450), .O(n9446) );
  NAND_GATE U9740 ( .I1(n9448), .I2(n9446), .O(n9442) );
  NAND_GATE U9741 ( .I1(B[13]), .I2(A[9]), .O(n9323) );
  INV_GATE U9742 ( .I1(n9323), .O(n9103) );
  OR_GATE U9743 ( .I1(n8998), .I2(n8995), .O(n8996) );
  AND_GATE U9744 ( .I1(n8997), .I2(n8996), .O(n9004) );
  NAND_GATE U9745 ( .I1(n1299), .I2(n8998), .O(n9002) );
  NAND3_GATE U9746 ( .I1(n9002), .I2(n9001), .I3(n9000), .O(n9003) );
  NAND_GATE U9747 ( .I1(B[13]), .I2(A[8]), .O(n9433) );
  INV_GATE U9748 ( .I1(n9433), .O(n9428) );
  NAND_GATE U9749 ( .I1(n769), .I2(n9428), .O(n9425) );
  NAND_GATE U9750 ( .I1(B[13]), .I2(A[7]), .O(n9334) );
  INV_GATE U9751 ( .I1(n9334), .O(n9087) );
  OR_GATE U9752 ( .I1(n9005), .I2(n9010), .O(n9008) );
  OR_GATE U9753 ( .I1(n9009), .I2(n9006), .O(n9007) );
  AND_GATE U9754 ( .I1(n9008), .I2(n9007), .O(n9015) );
  NAND_GATE U9755 ( .I1(n1072), .I2(n9009), .O(n9013) );
  NAND3_GATE U9756 ( .I1(n9013), .I2(n9012), .I3(n9011), .O(n9014) );
  NAND_GATE U9757 ( .I1(n9015), .I2(n9014), .O(n9409) );
  INV_GATE U9758 ( .I1(n9409), .O(n9412) );
  NAND_GATE U9759 ( .I1(B[13]), .I2(A[6]), .O(n9416) );
  INV_GATE U9760 ( .I1(n9416), .O(n9410) );
  NAND_GATE U9761 ( .I1(n9412), .I2(n9410), .O(n9406) );
  NAND_GATE U9762 ( .I1(B[13]), .I2(A[5]), .O(n9345) );
  INV_GATE U9763 ( .I1(n9345), .O(n9068) );
  OR_GATE U9764 ( .I1(n9016), .I2(n9021), .O(n9019) );
  OR_GATE U9765 ( .I1(n9020), .I2(n9017), .O(n9018) );
  AND_GATE U9766 ( .I1(n9019), .I2(n9018), .O(n9026) );
  NAND_GATE U9767 ( .I1(n1167), .I2(n9020), .O(n9024) );
  NAND3_GATE U9768 ( .I1(n9024), .I2(n9023), .I3(n9022), .O(n9025) );
  NAND_GATE U9769 ( .I1(n9026), .I2(n9025), .O(n9353) );
  INV_GATE U9770 ( .I1(n9353), .O(n9356) );
  NAND_GATE U9771 ( .I1(B[13]), .I2(A[4]), .O(n9360) );
  INV_GATE U9772 ( .I1(n9360), .O(n9354) );
  NAND_GATE U9773 ( .I1(n9356), .I2(n9354), .O(n9350) );
  OR_GATE U9774 ( .I1(n9028), .I2(n9027), .O(n9040) );
  NAND_GATE U9775 ( .I1(n9029), .I2(n9028), .O(n9034) );
  NAND_GATE U9776 ( .I1(n9030), .I2(n9034), .O(n9038) );
  NAND_GATE U9777 ( .I1(n9032), .I2(n9031), .O(n9033) );
  NAND_GATE U9778 ( .I1(n9034), .I2(n9033), .O(n9035) );
  NAND_GATE U9779 ( .I1(n9036), .I2(n9035), .O(n9037) );
  NAND_GATE U9780 ( .I1(n9038), .I2(n9037), .O(n9039) );
  NAND_GATE U9781 ( .I1(n9040), .I2(n9039), .O(n9393) );
  NAND3_GATE U9782 ( .I1(B[13]), .I2(B[14]), .I3(n1196), .O(n9367) );
  INV_GATE U9783 ( .I1(n9367), .O(n9370) );
  NAND_GATE U9784 ( .I1(n1378), .I2(A[0]), .O(n9041) );
  NAND_GATE U9785 ( .I1(n14781), .I2(n9041), .O(n9042) );
  NAND_GATE U9786 ( .I1(n1379), .I2(n9042), .O(n9046) );
  NAND_GATE U9787 ( .I1(n1380), .I2(A[1]), .O(n9043) );
  NAND_GATE U9788 ( .I1(n14784), .I2(n9043), .O(n9044) );
  NAND_GATE U9789 ( .I1(B[14]), .I2(n9044), .O(n9045) );
  NAND_GATE U9790 ( .I1(n9046), .I2(n9045), .O(n9369) );
  INV_GATE U9791 ( .I1(n9369), .O(n9366) );
  NAND_GATE U9792 ( .I1(B[13]), .I2(A[2]), .O(n9374) );
  NAND_GATE U9793 ( .I1(n9366), .I2(n9374), .O(n9047) );
  NAND_GATE U9794 ( .I1(n9370), .I2(n9047), .O(n9048) );
  INV_GATE U9795 ( .I1(n9374), .O(n9368) );
  NAND_GATE U9796 ( .I1(n9369), .I2(n9368), .O(n9365) );
  NAND_GATE U9797 ( .I1(n9048), .I2(n9365), .O(n9394) );
  NAND_GATE U9798 ( .I1(n9393), .I2(n9394), .O(n9050) );
  NAND_GATE U9799 ( .I1(B[13]), .I2(A[3]), .O(n9395) );
  INV_GATE U9800 ( .I1(n9395), .O(n9049) );
  NAND_GATE U9801 ( .I1(n9394), .I2(n9049), .O(n9390) );
  NAND_GATE U9802 ( .I1(n9393), .I2(n9049), .O(n9389) );
  NAND3_GATE U9803 ( .I1(n9050), .I2(n9390), .I3(n9389), .O(n9355) );
  NAND_GATE U9804 ( .I1(n9353), .I2(n9360), .O(n9051) );
  NAND_GATE U9805 ( .I1(n9355), .I2(n9051), .O(n9052) );
  NAND_GATE U9806 ( .I1(n9350), .I2(n9052), .O(n9344) );
  NAND_GATE U9807 ( .I1(n9068), .I2(n9344), .O(n9340) );
  INV_GATE U9808 ( .I1(n9053), .O(n9054) );
  NAND_GATE U9809 ( .I1(n9054), .I2(n9058), .O(n9067) );
  INV_GATE U9810 ( .I1(n9058), .O(n9055) );
  NAND_GATE U9811 ( .I1(n9056), .I2(n9055), .O(n9061) );
  NAND_GATE U9812 ( .I1(n9057), .I2(n9061), .O(n9065) );
  NAND_GATE U9813 ( .I1(n9059), .I2(n9058), .O(n9060) );
  NAND_GATE U9814 ( .I1(n9061), .I2(n9060), .O(n9062) );
  NAND_GATE U9815 ( .I1(n9063), .I2(n9062), .O(n9064) );
  NAND_GATE U9816 ( .I1(n9065), .I2(n9064), .O(n9066) );
  NAND_GATE U9817 ( .I1(n9067), .I2(n9066), .O(n9343) );
  NAND_GATE U9818 ( .I1(n9344), .I2(n9343), .O(n9069) );
  NAND_GATE U9819 ( .I1(n9068), .I2(n9343), .O(n9339) );
  NAND3_GATE U9820 ( .I1(n9340), .I2(n9069), .I3(n9339), .O(n9411) );
  NAND_GATE U9821 ( .I1(n9409), .I2(n9416), .O(n9070) );
  NAND_GATE U9822 ( .I1(n9411), .I2(n9070), .O(n9071) );
  NAND_GATE U9823 ( .I1(n9406), .I2(n9071), .O(n9333) );
  NAND_GATE U9824 ( .I1(n9087), .I2(n9333), .O(n9329) );
  INV_GATE U9825 ( .I1(n9072), .O(n9073) );
  NAND_GATE U9826 ( .I1(n9073), .I2(n9077), .O(n9086) );
  INV_GATE U9827 ( .I1(n9077), .O(n9074) );
  NAND_GATE U9828 ( .I1(n9075), .I2(n9074), .O(n9080) );
  NAND_GATE U9829 ( .I1(n9076), .I2(n9080), .O(n9084) );
  NAND_GATE U9830 ( .I1(n9078), .I2(n9077), .O(n9079) );
  NAND_GATE U9831 ( .I1(n9080), .I2(n9079), .O(n9081) );
  NAND_GATE U9832 ( .I1(n9082), .I2(n9081), .O(n9083) );
  NAND_GATE U9833 ( .I1(n9084), .I2(n9083), .O(n9085) );
  NAND_GATE U9834 ( .I1(n9086), .I2(n9085), .O(n9332) );
  NAND_GATE U9835 ( .I1(n9333), .I2(n9332), .O(n9088) );
  NAND_GATE U9836 ( .I1(n9087), .I2(n9332), .O(n9328) );
  NAND3_GATE U9837 ( .I1(n9329), .I2(n9088), .I3(n9328), .O(n9429) );
  NAND_GATE U9838 ( .I1(n9427), .I2(n9433), .O(n9089) );
  NAND_GATE U9839 ( .I1(n9429), .I2(n9089), .O(n9090) );
  NAND_GATE U9840 ( .I1(n9425), .I2(n9090), .O(n9322) );
  NAND_GATE U9841 ( .I1(n9103), .I2(n9322), .O(n9318) );
  INV_GATE U9842 ( .I1(n9091), .O(n9092) );
  NAND_GATE U9843 ( .I1(n9092), .I2(n9095), .O(n9102) );
  NAND_GATE U9844 ( .I1(n9093), .I2(n768), .O(n9097) );
  NAND_GATE U9845 ( .I1(n9094), .I2(n9097), .O(n9100) );
  NAND_GATE U9846 ( .I1(n9100), .I2(n9099), .O(n9101) );
  NAND_GATE U9847 ( .I1(n9102), .I2(n9101), .O(n9321) );
  NAND_GATE U9848 ( .I1(n9322), .I2(n9321), .O(n9104) );
  NAND_GATE U9849 ( .I1(n9103), .I2(n9321), .O(n9317) );
  NAND3_GATE U9850 ( .I1(n9318), .I2(n9104), .I3(n9317), .O(n9447) );
  NAND_GATE U9851 ( .I1(n9445), .I2(n9450), .O(n9105) );
  NAND_GATE U9852 ( .I1(n9447), .I2(n9105), .O(n9106) );
  NAND_GATE U9853 ( .I1(n9442), .I2(n9106), .O(n9313) );
  NAND_GATE U9854 ( .I1(n9308), .I2(n9313), .O(n9108) );
  NAND_GATE U9855 ( .I1(n9107), .I2(n9313), .O(n9307) );
  NAND_GATE U9856 ( .I1(n9299), .I2(n9459), .O(n9109) );
  NAND_GATE U9857 ( .I1(n9303), .I2(n9109), .O(n9110) );
  NAND_GATE U9858 ( .I1(n9302), .I2(n9110), .O(n9292) );
  NAND_GATE U9859 ( .I1(n9124), .I2(n9292), .O(n9286) );
  NAND_GATE U9860 ( .I1(n9113), .I2(n168), .O(n9111) );
  NAND_GATE U9861 ( .I1(n9112), .I2(n9111), .O(n9118) );
  NAND_GATE U9862 ( .I1(n1204), .I2(n9120), .O(n9114) );
  NAND_GATE U9863 ( .I1(n9114), .I2(n9111), .O(n9115) );
  NAND_GATE U9864 ( .I1(n9116), .I2(n9115), .O(n9117) );
  NAND_GATE U9865 ( .I1(n9118), .I2(n9117), .O(n9123) );
  INV_GATE U9866 ( .I1(n9119), .O(n9121) );
  NAND_GATE U9867 ( .I1(n9121), .I2(n9120), .O(n9122) );
  NAND_GATE U9868 ( .I1(n9123), .I2(n9122), .O(n9290) );
  NAND_GATE U9869 ( .I1(n9292), .I2(n9290), .O(n9125) );
  NAND_GATE U9870 ( .I1(n9124), .I2(n9290), .O(n9285) );
  OR_GATE U9871 ( .I1(n9126), .I2(n9128), .O(n9136) );
  INV_GATE U9872 ( .I1(n9133), .O(n9127) );
  NAND_GATE U9873 ( .I1(n9128), .I2(n9127), .O(n9130) );
  NAND_GATE U9874 ( .I1(n1341), .I2(n9133), .O(n9129) );
  NAND3_GATE U9875 ( .I1(n9131), .I2(n9130), .I3(n9129), .O(n9135) );
  OR_GATE U9876 ( .I1(n9133), .I2(n9132), .O(n9134) );
  NAND3_GATE U9877 ( .I1(n9136), .I2(n9135), .I3(n9134), .O(n9470) );
  INV_GATE U9878 ( .I1(n9470), .O(n9469) );
  NAND_GATE U9879 ( .I1(n9834), .I2(n632), .O(n9137) );
  NAND_GATE U9880 ( .I1(n9469), .I2(n9137), .O(n9138) );
  NAND_GATE U9881 ( .I1(n9467), .I2(n9138), .O(n9278) );
  NAND_GATE U9882 ( .I1(n9153), .I2(n9278), .O(n9280) );
  NAND_GATE U9883 ( .I1(n9139), .I2(n9149), .O(n9140) );
  NAND_GATE U9884 ( .I1(n9144), .I2(n9140), .O(n9141) );
  NAND_GATE U9885 ( .I1(n9142), .I2(n9141), .O(n9147) );
  NAND_GATE U9886 ( .I1(n9145), .I2(n9144), .O(n9146) );
  NAND_GATE U9887 ( .I1(n9147), .I2(n9146), .O(n9152) );
  INV_GATE U9888 ( .I1(n9148), .O(n9150) );
  NAND_GATE U9889 ( .I1(n9150), .I2(n9149), .O(n9151) );
  NAND_GATE U9890 ( .I1(n9152), .I2(n9151), .O(n9281) );
  NAND_GATE U9891 ( .I1(n9278), .I2(n9281), .O(n9154) );
  NAND_GATE U9892 ( .I1(n9153), .I2(n9281), .O(n9279) );
  NAND3_GATE U9893 ( .I1(n9280), .I2(n9154), .I3(n9279), .O(n9272) );
  NAND3_GATE U9894 ( .I1(n9156), .I2(n9155), .I3(n9272), .O(n9157) );
  NAND_GATE U9895 ( .I1(n9269), .I2(n9157), .O(n9261) );
  NAND_GATE U9896 ( .I1(n9164), .I2(n9261), .O(n9252) );
  NAND3_GATE U9897 ( .I1(n9160), .I2(n9161), .I3(n9158), .O(n9255) );
  NAND_GATE U9898 ( .I1(n1301), .I2(n9255), .O(n9260) );
  NAND_GATE U9899 ( .I1(n9159), .I2(n1200), .O(n9163) );
  NAND_GATE U9900 ( .I1(n9161), .I2(n9160), .O(n9162) );
  NAND_GATE U9901 ( .I1(n9163), .I2(n9162), .O(n9257) );
  NAND_GATE U9902 ( .I1(n9258), .I2(n9257), .O(n9256) );
  NAND3_GATE U9903 ( .I1(n9261), .I2(n9260), .I3(n9256), .O(n9166) );
  NAND_GATE U9904 ( .I1(n9256), .I2(n950), .O(n9165) );
  NAND3_GATE U9905 ( .I1(n9252), .I2(n9166), .I3(n9165), .O(n9493) );
  NAND_GATE U9906 ( .I1(n9484), .I2(n9498), .O(n9167) );
  NAND_GATE U9907 ( .I1(n9493), .I2(n9167), .O(n9168) );
  NAND_GATE U9908 ( .I1(n9482), .I2(n9168), .O(n9245) );
  NAND_GATE U9909 ( .I1(n9176), .I2(n9245), .O(n9247) );
  NAND3_GATE U9910 ( .I1(n9171), .I2(n9172), .I3(n9169), .O(n9238) );
  NAND_GATE U9911 ( .I1(n9169), .I2(n9174), .O(n9236) );
  NAND_GATE U9912 ( .I1(n9170), .I2(n822), .O(n9174) );
  NAND_GATE U9913 ( .I1(n9172), .I2(n9171), .O(n9173) );
  NAND_GATE U9914 ( .I1(n9174), .I2(n9173), .O(n9234) );
  NAND_GATE U9915 ( .I1(n9236), .I2(n9240), .O(n9175) );
  NAND_GATE U9916 ( .I1(n9238), .I2(n9175), .O(n9248) );
  NAND_GATE U9917 ( .I1(n9176), .I2(n9248), .O(n9246) );
  NAND_GATE U9918 ( .I1(n9245), .I2(n9248), .O(n9177) );
  NAND3_GATE U9919 ( .I1(n9247), .I2(n9246), .I3(n9177), .O(n9506) );
  NAND_GATE U9920 ( .I1(B[13]), .I2(A[20]), .O(n9779) );
  NAND_GATE U9921 ( .I1(n9179), .I2(n9178), .O(n9182) );
  INV_GATE U9922 ( .I1(n9185), .O(n9190) );
  NAND_GATE U9923 ( .I1(n186), .I2(n9181), .O(n9183) );
  NAND3_GATE U9924 ( .I1(n9182), .I2(n9190), .I3(n9183), .O(n9188) );
  NAND_GATE U9925 ( .I1(n9183), .I2(n9182), .O(n9184) );
  NAND_GATE U9926 ( .I1(n9185), .I2(n9184), .O(n9187) );
  NAND3_GATE U9927 ( .I1(n9188), .I2(n9187), .I3(n9186), .O(n9195) );
  NAND3_GATE U9928 ( .I1(n9190), .I2(n9189), .I3(n9192), .O(n9194) );
  OR_GATE U9929 ( .I1(n9192), .I2(n9191), .O(n9193) );
  NAND3_GATE U9930 ( .I1(n9195), .I2(n9194), .I3(n9193), .O(n9507) );
  NAND_GATE U9931 ( .I1(n9779), .I2(n9507), .O(n9196) );
  NAND_GATE U9932 ( .I1(n9506), .I2(n9196), .O(n9198) );
  INV_GATE U9933 ( .I1(n9779), .O(n9503) );
  NAND_GATE U9934 ( .I1(n9503), .I2(n9505), .O(n9197) );
  NAND_GATE U9935 ( .I1(n9198), .I2(n9197), .O(n9233) );
  NAND_GATE U9936 ( .I1(n9764), .I2(n9232), .O(n9199) );
  NAND4_GATE U9937 ( .I1(n9201), .I2(n9200), .I3(n9202), .I4(n9229), .O(n9204)
         );
  NAND_GATE U9938 ( .I1(B[13]), .I2(A[22]), .O(n9226) );
  INV_GATE U9939 ( .I1(n9226), .O(n9749) );
  NAND_GATE U9940 ( .I1(n9749), .I2(n9229), .O(n9203) );
  NAND3_GATE U9941 ( .I1(n9202), .I2(n9201), .I3(n9200), .O(n9227) );
  NAND_GATE U9942 ( .I1(n9749), .I2(n210), .O(n9228) );
  NAND3_GATE U9943 ( .I1(n9204), .I2(n9203), .I3(n9228), .O(n9529) );
  NAND_GATE U9944 ( .I1(n9522), .I2(n9524), .O(n9205) );
  NAND_GATE U9945 ( .I1(n9529), .I2(n9205), .O(n9206) );
  NAND_GATE U9946 ( .I1(n9720), .I2(n9538), .O(n9207) );
  NAND_GATE U9947 ( .I1(n9536), .I2(n9207), .O(n9208) );
  NAND_GATE U9948 ( .I1(n9209), .I2(n9208), .O(n9548) );
  NAND_GATE U9949 ( .I1(n9552), .I2(n9550), .O(n9210) );
  NAND_GATE U9950 ( .I1(n9548), .I2(n9210), .O(n9211) );
  NAND_GATE U9951 ( .I1(n9544), .I2(n9211), .O(n9563) );
  NAND_GATE U9952 ( .I1(n9564), .I2(n9567), .O(n9212) );
  NAND_GATE U9953 ( .I1(n9563), .I2(n9212), .O(n9213) );
  NAND_GATE U9954 ( .I1(n9560), .I2(n9213), .O(n9575) );
  NAND_GATE U9955 ( .I1(n9578), .I2(n9580), .O(n9214) );
  NAND_GATE U9956 ( .I1(n9575), .I2(n9214), .O(n9215) );
  NAND_GATE U9957 ( .I1(n9572), .I2(n9215), .O(n9590) );
  NAND_GATE U9958 ( .I1(n9591), .I2(n9594), .O(n9216) );
  NAND_GATE U9959 ( .I1(n9590), .I2(n9216), .O(n9217) );
  NAND_GATE U9960 ( .I1(n9586), .I2(n9217), .O(n9605) );
  NAND_GATE U9961 ( .I1(n9607), .I2(n9610), .O(n9218) );
  NAND_GATE U9962 ( .I1(n9605), .I2(n9218), .O(n9219) );
  NAND_GATE U9963 ( .I1(n9601), .I2(n9219), .O(n9621) );
  NAND_GATE U9964 ( .I1(n9619), .I2(n9626), .O(n9220) );
  NAND_GATE U9965 ( .I1(n9621), .I2(n9220), .O(n9221) );
  NAND_GATE U9966 ( .I1(n9617), .I2(n9221), .O(n9637) );
  NAND_GATE U9967 ( .I1(n9635), .I2(n9642), .O(n9222) );
  NAND_GATE U9968 ( .I1(n9637), .I2(n9222), .O(n9223) );
  NAND_GATE U9969 ( .I1(n9224), .I2(n284), .O(n9225) );
  AND_GATE U9970 ( .I1(n15331), .I2(n9225), .O(\A1[43] ) );
  NAND_GATE U9971 ( .I1(B[12]), .I2(A[31]), .O(n9657) );
  INV_GATE U9972 ( .I1(n9657), .O(n9631) );
  NAND_GATE U9973 ( .I1(B[12]), .I2(A[30]), .O(n9668) );
  INV_GATE U9974 ( .I1(n9668), .O(n9615) );
  NAND_GATE U9975 ( .I1(B[12]), .I2(A[29]), .O(n9673) );
  INV_GATE U9976 ( .I1(n9673), .O(n9599) );
  NAND_GATE U9977 ( .I1(B[12]), .I2(A[28]), .O(n9683) );
  INV_GATE U9978 ( .I1(n9683), .O(n9584) );
  NAND_GATE U9979 ( .I1(B[12]), .I2(A[27]), .O(n9702) );
  INV_GATE U9980 ( .I1(n9702), .O(n9570) );
  NAND_GATE U9981 ( .I1(B[12]), .I2(A[26]), .O(n9707) );
  INV_GATE U9982 ( .I1(n9707), .O(n9710) );
  NAND_GATE U9983 ( .I1(B[12]), .I2(A[25]), .O(n9730) );
  INV_GATE U9984 ( .I1(n9730), .O(n9723) );
  NAND_GATE U9985 ( .I1(B[12]), .I2(A[24]), .O(n9745) );
  INV_GATE U9986 ( .I1(n9745), .O(n9736) );
  NAND3_GATE U9987 ( .I1(n9227), .I2(n14), .I3(n9226), .O(n9750) );
  NAND3_GATE U9988 ( .I1(n210), .I2(n9229), .I3(n9226), .O(n9752) );
  NAND_GATE U9989 ( .I1(n9227), .I2(n14), .O(n9748) );
  NAND3_GATE U9990 ( .I1(n9749), .I2(n9748), .I3(n9755), .O(n9759) );
  NAND_GATE U9991 ( .I1(B[12]), .I2(A[22]), .O(n9768) );
  INV_GATE U9992 ( .I1(n9768), .O(n9513) );
  NAND_GATE U9993 ( .I1(n9232), .I2(n921), .O(n9231) );
  NAND_GATE U9994 ( .I1(n9231), .I2(n9230), .O(n9763) );
  NAND_GATE U9995 ( .I1(n1212), .I2(n9233), .O(n9515) );
  NAND_GATE U9996 ( .I1(n876), .I2(n9515), .O(n9766) );
  NAND3_GATE U9997 ( .I1(n9513), .I2(n9765), .I3(n9766), .O(n9773) );
  NAND_GATE U9998 ( .I1(B[12]), .I2(A[21]), .O(n9782) );
  INV_GATE U9999 ( .I1(n9782), .O(n9504) );
  NAND_GATE U10000 ( .I1(B[12]), .I2(A[20]), .O(n10078) );
  INV_GATE U10001 ( .I1(n10078), .O(n10066) );
  NAND_GATE U10002 ( .I1(n9235), .I2(n9234), .O(n9240) );
  INV_GATE U10003 ( .I1(n9236), .O(n9237) );
  NAND_GATE U10004 ( .I1(n9238), .I2(n9237), .O(n9241) );
  NAND_GATE U10005 ( .I1(n9240), .I2(n9241), .O(n9239) );
  NAND_GATE U10006 ( .I1(n9245), .I2(n9239), .O(n9243) );
  NAND3_GATE U10007 ( .I1(n9241), .I2(n246), .I3(n9240), .O(n9242) );
  NAND3_GATE U10008 ( .I1(n9244), .I2(n9243), .I3(n9242), .O(n9251) );
  OR_GATE U10009 ( .I1(n9248), .I2(n9247), .O(n9249) );
  NAND3_GATE U10010 ( .I1(n9251), .I2(n9250), .I3(n9249), .O(n10069) );
  NAND_GATE U10011 ( .I1(n10066), .I2(n10067), .O(n10071) );
  NAND_GATE U10012 ( .I1(B[12]), .I2(A[19]), .O(n9797) );
  INV_GATE U10013 ( .I1(n9797), .O(n9492) );
  INV_GATE U10014 ( .I1(n9252), .O(n9253) );
  NAND3_GATE U10015 ( .I1(n9255), .I2(n9254), .I3(n9253), .O(n9268) );
  NAND3_GATE U10016 ( .I1(n671), .I2(n950), .I3(n9256), .O(n9267) );
  NAND_GATE U10017 ( .I1(n9260), .I2(n9259), .O(n9262) );
  NAND_GATE U10018 ( .I1(n9261), .I2(n9262), .O(n9264) );
  NAND3_GATE U10019 ( .I1(n9265), .I2(n9264), .I3(n9263), .O(n9266) );
  NAND3_GATE U10020 ( .I1(n9268), .I2(n9267), .I3(n9266), .O(n10055) );
  NAND_GATE U10021 ( .I1(B[12]), .I2(A[18]), .O(n10052) );
  INV_GATE U10022 ( .I1(n10052), .O(n10057) );
  NAND_GATE U10023 ( .I1(n672), .I2(n10057), .O(n10051) );
  NAND_GATE U10024 ( .I1(B[12]), .I2(A[17]), .O(n9811) );
  INV_GATE U10025 ( .I1(n9811), .O(n9478) );
  INV_GATE U10026 ( .I1(n9272), .O(n9270) );
  NAND_GATE U10027 ( .I1(n9271), .I2(n9270), .O(n9274) );
  NAND_GATE U10028 ( .I1(n9274), .I2(n9273), .O(n9816) );
  NAND_GATE U10029 ( .I1(n9817), .I2(n9816), .O(n9808) );
  NAND3_GATE U10030 ( .I1(n9478), .I2(n9809), .I3(n9808), .O(n9815) );
  NAND_GATE U10031 ( .I1(n967), .I2(n9281), .O(n9276) );
  NAND3_GATE U10032 ( .I1(n9277), .I2(n9276), .I3(n9275), .O(n9284) );
  OR_GATE U10033 ( .I1(n9279), .I2(n9278), .O(n9283) );
  OR_GATE U10034 ( .I1(n9281), .I2(n9280), .O(n9282) );
  NAND3_GATE U10035 ( .I1(n9284), .I2(n9283), .I3(n9282), .O(n10040) );
  NAND_GATE U10036 ( .I1(B[12]), .I2(A[16]), .O(n10039) );
  NAND_GATE U10037 ( .I1(B[12]), .I2(A[14]), .O(n10025) );
  INV_GATE U10038 ( .I1(n10025), .O(n10020) );
  OR_GATE U10039 ( .I1(n9285), .I2(n9292), .O(n9288) );
  OR_GATE U10040 ( .I1(n9290), .I2(n9286), .O(n9287) );
  AND_GATE U10041 ( .I1(n9288), .I2(n9287), .O(n9297) );
  INV_GATE U10042 ( .I1(n9292), .O(n9289) );
  NAND_GATE U10043 ( .I1(n9289), .I2(n9290), .O(n9294) );
  INV_GATE U10044 ( .I1(n9290), .O(n9291) );
  NAND_GATE U10045 ( .I1(n9292), .I2(n9291), .O(n9293) );
  NAND3_GATE U10046 ( .I1(n9295), .I2(n9294), .I3(n9293), .O(n9296) );
  NAND_GATE U10047 ( .I1(n9297), .I2(n9296), .O(n10022) );
  NAND_GATE U10048 ( .I1(n10020), .I2(n1203), .O(n10028) );
  NAND_GATE U10049 ( .I1(n9300), .I2(n9298), .O(n9458) );
  NAND_GATE U10050 ( .I1(n9459), .I2(n9458), .O(n9306) );
  NAND_GATE U10051 ( .I1(n9299), .I2(n844), .O(n9300) );
  NAND_GATE U10052 ( .I1(n9301), .I2(n9300), .O(n9460) );
  INV_GATE U10053 ( .I1(n9460), .O(n9304) );
  NAND_GATE U10054 ( .I1(n9304), .I2(n9462), .O(n9305) );
  NAND4_GATE U10055 ( .I1(n9306), .I2(n9305), .I3(A[13]), .I4(B[12]), .O(n9848) );
  NAND_GATE U10056 ( .I1(B[12]), .I2(A[12]), .O(n9860) );
  INV_GATE U10057 ( .I1(n9860), .O(n9855) );
  OR_GATE U10058 ( .I1(n9307), .I2(n9308), .O(n9316) );
  NAND_GATE U10059 ( .I1(n9308), .I2(n940), .O(n9311) );
  NAND3_GATE U10060 ( .I1(n9311), .I2(n9310), .I3(n9309), .O(n9315) );
  OR_GATE U10061 ( .I1(n9313), .I2(n9312), .O(n9314) );
  NAND3_GATE U10062 ( .I1(n9316), .I2(n9315), .I3(n9314), .O(n9853) );
  NAND_GATE U10063 ( .I1(B[12]), .I2(A[11]), .O(n10010) );
  INV_GATE U10064 ( .I1(n10010), .O(n9455) );
  OR_GATE U10065 ( .I1(n9321), .I2(n9318), .O(n9319) );
  AND_GATE U10066 ( .I1(n9320), .I2(n9319), .O(n9327) );
  NAND_GATE U10067 ( .I1(n971), .I2(n9321), .O(n9325) );
  NAND3_GATE U10068 ( .I1(n9325), .I2(n9324), .I3(n9323), .O(n9326) );
  NAND_GATE U10069 ( .I1(n9327), .I2(n9326), .O(n9990) );
  INV_GATE U10070 ( .I1(n9990), .O(n9993) );
  NAND_GATE U10071 ( .I1(B[12]), .I2(A[10]), .O(n9997) );
  INV_GATE U10072 ( .I1(n9997), .O(n9991) );
  NAND_GATE U10073 ( .I1(n9993), .I2(n9991), .O(n9987) );
  NAND_GATE U10074 ( .I1(B[12]), .I2(A[9]), .O(n9869) );
  INV_GATE U10075 ( .I1(n9869), .O(n9438) );
  OR_GATE U10076 ( .I1(n9332), .I2(n9329), .O(n9330) );
  AND_GATE U10077 ( .I1(n9331), .I2(n9330), .O(n9338) );
  NAND_GATE U10078 ( .I1(n944), .I2(n9332), .O(n9336) );
  NAND3_GATE U10079 ( .I1(n9336), .I2(n9335), .I3(n9334), .O(n9337) );
  NAND_GATE U10080 ( .I1(B[12]), .I2(A[8]), .O(n9978) );
  INV_GATE U10081 ( .I1(n9978), .O(n9974) );
  NAND_GATE U10082 ( .I1(n633), .I2(n9974), .O(n9971) );
  NAND_GATE U10083 ( .I1(B[12]), .I2(A[7]), .O(n9880) );
  INV_GATE U10084 ( .I1(n9880), .O(n9421) );
  OR_GATE U10085 ( .I1(n9339), .I2(n9344), .O(n9342) );
  OR_GATE U10086 ( .I1(n9343), .I2(n9340), .O(n9341) );
  AND_GATE U10087 ( .I1(n9342), .I2(n9341), .O(n9349) );
  NAND_GATE U10088 ( .I1(n1089), .I2(n9343), .O(n9347) );
  NAND3_GATE U10089 ( .I1(n9347), .I2(n9346), .I3(n9345), .O(n9348) );
  NAND_GATE U10090 ( .I1(n9349), .I2(n9348), .O(n9888) );
  INV_GATE U10091 ( .I1(n9888), .O(n9891) );
  NAND_GATE U10092 ( .I1(B[12]), .I2(A[6]), .O(n9895) );
  INV_GATE U10093 ( .I1(n9895), .O(n9889) );
  NAND_GATE U10094 ( .I1(n9891), .I2(n9889), .O(n9885) );
  INV_GATE U10095 ( .I1(n9350), .O(n9351) );
  NAND_GATE U10096 ( .I1(n9351), .I2(n9355), .O(n9364) );
  INV_GATE U10097 ( .I1(n9355), .O(n9352) );
  NAND_GATE U10098 ( .I1(n9353), .I2(n9352), .O(n9358) );
  NAND_GATE U10099 ( .I1(n9354), .I2(n9358), .O(n9362) );
  NAND_GATE U10100 ( .I1(n9356), .I2(n9355), .O(n9357) );
  NAND_GATE U10101 ( .I1(n9358), .I2(n9357), .O(n9359) );
  NAND_GATE U10102 ( .I1(n9360), .I2(n9359), .O(n9361) );
  NAND_GATE U10103 ( .I1(n9362), .I2(n9361), .O(n9363) );
  NAND_GATE U10104 ( .I1(n9364), .I2(n9363), .O(n9958) );
  OR_GATE U10105 ( .I1(n9365), .I2(n9367), .O(n9378) );
  NAND_GATE U10106 ( .I1(n9367), .I2(n9366), .O(n9372) );
  NAND_GATE U10107 ( .I1(n9368), .I2(n9372), .O(n9376) );
  NAND_GATE U10108 ( .I1(n9370), .I2(n9369), .O(n9371) );
  NAND_GATE U10109 ( .I1(n9372), .I2(n9371), .O(n9373) );
  NAND_GATE U10110 ( .I1(n9374), .I2(n9373), .O(n9375) );
  NAND_GATE U10111 ( .I1(n9376), .I2(n9375), .O(n9377) );
  NAND_GATE U10112 ( .I1(n9378), .I2(n9377), .O(n9943) );
  NAND3_GATE U10113 ( .I1(B[12]), .I2(B[13]), .I3(n1196), .O(n9917) );
  INV_GATE U10114 ( .I1(n9917), .O(n9920) );
  NAND_GATE U10115 ( .I1(n1377), .I2(A[0]), .O(n9379) );
  NAND_GATE U10116 ( .I1(n14781), .I2(n9379), .O(n9380) );
  NAND_GATE U10117 ( .I1(B[14]), .I2(n9380), .O(n9384) );
  NAND_GATE U10118 ( .I1(n1378), .I2(A[1]), .O(n9381) );
  NAND_GATE U10119 ( .I1(n14784), .I2(n9381), .O(n9382) );
  NAND_GATE U10120 ( .I1(B[13]), .I2(n9382), .O(n9383) );
  NAND_GATE U10121 ( .I1(n9384), .I2(n9383), .O(n9919) );
  INV_GATE U10122 ( .I1(n9919), .O(n9916) );
  NAND_GATE U10123 ( .I1(B[12]), .I2(A[2]), .O(n9924) );
  NAND_GATE U10124 ( .I1(n9916), .I2(n9924), .O(n9385) );
  NAND_GATE U10125 ( .I1(n9920), .I2(n9385), .O(n9386) );
  INV_GATE U10126 ( .I1(n9924), .O(n9918) );
  NAND_GATE U10127 ( .I1(n9919), .I2(n9918), .O(n9915) );
  NAND_GATE U10128 ( .I1(n9386), .I2(n9915), .O(n9944) );
  NAND_GATE U10129 ( .I1(n9943), .I2(n9944), .O(n9388) );
  NAND_GATE U10130 ( .I1(B[12]), .I2(A[3]), .O(n9945) );
  INV_GATE U10131 ( .I1(n9945), .O(n9387) );
  NAND_GATE U10132 ( .I1(n9944), .I2(n9387), .O(n9940) );
  NAND_GATE U10133 ( .I1(n9943), .I2(n9387), .O(n9939) );
  NAND3_GATE U10134 ( .I1(n9388), .I2(n9940), .I3(n9939), .O(n9906) );
  NAND_GATE U10135 ( .I1(B[12]), .I2(A[4]), .O(n9910) );
  OR_GATE U10136 ( .I1(n9389), .I2(n9394), .O(n9392) );
  OR_GATE U10137 ( .I1(n9390), .I2(n9393), .O(n9391) );
  AND_GATE U10138 ( .I1(n9392), .I2(n9391), .O(n9399) );
  NAND_GATE U10139 ( .I1(n9393), .I2(n1169), .O(n9397) );
  NAND3_GATE U10140 ( .I1(n9397), .I2(n9396), .I3(n9395), .O(n9398) );
  NAND_GATE U10141 ( .I1(n9399), .I2(n9398), .O(n9902) );
  NAND_GATE U10142 ( .I1(n9910), .I2(n9902), .O(n9400) );
  NAND_GATE U10143 ( .I1(n9906), .I2(n9400), .O(n9401) );
  INV_GATE U10144 ( .I1(n9910), .O(n9904) );
  INV_GATE U10145 ( .I1(n9902), .O(n9905) );
  NAND_GATE U10146 ( .I1(n9904), .I2(n9905), .O(n9900) );
  NAND_GATE U10147 ( .I1(n9401), .I2(n9900), .O(n9959) );
  NAND_GATE U10148 ( .I1(n9958), .I2(n9959), .O(n9403) );
  NAND_GATE U10149 ( .I1(B[12]), .I2(A[5]), .O(n9960) );
  INV_GATE U10150 ( .I1(n9960), .O(n9402) );
  NAND_GATE U10151 ( .I1(n9959), .I2(n9402), .O(n9955) );
  NAND_GATE U10152 ( .I1(n9958), .I2(n9402), .O(n9954) );
  NAND3_GATE U10153 ( .I1(n9403), .I2(n9955), .I3(n9954), .O(n9890) );
  NAND_GATE U10154 ( .I1(n9888), .I2(n9895), .O(n9404) );
  NAND_GATE U10155 ( .I1(n9890), .I2(n9404), .O(n9405) );
  NAND_GATE U10156 ( .I1(n9885), .I2(n9405), .O(n9879) );
  NAND_GATE U10157 ( .I1(n9421), .I2(n9879), .O(n9875) );
  INV_GATE U10158 ( .I1(n9406), .O(n9407) );
  NAND_GATE U10159 ( .I1(n9407), .I2(n9411), .O(n9420) );
  INV_GATE U10160 ( .I1(n9411), .O(n9408) );
  NAND_GATE U10161 ( .I1(n9409), .I2(n9408), .O(n9414) );
  NAND_GATE U10162 ( .I1(n9410), .I2(n9414), .O(n9418) );
  NAND_GATE U10163 ( .I1(n9412), .I2(n9411), .O(n9413) );
  NAND_GATE U10164 ( .I1(n9414), .I2(n9413), .O(n9415) );
  NAND_GATE U10165 ( .I1(n9416), .I2(n9415), .O(n9417) );
  NAND_GATE U10166 ( .I1(n9418), .I2(n9417), .O(n9419) );
  NAND_GATE U10167 ( .I1(n9420), .I2(n9419), .O(n9878) );
  NAND_GATE U10168 ( .I1(n9879), .I2(n9878), .O(n9422) );
  NAND_GATE U10169 ( .I1(n9421), .I2(n9878), .O(n9874) );
  NAND3_GATE U10170 ( .I1(n9875), .I2(n9422), .I3(n9874), .O(n9975) );
  NAND_GATE U10171 ( .I1(n9973), .I2(n9978), .O(n9423) );
  NAND_GATE U10172 ( .I1(n9975), .I2(n9423), .O(n9424) );
  NAND_GATE U10173 ( .I1(n9971), .I2(n9424), .O(n9868) );
  NAND_GATE U10174 ( .I1(n9438), .I2(n9868), .O(n9864) );
  INV_GATE U10175 ( .I1(n9425), .O(n9426) );
  NAND_GATE U10176 ( .I1(n9426), .I2(n9429), .O(n9437) );
  NAND_GATE U10177 ( .I1(n9428), .I2(n9431), .O(n9435) );
  NAND_GATE U10178 ( .I1(n769), .I2(n9429), .O(n9430) );
  NAND_GATE U10179 ( .I1(n9431), .I2(n9430), .O(n9432) );
  NAND_GATE U10180 ( .I1(n9433), .I2(n9432), .O(n9434) );
  NAND_GATE U10181 ( .I1(n9435), .I2(n9434), .O(n9436) );
  NAND_GATE U10182 ( .I1(n9437), .I2(n9436), .O(n9867) );
  NAND_GATE U10183 ( .I1(n9868), .I2(n9867), .O(n9439) );
  NAND_GATE U10184 ( .I1(n9438), .I2(n9867), .O(n9863) );
  NAND3_GATE U10185 ( .I1(n9864), .I2(n9439), .I3(n9863), .O(n9992) );
  NAND_GATE U10186 ( .I1(n9990), .I2(n9997), .O(n9440) );
  NAND_GATE U10187 ( .I1(n9992), .I2(n9440), .O(n9441) );
  NAND_GATE U10188 ( .I1(n9987), .I2(n9441), .O(n10009) );
  NAND_GATE U10189 ( .I1(n9455), .I2(n10009), .O(n10005) );
  INV_GATE U10190 ( .I1(n9442), .O(n9443) );
  NAND_GATE U10191 ( .I1(n9443), .I2(n9447), .O(n9454) );
  INV_GATE U10192 ( .I1(n9447), .O(n9444) );
  NAND_GATE U10193 ( .I1(n9445), .I2(n9444), .O(n9449) );
  NAND_GATE U10194 ( .I1(n9446), .I2(n9449), .O(n9452) );
  NAND_GATE U10195 ( .I1(n9452), .I2(n9451), .O(n9453) );
  NAND_GATE U10196 ( .I1(n9454), .I2(n9453), .O(n10008) );
  NAND_GATE U10197 ( .I1(n10009), .I2(n10008), .O(n9456) );
  NAND_GATE U10198 ( .I1(n9455), .I2(n10008), .O(n10004) );
  NAND3_GATE U10199 ( .I1(n10005), .I2(n9456), .I3(n10004), .O(n9856) );
  NAND_GATE U10200 ( .I1(n9860), .I2(n9853), .O(n9457) );
  NAND_GATE U10201 ( .I1(n9460), .I2(n9306), .O(n9461) );
  NAND_GATE U10202 ( .I1(n9462), .I2(n9461), .O(n9844) );
  NAND_GATE U10203 ( .I1(n9849), .I2(n9844), .O(n9464) );
  NAND_GATE U10204 ( .I1(B[12]), .I2(A[13]), .O(n9847) );
  INV_GATE U10205 ( .I1(n9847), .O(n9463) );
  NAND_GATE U10206 ( .I1(n9849), .I2(n9463), .O(n9843) );
  NAND3_GATE U10207 ( .I1(n9848), .I2(n9464), .I3(n9843), .O(n10029) );
  NAND_GATE U10208 ( .I1(n10025), .I2(n10022), .O(n9465) );
  NAND_GATE U10209 ( .I1(n10029), .I2(n9465), .O(n9466) );
  NAND_GATE U10210 ( .I1(n10028), .I2(n9466), .O(n9836) );
  NAND_GATE U10211 ( .I1(n9468), .I2(n9471), .O(n9831) );
  NAND_GATE U10212 ( .I1(n632), .I2(n9470), .O(n9471) );
  NAND_GATE U10213 ( .I1(n9472), .I2(n9471), .O(n9833) );
  NAND_GATE U10214 ( .I1(n9834), .I2(n9833), .O(n9473) );
  NAND_GATE U10215 ( .I1(n9831), .I2(n9473), .O(n9474) );
  NAND_GATE U10216 ( .I1(n9832), .I2(n9474), .O(n9828) );
  NAND_GATE U10217 ( .I1(n9836), .I2(n9828), .O(n9476) );
  NAND_GATE U10218 ( .I1(B[12]), .I2(A[15]), .O(n9838) );
  INV_GATE U10219 ( .I1(n9838), .O(n9475) );
  NAND_GATE U10220 ( .I1(n9475), .I2(n9828), .O(n9826) );
  NAND_GATE U10221 ( .I1(n9475), .I2(n9836), .O(n9827) );
  NAND_GATE U10222 ( .I1(n10040), .I2(n10039), .O(n9477) );
  NAND3_GATE U10223 ( .I1(n9809), .I2(n9808), .I3(n9814), .O(n9479) );
  NAND_GATE U10224 ( .I1(n9478), .I2(n9814), .O(n9819) );
  NAND3_GATE U10225 ( .I1(n9815), .I2(n9479), .I3(n9819), .O(n10053) );
  NAND_GATE U10226 ( .I1(n10055), .I2(n10052), .O(n9480) );
  NAND_GATE U10227 ( .I1(n10053), .I2(n9480), .O(n9481) );
  NAND_GATE U10228 ( .I1(n10051), .I2(n9481), .O(n9796) );
  NAND_GATE U10229 ( .I1(n9492), .I2(n9796), .O(n9802) );
  INV_GATE U10230 ( .I1(n9493), .O(n9483) );
  NAND3_GATE U10231 ( .I1(n9484), .I2(n9483), .I3(n9498), .O(n9486) );
  NAND_GATE U10232 ( .I1(n9484), .I2(n9483), .O(n9496) );
  NAND_GATE U10233 ( .I1(n9485), .I2(n9496), .O(n9488) );
  NAND3_GATE U10234 ( .I1(n9486), .I2(n9495), .I3(n9488), .O(n9487) );
  NAND_GATE U10235 ( .I1(n9490), .I2(n9487), .O(n9803) );
  NAND_GATE U10236 ( .I1(n9796), .I2(n9803), .O(n9500) );
  INV_GATE U10237 ( .I1(n9488), .O(n9489) );
  NAND_GATE U10238 ( .I1(n9490), .I2(n9489), .O(n9491) );
  AND_GATE U10239 ( .I1(n9492), .I2(n9491), .O(n9801) );
  NAND_GATE U10240 ( .I1(n9494), .I2(n9493), .O(n9495) );
  NAND_GATE U10241 ( .I1(n9496), .I2(n9495), .O(n9497) );
  NAND_GATE U10242 ( .I1(n9498), .I2(n9497), .O(n9800) );
  NAND_GATE U10243 ( .I1(n9801), .I2(n9800), .O(n9499) );
  NAND3_GATE U10244 ( .I1(n9802), .I2(n9500), .I3(n9499), .O(n10072) );
  NAND_GATE U10245 ( .I1(n10078), .I2(n10069), .O(n9501) );
  NAND_GATE U10246 ( .I1(n10072), .I2(n9501), .O(n9502) );
  NAND_GATE U10247 ( .I1(n10071), .I2(n9502), .O(n9785) );
  NAND_GATE U10248 ( .I1(n9504), .I2(n9785), .O(n9789) );
  INV_GATE U10249 ( .I1(n9506), .O(n9508) );
  NAND_GATE U10250 ( .I1(n9503), .I2(n9509), .O(n9788) );
  NAND3_GATE U10251 ( .I1(n9506), .I2(n9503), .I3(n9505), .O(n9792) );
  NAND_GATE U10252 ( .I1(n9506), .I2(n9505), .O(n9510) );
  NAND_GATE U10253 ( .I1(n9508), .I2(n9507), .O(n9509) );
  NAND_GATE U10254 ( .I1(n9510), .I2(n9509), .O(n9778) );
  NAND_GATE U10255 ( .I1(n9779), .I2(n9778), .O(n9787) );
  NAND_GATE U10256 ( .I1(n916), .I2(n9787), .O(n9512) );
  NAND3_GATE U10257 ( .I1(n9785), .I2(n9780), .I3(n9787), .O(n9511) );
  NAND3_GATE U10258 ( .I1(n9789), .I2(n9512), .I3(n9511), .O(n9774) );
  NAND_GATE U10259 ( .I1(n9513), .I2(n9774), .O(n9771) );
  AND_GATE U10260 ( .I1(n9773), .I2(n9771), .O(n9517) );
  NAND_GATE U10261 ( .I1(n9515), .I2(n9514), .O(n9772) );
  NAND_GATE U10262 ( .I1(n9774), .I2(n9772), .O(n9516) );
  NAND_GATE U10263 ( .I1(n9517), .I2(n9516), .O(n9753) );
  NAND4_GATE U10264 ( .I1(n9750), .I2(n9752), .I3(n9759), .I4(n9753), .O(n9519) );
  NAND_GATE U10265 ( .I1(B[12]), .I2(A[23]), .O(n10091) );
  INV_GATE U10266 ( .I1(n10091), .O(n9758) );
  NAND3_GATE U10267 ( .I1(n949), .I2(n9759), .I3(n9758), .O(n9518) );
  NAND3_GATE U10268 ( .I1(n9519), .I2(n9518), .I3(n9756), .O(n9742) );
  NAND_GATE U10269 ( .I1(n9736), .I2(n9742), .O(n9737) );
  INV_GATE U10270 ( .I1(n9529), .O(n9523) );
  NAND_GATE U10271 ( .I1(n9524), .I2(n9523), .O(n9520) );
  NAND_GATE U10272 ( .I1(n9521), .I2(n9520), .O(n9527) );
  NAND_GATE U10273 ( .I1(n4), .I2(n9529), .O(n9526) );
  NAND3_GATE U10274 ( .I1(n9524), .I2(n9523), .I3(n9522), .O(n9525) );
  NAND3_GATE U10275 ( .I1(n9527), .I2(n9526), .I3(n9525), .O(n9532) );
  INV_GATE U10276 ( .I1(n9528), .O(n9530) );
  NAND_GATE U10277 ( .I1(n9530), .I2(n9529), .O(n9531) );
  NAND_GATE U10278 ( .I1(n9532), .I2(n9531), .O(n9741) );
  NAND_GATE U10279 ( .I1(n9736), .I2(n9741), .O(n9534) );
  NAND_GATE U10280 ( .I1(n9742), .I2(n9741), .O(n9533) );
  NAND3_GATE U10281 ( .I1(n9737), .I2(n9534), .I3(n9533), .O(n9731) );
  NAND_GATE U10282 ( .I1(n9723), .I2(n9731), .O(n9724) );
  NAND3_GATE U10283 ( .I1(n9535), .I2(n9536), .I3(n9537), .O(n9718) );
  NAND_GATE U10284 ( .I1(n9535), .I2(n9539), .O(n9717) );
  NAND_GATE U10285 ( .I1(n9538), .I2(n176), .O(n9539) );
  NAND_GATE U10286 ( .I1(n9540), .I2(n9539), .O(n9719) );
  NAND_GATE U10287 ( .I1(n9720), .I2(n9719), .O(n9541) );
  NAND_GATE U10288 ( .I1(n9717), .I2(n9541), .O(n9542) );
  NAND_GATE U10289 ( .I1(n9718), .I2(n9542), .O(n9725) );
  NAND_GATE U10290 ( .I1(n9731), .I2(n9725), .O(n9543) );
  NAND3_GATE U10291 ( .I1(n9724), .I2(n9732), .I3(n9543), .O(n9706) );
  NAND_GATE U10292 ( .I1(n9710), .I2(n9706), .O(n9712) );
  INV_GATE U10293 ( .I1(n9544), .O(n9545) );
  NAND_GATE U10294 ( .I1(n9545), .I2(n9548), .O(n9557) );
  NAND_GATE U10295 ( .I1(n9552), .I2(n9551), .O(n9546) );
  NAND_GATE U10296 ( .I1(n9547), .I2(n9546), .O(n9555) );
  NAND_GATE U10297 ( .I1(n9549), .I2(n9548), .O(n9554) );
  NAND3_GATE U10298 ( .I1(n9552), .I2(n9551), .I3(n9550), .O(n9553) );
  NAND3_GATE U10299 ( .I1(n9555), .I2(n9554), .I3(n9553), .O(n9556) );
  NAND_GATE U10300 ( .I1(n9557), .I2(n9556), .O(n9713) );
  NAND_GATE U10301 ( .I1(n9710), .I2(n9713), .O(n9559) );
  NAND_GATE U10302 ( .I1(n9706), .I2(n9713), .O(n9558) );
  NAND3_GATE U10303 ( .I1(n9712), .I2(n9559), .I3(n9558), .O(n9700) );
  NAND_GATE U10304 ( .I1(n9570), .I2(n9700), .O(n9694) );
  NAND_GATE U10305 ( .I1(n9564), .I2(n513), .O(n9561) );
  NAND_GATE U10306 ( .I1(n9562), .I2(n9561), .O(n9569) );
  NAND_GATE U10307 ( .I1(n630), .I2(n9563), .O(n9565) );
  NAND_GATE U10308 ( .I1(n9565), .I2(n9561), .O(n9566) );
  NAND_GATE U10309 ( .I1(n9567), .I2(n9566), .O(n9568) );
  NAND_GATE U10310 ( .I1(n9569), .I2(n9568), .O(n9699) );
  NAND_GATE U10311 ( .I1(n9701), .I2(n9699), .O(n9697) );
  NAND_GATE U10312 ( .I1(n9570), .I2(n9697), .O(n9693) );
  NAND_GATE U10313 ( .I1(n9700), .I2(n9697), .O(n9571) );
  NAND3_GATE U10314 ( .I1(n9694), .I2(n9693), .I3(n9571), .O(n9686) );
  NAND_GATE U10315 ( .I1(n9584), .I2(n9686), .O(n9688) );
  INV_GATE U10316 ( .I1(n9572), .O(n9573) );
  NAND_GATE U10317 ( .I1(n9573), .I2(n9575), .O(n9583) );
  NAND_GATE U10318 ( .I1(n9574), .I2(n9579), .O(n9581) );
  NAND_GATE U10319 ( .I1(n9578), .I2(n9577), .O(n9579) );
  NAND_GATE U10320 ( .I1(n9583), .I2(n9582), .O(n9689) );
  NAND_GATE U10321 ( .I1(n9584), .I2(n9689), .O(n9687) );
  NAND_GATE U10322 ( .I1(n9686), .I2(n9689), .O(n9585) );
  NAND3_GATE U10323 ( .I1(n9688), .I2(n9687), .I3(n9585), .O(n9676) );
  NAND_GATE U10324 ( .I1(n9599), .I2(n9676), .O(n9678) );
  INV_GATE U10325 ( .I1(n9586), .O(n9587) );
  NAND_GATE U10326 ( .I1(n9587), .I2(n9590), .O(n9598) );
  NAND_GATE U10327 ( .I1(n9591), .I2(n662), .O(n9588) );
  NAND_GATE U10328 ( .I1(n9589), .I2(n9588), .O(n9596) );
  NAND_GATE U10329 ( .I1(n830), .I2(n9590), .O(n9592) );
  NAND_GATE U10330 ( .I1(n9592), .I2(n9588), .O(n9593) );
  NAND_GATE U10331 ( .I1(n9594), .I2(n9593), .O(n9595) );
  NAND_GATE U10332 ( .I1(n9596), .I2(n9595), .O(n9597) );
  NAND_GATE U10333 ( .I1(n9598), .I2(n9597), .O(n9679) );
  NAND_GATE U10334 ( .I1(n9599), .I2(n9679), .O(n9677) );
  NAND_GATE U10335 ( .I1(n9676), .I2(n9679), .O(n9600) );
  NAND3_GATE U10336 ( .I1(n9678), .I2(n9677), .I3(n9600), .O(n9667) );
  NAND_GATE U10337 ( .I1(n9615), .I2(n9667), .O(n9663) );
  INV_GATE U10338 ( .I1(n9601), .O(n9602) );
  NAND_GATE U10339 ( .I1(n9602), .I2(n9605), .O(n9614) );
  INV_GATE U10340 ( .I1(n9605), .O(n9606) );
  NAND_GATE U10341 ( .I1(n9607), .I2(n9606), .O(n9603) );
  NAND_GATE U10342 ( .I1(n9604), .I2(n9603), .O(n9612) );
  NAND_GATE U10343 ( .I1(n617), .I2(n9605), .O(n9608) );
  NAND_GATE U10344 ( .I1(n9608), .I2(n9603), .O(n9609) );
  NAND_GATE U10345 ( .I1(n9610), .I2(n9609), .O(n9611) );
  NAND_GATE U10346 ( .I1(n9612), .I2(n9611), .O(n9613) );
  NAND_GATE U10347 ( .I1(n9614), .I2(n9613), .O(n9666) );
  NAND_GATE U10348 ( .I1(n9667), .I2(n9666), .O(n9616) );
  NAND3_GATE U10349 ( .I1(n9663), .I2(n9662), .I3(n9616), .O(n9656) );
  NAND_GATE U10350 ( .I1(n9631), .I2(n9656), .O(n9652) );
  INV_GATE U10351 ( .I1(n9617), .O(n9618) );
  NAND_GATE U10352 ( .I1(n9618), .I2(n9621), .O(n9630) );
  NAND_GATE U10353 ( .I1(n9620), .I2(n9624), .O(n9628) );
  NAND_GATE U10354 ( .I1(n9622), .I2(n9621), .O(n9623) );
  NAND_GATE U10355 ( .I1(n9624), .I2(n9623), .O(n9625) );
  NAND_GATE U10356 ( .I1(n9626), .I2(n9625), .O(n9627) );
  NAND_GATE U10357 ( .I1(n9628), .I2(n9627), .O(n9629) );
  NAND_GATE U10358 ( .I1(n9630), .I2(n9629), .O(n9655) );
  NAND_GATE U10359 ( .I1(n9656), .I2(n9655), .O(n9632) );
  NAND3_GATE U10360 ( .I1(n9652), .I2(n9651), .I3(n9632), .O(n15333) );
  INV_GATE U10361 ( .I1(n15333), .O(n9647) );
  INV_GATE U10362 ( .I1(n9633), .O(n9634) );
  NAND_GATE U10363 ( .I1(n9634), .I2(n9637), .O(n9646) );
  NAND_GATE U10364 ( .I1(n9636), .I2(n9640), .O(n9644) );
  NAND_GATE U10365 ( .I1(n9638), .I2(n9637), .O(n9639) );
  NAND_GATE U10366 ( .I1(n9640), .I2(n9639), .O(n9641) );
  NAND_GATE U10367 ( .I1(n9642), .I2(n9641), .O(n9643) );
  NAND_GATE U10368 ( .I1(n9644), .I2(n9643), .O(n9645) );
  NAND_GATE U10369 ( .I1(n9646), .I2(n9645), .O(n15332) );
  NAND_GATE U10370 ( .I1(n9647), .I2(n15332), .O(n9650) );
  INV_GATE U10371 ( .I1(n15332), .O(n9648) );
  NAND_GATE U10372 ( .I1(n15333), .I2(n9648), .O(n9649) );
  NAND_GATE U10373 ( .I1(n9650), .I2(n9649), .O(\A1[42] ) );
  OR_GATE U10374 ( .I1(n9651), .I2(n9656), .O(n9654) );
  OR_GATE U10375 ( .I1(n9655), .I2(n9652), .O(n9653) );
  AND_GATE U10376 ( .I1(n9654), .I2(n9653), .O(n9661) );
  NAND_GATE U10377 ( .I1(n902), .I2(n9655), .O(n9659) );
  NAND3_GATE U10378 ( .I1(n9659), .I2(n9658), .I3(n9657), .O(n9660) );
  OR_GATE U10379 ( .I1(n9662), .I2(n9667), .O(n9665) );
  OR_GATE U10380 ( .I1(n9666), .I2(n9663), .O(n9664) );
  AND_GATE U10381 ( .I1(n9665), .I2(n9664), .O(n9672) );
  NAND_GATE U10382 ( .I1(n890), .I2(n9666), .O(n9670) );
  NAND3_GATE U10383 ( .I1(n9670), .I2(n9669), .I3(n9668), .O(n9671) );
  NAND_GATE U10384 ( .I1(n9672), .I2(n9671), .O(n10490) );
  NAND_GATE U10385 ( .I1(B[11]), .I2(A[31]), .O(n15336) );
  INV_GATE U10386 ( .I1(n15336), .O(n10491) );
  NAND_GATE U10387 ( .I1(n10487), .I2(n10491), .O(n10492) );
  NAND_GATE U10388 ( .I1(n889), .I2(n9679), .O(n9675) );
  NAND3_GATE U10389 ( .I1(n9675), .I2(n9674), .I3(n9673), .O(n9682) );
  OR_GATE U10390 ( .I1(n9677), .I2(n9676), .O(n9681) );
  OR_GATE U10391 ( .I1(n9679), .I2(n9678), .O(n9680) );
  NAND3_GATE U10392 ( .I1(n9682), .I2(n9681), .I3(n9680), .O(n10477) );
  INV_GATE U10393 ( .I1(n10477), .O(n10476) );
  NAND_GATE U10394 ( .I1(B[11]), .I2(A[30]), .O(n10480) );
  INV_GATE U10395 ( .I1(n10480), .O(n10474) );
  NAND_GATE U10396 ( .I1(n10476), .I2(n10474), .O(n10471) );
  NAND_GATE U10397 ( .I1(n1198), .I2(n9689), .O(n9685) );
  NAND3_GATE U10398 ( .I1(n9685), .I2(n9684), .I3(n9683), .O(n9692) );
  OR_GATE U10399 ( .I1(n9687), .I2(n9686), .O(n9691) );
  OR_GATE U10400 ( .I1(n9689), .I2(n9688), .O(n9690) );
  NAND3_GATE U10401 ( .I1(n9692), .I2(n9691), .I3(n9690), .O(n10465) );
  NAND_GATE U10402 ( .I1(B[11]), .I2(A[29]), .O(n10506) );
  OR_GATE U10403 ( .I1(n9693), .I2(n9700), .O(n9696) );
  OR_GATE U10404 ( .I1(n9697), .I2(n9694), .O(n9695) );
  INV_GATE U10405 ( .I1(n9700), .O(n9698) );
  NAND_GATE U10406 ( .I1(n9698), .I2(n9697), .O(n9704) );
  NAND3_GATE U10407 ( .I1(n9701), .I2(n9700), .I3(n9699), .O(n9703) );
  NAND3_GATE U10408 ( .I1(n9704), .I2(n9703), .I3(n9702), .O(n9705) );
  INV_GATE U10409 ( .I1(n10456), .O(n10454) );
  NAND_GATE U10410 ( .I1(B[11]), .I2(A[28]), .O(n10457) );
  INV_GATE U10411 ( .I1(n10457), .O(n10452) );
  NAND_GATE U10412 ( .I1(n10454), .I2(n10452), .O(n10450) );
  NAND_GATE U10413 ( .I1(B[11]), .I2(A[27]), .O(n10936) );
  INV_GATE U10414 ( .I1(n10936), .O(n10441) );
  NAND_GATE U10415 ( .I1(n9711), .I2(n9713), .O(n9709) );
  NAND3_GATE U10416 ( .I1(n9709), .I2(n9708), .I3(n9707), .O(n9716) );
  NAND3_GATE U10417 ( .I1(n9711), .I2(n9713), .I3(n9710), .O(n9715) );
  OR_GATE U10418 ( .I1(n9713), .I2(n9712), .O(n9714) );
  NAND3_GATE U10419 ( .I1(n9716), .I2(n9715), .I3(n9714), .O(n10445) );
  NAND_GATE U10420 ( .I1(n10441), .I2(n10443), .O(n10105) );
  NAND_GATE U10421 ( .I1(B[11]), .I2(A[26]), .O(n10530) );
  INV_GATE U10422 ( .I1(n10530), .O(n10432) );
  NAND_GATE U10423 ( .I1(n9718), .I2(n588), .O(n9722) );
  NAND_GATE U10424 ( .I1(n9722), .I2(n9541), .O(n9721) );
  NAND_GATE U10425 ( .I1(n9731), .I2(n9721), .O(n9729) );
  NAND3_GATE U10426 ( .I1(n218), .I2(n9722), .I3(n9541), .O(n9728) );
  NAND3_GATE U10427 ( .I1(n9729), .I2(n9728), .I3(n9730), .O(n9727) );
  NAND3_GATE U10428 ( .I1(n9723), .I2(n218), .I3(n9725), .O(n9726) );
  NAND3_GATE U10429 ( .I1(n9727), .I2(n9726), .I3(n9734), .O(n10435) );
  NAND_GATE U10430 ( .I1(n10432), .I2(n10434), .O(n10102) );
  NAND4_GATE U10431 ( .I1(n9730), .I2(n9729), .I3(n10530), .I4(n9728), .O(
        n10100) );
  OR_GATE U10432 ( .I1(n9732), .I2(n9731), .O(n9733) );
  NAND_GATE U10433 ( .I1(n9734), .I2(n9733), .O(n9735) );
  NAND_GATE U10434 ( .I1(n10530), .I2(n9735), .O(n10099) );
  NAND_GATE U10435 ( .I1(B[11]), .I2(A[25]), .O(n10545) );
  INV_GATE U10436 ( .I1(n10545), .O(n10120) );
  INV_GATE U10437 ( .I1(n9742), .O(n9740) );
  NAND3_GATE U10438 ( .I1(n9740), .I2(n9741), .I3(n9736), .O(n9739) );
  OR_GATE U10439 ( .I1(n9741), .I2(n9737), .O(n9738) );
  AND_GATE U10440 ( .I1(n9739), .I2(n9738), .O(n9747) );
  NAND_GATE U10441 ( .I1(n9740), .I2(n9741), .O(n9744) );
  NAND3_GATE U10442 ( .I1(n9745), .I2(n9744), .I3(n9743), .O(n9746) );
  NAND_GATE U10443 ( .I1(n9747), .I2(n9746), .O(n10115) );
  NAND_GATE U10444 ( .I1(n10120), .I2(n736), .O(n10098) );
  NAND_GATE U10445 ( .I1(B[11]), .I2(A[24]), .O(n10568) );
  INV_GATE U10446 ( .I1(n10568), .O(n10420) );
  NAND_GATE U10447 ( .I1(n9749), .I2(n9748), .O(n9751) );
  NAND3_GATE U10448 ( .I1(n9752), .I2(n9751), .I3(n9750), .O(n9754) );
  NAND3_GATE U10449 ( .I1(n9754), .I2(n9755), .I3(n9753), .O(n10090) );
  NAND_GATE U10450 ( .I1(n9755), .I2(n9754), .O(n9757) );
  NAND_GATE U10451 ( .I1(n19), .I2(n9757), .O(n10089) );
  AND3_GATE U10452 ( .I1(n10090), .I2(n10089), .I3(n10091), .O(n9762) );
  OR_GATE U10453 ( .I1(n9757), .I2(n9756), .O(n9761) );
  NAND4_GATE U10454 ( .I1(n19), .I2(n9759), .I3(n949), .I4(n9758), .O(n9760)
         );
  NAND_GATE U10455 ( .I1(n9761), .I2(n9760), .O(n10092) );
  OR_GATE U10456 ( .I1(n9762), .I2(n10092), .O(n10424) );
  INV_GATE U10457 ( .I1(n10424), .O(n10423) );
  NAND_GATE U10458 ( .I1(n10420), .I2(n10423), .O(n10421) );
  NAND_GATE U10459 ( .I1(n9764), .I2(n9763), .O(n9765) );
  NAND_GATE U10460 ( .I1(n9766), .I2(n9765), .O(n9767) );
  OR_GATE U10461 ( .I1(n9767), .I2(n9774), .O(n9770) );
  NAND_GATE U10462 ( .I1(n9774), .I2(n9767), .O(n9769) );
  NAND3_GATE U10463 ( .I1(n9770), .I2(n9769), .I3(n9768), .O(n9777) );
  OR_GATE U10464 ( .I1(n9772), .I2(n9771), .O(n9776) );
  OR_GATE U10465 ( .I1(n9774), .I2(n9773), .O(n9775) );
  NAND3_GATE U10466 ( .I1(n9777), .I2(n9776), .I3(n9775), .O(n10413) );
  NAND_GATE U10467 ( .I1(B[11]), .I2(A[23]), .O(n10593) );
  INV_GATE U10468 ( .I1(n10593), .O(n10415) );
  NAND_GATE U10469 ( .I1(n806), .I2(n10415), .O(n10088) );
  NAND_GATE U10470 ( .I1(B[11]), .I2(A[22]), .O(n10122) );
  INV_GATE U10471 ( .I1(n10122), .O(n10404) );
  NAND_GATE U10472 ( .I1(n9780), .I2(n9787), .O(n9781) );
  OR_GATE U10473 ( .I1(n9781), .I2(n9785), .O(n9784) );
  NAND_GATE U10474 ( .I1(n9785), .I2(n9781), .O(n9783) );
  NAND3_GATE U10475 ( .I1(n9784), .I2(n9783), .I3(n9782), .O(n9795) );
  INV_GATE U10476 ( .I1(n9785), .O(n9786) );
  NAND3_GATE U10477 ( .I1(n916), .I2(n9787), .I3(n9786), .O(n9794) );
  NAND_GATE U10478 ( .I1(n9788), .I2(n9787), .O(n9791) );
  INV_GATE U10479 ( .I1(n9789), .O(n9790) );
  NAND3_GATE U10480 ( .I1(n9792), .I2(n9791), .I3(n9790), .O(n9793) );
  NAND3_GATE U10481 ( .I1(n9795), .I2(n9794), .I3(n9793), .O(n10125) );
  NAND_GATE U10482 ( .I1(n10404), .I2(n10123), .O(n10085) );
  NAND_GATE U10483 ( .I1(B[11]), .I2(A[21]), .O(n10136) );
  INV_GATE U10484 ( .I1(n10136), .O(n10081) );
  NAND_GATE U10485 ( .I1(n936), .I2(n9803), .O(n9799) );
  NAND3_GATE U10486 ( .I1(n9799), .I2(n9798), .I3(n9797), .O(n9806) );
  NAND3_GATE U10487 ( .I1(n9801), .I2(n9800), .I3(n936), .O(n9805) );
  OR_GATE U10488 ( .I1(n9803), .I2(n9802), .O(n9804) );
  NAND3_GATE U10489 ( .I1(n9806), .I2(n9805), .I3(n9804), .O(n10394) );
  NAND_GATE U10490 ( .I1(B[11]), .I2(A[20]), .O(n10615) );
  INV_GATE U10491 ( .I1(n10615), .O(n10392) );
  NAND_GATE U10492 ( .I1(n670), .I2(n10392), .O(n10391) );
  INV_GATE U10493 ( .I1(n9814), .O(n9807) );
  NAND3_GATE U10494 ( .I1(n9809), .I2(n9808), .I3(n9807), .O(n9813) );
  NAND_GATE U10495 ( .I1(n9809), .I2(n9808), .O(n9810) );
  NAND_GATE U10496 ( .I1(n9814), .I2(n9810), .O(n9812) );
  NAND3_GATE U10497 ( .I1(n9813), .I2(n9812), .I3(n9811), .O(n9825) );
  OR_GATE U10498 ( .I1(n9815), .I2(n9814), .O(n9824) );
  NAND_GATE U10499 ( .I1(n9818), .I2(n9808), .O(n9821) );
  INV_GATE U10500 ( .I1(n9819), .O(n9820) );
  NAND3_GATE U10501 ( .I1(n9822), .I2(n9821), .I3(n9820), .O(n9823) );
  NAND3_GATE U10502 ( .I1(n9825), .I2(n9824), .I3(n9823), .O(n10380) );
  NAND_GATE U10503 ( .I1(B[11]), .I2(A[18]), .O(n10387) );
  INV_GATE U10504 ( .I1(n10387), .O(n10381) );
  NAND_GATE U10505 ( .I1(n741), .I2(n10381), .O(n10382) );
  NAND_GATE U10506 ( .I1(B[11]), .I2(A[16]), .O(n10653) );
  INV_GATE U10507 ( .I1(n10653), .O(n10164) );
  OR_GATE U10508 ( .I1(n9826), .I2(n9836), .O(n9830) );
  OR_GATE U10509 ( .I1(n9828), .I2(n9827), .O(n9829) );
  AND_GATE U10510 ( .I1(n9830), .I2(n9829), .O(n9842) );
  NAND_GATE U10511 ( .I1(n9837), .I2(n9473), .O(n9835) );
  NAND_GATE U10512 ( .I1(n9836), .I2(n9835), .O(n9840) );
  NAND3_GATE U10513 ( .I1(n9840), .I2(n9839), .I3(n9838), .O(n9841) );
  NAND_GATE U10514 ( .I1(n10164), .I2(n1328), .O(n10037) );
  NAND_GATE U10515 ( .I1(B[11]), .I2(A[15]), .O(n10175) );
  INV_GATE U10516 ( .I1(n10175), .O(n10033) );
  NAND_GATE U10517 ( .I1(B[11]), .I2(A[14]), .O(n10180) );
  INV_GATE U10518 ( .I1(n10180), .O(n10183) );
  OR_GATE U10519 ( .I1(n9843), .I2(n9844), .O(n9852) );
  NAND_GATE U10520 ( .I1(n941), .I2(n9844), .O(n9846) );
  NAND3_GATE U10521 ( .I1(n9847), .I2(n9846), .I3(n9845), .O(n9851) );
  OR_GATE U10522 ( .I1(n9849), .I2(n9848), .O(n9850) );
  NAND3_GATE U10523 ( .I1(n9852), .I2(n9851), .I3(n9850), .O(n10181) );
  NAND_GATE U10524 ( .I1(n1353), .I2(n9856), .O(n9854) );
  NAND3_GATE U10525 ( .I1(n9855), .I2(n9854), .I3(n9858), .O(n9862) );
  NAND_GATE U10526 ( .I1(n1197), .I2(n9856), .O(n9857) );
  NAND_GATE U10527 ( .I1(n9858), .I2(n9857), .O(n9859) );
  NAND_GATE U10528 ( .I1(n9860), .I2(n9859), .O(n9861) );
  NAND_GATE U10529 ( .I1(n9862), .I2(n9861), .O(n10194) );
  INV_GATE U10530 ( .I1(n10194), .O(n10193) );
  NAND_GATE U10531 ( .I1(B[11]), .I2(A[13]), .O(n10195) );
  NAND_GATE U10532 ( .I1(B[11]), .I2(A[12]), .O(n10360) );
  INV_GATE U10533 ( .I1(n10360), .O(n10355) );
  NAND_GATE U10534 ( .I1(B[11]), .I2(A[11]), .O(n10209) );
  INV_GATE U10535 ( .I1(n10209), .O(n10002) );
  OR_GATE U10536 ( .I1(n9863), .I2(n9868), .O(n9866) );
  OR_GATE U10537 ( .I1(n9867), .I2(n9864), .O(n9865) );
  AND_GATE U10538 ( .I1(n9866), .I2(n9865), .O(n9873) );
  NAND_GATE U10539 ( .I1(n986), .I2(n9867), .O(n9871) );
  NAND3_GATE U10540 ( .I1(n9871), .I2(n9870), .I3(n9869), .O(n9872) );
  NAND_GATE U10541 ( .I1(n9873), .I2(n9872), .O(n10216) );
  NAND_GATE U10542 ( .I1(B[11]), .I2(A[10]), .O(n10220) );
  INV_GATE U10543 ( .I1(n10220), .O(n10217) );
  NAND_GATE U10544 ( .I1(n552), .I2(n10217), .O(n10213) );
  NAND_GATE U10545 ( .I1(B[11]), .I2(A[9]), .O(n10343) );
  INV_GATE U10546 ( .I1(n10343), .O(n9983) );
  OR_GATE U10547 ( .I1(n9874), .I2(n9879), .O(n9877) );
  OR_GATE U10548 ( .I1(n9878), .I2(n9875), .O(n9876) );
  AND_GATE U10549 ( .I1(n9877), .I2(n9876), .O(n9884) );
  NAND_GATE U10550 ( .I1(n974), .I2(n9878), .O(n9882) );
  NAND3_GATE U10551 ( .I1(n9882), .I2(n9881), .I3(n9880), .O(n9883) );
  NAND_GATE U10552 ( .I1(n9884), .I2(n9883), .O(n10228) );
  INV_GATE U10553 ( .I1(n10228), .O(n10231) );
  NAND_GATE U10554 ( .I1(B[11]), .I2(A[8]), .O(n10233) );
  INV_GATE U10555 ( .I1(n10233), .O(n10229) );
  NAND_GATE U10556 ( .I1(n10231), .I2(n10229), .O(n10225) );
  INV_GATE U10557 ( .I1(n9885), .O(n9886) );
  NAND_GATE U10558 ( .I1(n9886), .I2(n9890), .O(n9899) );
  INV_GATE U10559 ( .I1(n9890), .O(n9887) );
  NAND_GATE U10560 ( .I1(n9888), .I2(n9887), .O(n9893) );
  NAND_GATE U10561 ( .I1(n9889), .I2(n9893), .O(n9897) );
  NAND_GATE U10562 ( .I1(n9891), .I2(n9890), .O(n9892) );
  NAND_GATE U10563 ( .I1(n9893), .I2(n9892), .O(n9894) );
  NAND_GATE U10564 ( .I1(n9895), .I2(n9894), .O(n9896) );
  NAND_GATE U10565 ( .I1(n9897), .I2(n9896), .O(n9898) );
  NAND_GATE U10566 ( .I1(n9899), .I2(n9898), .O(n10242) );
  INV_GATE U10567 ( .I1(n9900), .O(n9901) );
  NAND_GATE U10568 ( .I1(n9906), .I2(n9901), .O(n9914) );
  INV_GATE U10569 ( .I1(n9906), .O(n9903) );
  NAND_GATE U10570 ( .I1(n9903), .I2(n9902), .O(n9908) );
  NAND_GATE U10571 ( .I1(n9904), .I2(n9908), .O(n9912) );
  NAND_GATE U10572 ( .I1(n9906), .I2(n9905), .O(n9907) );
  NAND_GATE U10573 ( .I1(n9908), .I2(n9907), .O(n9909) );
  NAND_GATE U10574 ( .I1(n9910), .I2(n9909), .O(n9911) );
  NAND_GATE U10575 ( .I1(n9912), .I2(n9911), .O(n9913) );
  NAND_GATE U10576 ( .I1(n9914), .I2(n9913), .O(n10268) );
  OR_GATE U10577 ( .I1(n9915), .I2(n9917), .O(n9928) );
  NAND_GATE U10578 ( .I1(n9917), .I2(n9916), .O(n9922) );
  NAND_GATE U10579 ( .I1(n9918), .I2(n9922), .O(n9926) );
  NAND_GATE U10580 ( .I1(n9920), .I2(n9919), .O(n9921) );
  NAND_GATE U10581 ( .I1(n9922), .I2(n9921), .O(n9923) );
  NAND_GATE U10582 ( .I1(n9924), .I2(n9923), .O(n9925) );
  NAND_GATE U10583 ( .I1(n9926), .I2(n9925), .O(n9927) );
  NAND_GATE U10584 ( .I1(n9928), .I2(n9927), .O(n10294) );
  NAND3_GATE U10585 ( .I1(B[11]), .I2(B[12]), .I3(n1196), .O(n10303) );
  INV_GATE U10586 ( .I1(n10303), .O(n10306) );
  NAND_GATE U10587 ( .I1(n1376), .I2(A[0]), .O(n9929) );
  NAND_GATE U10588 ( .I1(n14781), .I2(n9929), .O(n9930) );
  NAND_GATE U10589 ( .I1(B[13]), .I2(n9930), .O(n9934) );
  NAND_GATE U10590 ( .I1(n1377), .I2(A[1]), .O(n9931) );
  NAND_GATE U10591 ( .I1(n14784), .I2(n9931), .O(n9932) );
  NAND_GATE U10592 ( .I1(B[12]), .I2(n9932), .O(n9933) );
  NAND_GATE U10593 ( .I1(n9934), .I2(n9933), .O(n10305) );
  INV_GATE U10594 ( .I1(n10305), .O(n10302) );
  NAND_GATE U10595 ( .I1(B[11]), .I2(A[2]), .O(n10310) );
  NAND_GATE U10596 ( .I1(n10302), .I2(n10310), .O(n9935) );
  NAND_GATE U10597 ( .I1(n10306), .I2(n9935), .O(n9936) );
  INV_GATE U10598 ( .I1(n10310), .O(n10304) );
  NAND_GATE U10599 ( .I1(n10305), .I2(n10304), .O(n10301) );
  NAND_GATE U10600 ( .I1(n9936), .I2(n10301), .O(n10295) );
  NAND_GATE U10601 ( .I1(n10294), .I2(n10295), .O(n9938) );
  NAND_GATE U10602 ( .I1(B[11]), .I2(A[3]), .O(n10296) );
  INV_GATE U10603 ( .I1(n10296), .O(n9937) );
  NAND_GATE U10604 ( .I1(n10295), .I2(n9937), .O(n10291) );
  NAND_GATE U10605 ( .I1(n10294), .I2(n9937), .O(n10290) );
  NAND3_GATE U10606 ( .I1(n9938), .I2(n10291), .I3(n10290), .O(n10281) );
  NAND_GATE U10607 ( .I1(B[11]), .I2(A[4]), .O(n10285) );
  OR_GATE U10608 ( .I1(n9939), .I2(n9944), .O(n9942) );
  OR_GATE U10609 ( .I1(n9940), .I2(n9943), .O(n9941) );
  AND_GATE U10610 ( .I1(n9942), .I2(n9941), .O(n9949) );
  NAND_GATE U10611 ( .I1(n9943), .I2(n1170), .O(n9947) );
  NAND3_GATE U10612 ( .I1(n9947), .I2(n9946), .I3(n9945), .O(n9948) );
  NAND_GATE U10613 ( .I1(n9949), .I2(n9948), .O(n10277) );
  NAND_GATE U10614 ( .I1(n10285), .I2(n10277), .O(n9950) );
  NAND_GATE U10615 ( .I1(n10281), .I2(n9950), .O(n9951) );
  INV_GATE U10616 ( .I1(n10285), .O(n10279) );
  INV_GATE U10617 ( .I1(n10277), .O(n10280) );
  NAND_GATE U10618 ( .I1(n10279), .I2(n10280), .O(n10275) );
  NAND_GATE U10619 ( .I1(n9951), .I2(n10275), .O(n10269) );
  NAND_GATE U10620 ( .I1(n10268), .I2(n10269), .O(n9953) );
  NAND_GATE U10621 ( .I1(B[11]), .I2(A[5]), .O(n10270) );
  INV_GATE U10622 ( .I1(n10270), .O(n9952) );
  NAND_GATE U10623 ( .I1(n10269), .I2(n9952), .O(n10265) );
  NAND_GATE U10624 ( .I1(n10268), .I2(n9952), .O(n10264) );
  NAND3_GATE U10625 ( .I1(n9953), .I2(n10265), .I3(n10264), .O(n10255) );
  NAND_GATE U10626 ( .I1(B[11]), .I2(A[6]), .O(n10259) );
  OR_GATE U10627 ( .I1(n9954), .I2(n9959), .O(n9957) );
  OR_GATE U10628 ( .I1(n9955), .I2(n9958), .O(n9956) );
  AND_GATE U10629 ( .I1(n9957), .I2(n9956), .O(n9964) );
  NAND_GATE U10630 ( .I1(n9958), .I2(n1098), .O(n9962) );
  NAND3_GATE U10631 ( .I1(n9962), .I2(n9961), .I3(n9960), .O(n9963) );
  NAND_GATE U10632 ( .I1(n9964), .I2(n9963), .O(n10251) );
  NAND_GATE U10633 ( .I1(n10259), .I2(n10251), .O(n9965) );
  NAND_GATE U10634 ( .I1(n10255), .I2(n9965), .O(n9966) );
  INV_GATE U10635 ( .I1(n10259), .O(n10253) );
  INV_GATE U10636 ( .I1(n10251), .O(n10254) );
  NAND_GATE U10637 ( .I1(n10253), .I2(n10254), .O(n10249) );
  NAND_GATE U10638 ( .I1(n9966), .I2(n10249), .O(n10243) );
  NAND_GATE U10639 ( .I1(n10242), .I2(n10243), .O(n9968) );
  NAND_GATE U10640 ( .I1(B[11]), .I2(A[7]), .O(n10244) );
  INV_GATE U10641 ( .I1(n10244), .O(n9967) );
  NAND_GATE U10642 ( .I1(n10243), .I2(n9967), .O(n10239) );
  NAND_GATE U10643 ( .I1(n10242), .I2(n9967), .O(n10238) );
  NAND3_GATE U10644 ( .I1(n9968), .I2(n10239), .I3(n10238), .O(n10230) );
  NAND_GATE U10645 ( .I1(n10228), .I2(n10233), .O(n9969) );
  NAND_GATE U10646 ( .I1(n10230), .I2(n9969), .O(n9970) );
  NAND_GATE U10647 ( .I1(n10225), .I2(n9970), .O(n10342) );
  NAND_GATE U10648 ( .I1(n9983), .I2(n10342), .O(n10338) );
  INV_GATE U10649 ( .I1(n9971), .O(n9972) );
  NAND_GATE U10650 ( .I1(n9972), .I2(n9975), .O(n9982) );
  NAND_GATE U10651 ( .I1(n9974), .I2(n9977), .O(n9980) );
  NAND_GATE U10652 ( .I1(n633), .I2(n9975), .O(n9976) );
  NAND_GATE U10653 ( .I1(n9980), .I2(n9979), .O(n9981) );
  NAND_GATE U10654 ( .I1(n9982), .I2(n9981), .O(n10341) );
  NAND_GATE U10655 ( .I1(n10342), .I2(n10341), .O(n9984) );
  NAND_GATE U10656 ( .I1(n9983), .I2(n10341), .O(n10337) );
  NAND3_GATE U10657 ( .I1(n10338), .I2(n9984), .I3(n10337), .O(n10218) );
  NAND_GATE U10658 ( .I1(n10216), .I2(n10220), .O(n9985) );
  NAND_GATE U10659 ( .I1(n10218), .I2(n9985), .O(n9986) );
  NAND_GATE U10660 ( .I1(n10213), .I2(n9986), .O(n10208) );
  NAND_GATE U10661 ( .I1(n10002), .I2(n10208), .O(n10204) );
  INV_GATE U10662 ( .I1(n9987), .O(n9988) );
  NAND_GATE U10663 ( .I1(n9988), .I2(n9992), .O(n10001) );
  INV_GATE U10664 ( .I1(n9992), .O(n9989) );
  NAND_GATE U10665 ( .I1(n9990), .I2(n9989), .O(n9995) );
  NAND_GATE U10666 ( .I1(n9991), .I2(n9995), .O(n9999) );
  NAND_GATE U10667 ( .I1(n9993), .I2(n9992), .O(n9994) );
  NAND_GATE U10668 ( .I1(n9995), .I2(n9994), .O(n9996) );
  NAND_GATE U10669 ( .I1(n9997), .I2(n9996), .O(n9998) );
  NAND_GATE U10670 ( .I1(n9999), .I2(n9998), .O(n10000) );
  NAND_GATE U10671 ( .I1(n10001), .I2(n10000), .O(n10207) );
  NAND_GATE U10672 ( .I1(n10208), .I2(n10207), .O(n10003) );
  NAND_GATE U10673 ( .I1(n10002), .I2(n10207), .O(n10203) );
  NAND_GATE U10674 ( .I1(n10355), .I2(n10356), .O(n10353) );
  OR_GATE U10675 ( .I1(n10008), .I2(n10005), .O(n10006) );
  AND_GATE U10676 ( .I1(n10007), .I2(n10006), .O(n10014) );
  NAND_GATE U10677 ( .I1(n943), .I2(n10008), .O(n10012) );
  NAND3_GATE U10678 ( .I1(n10012), .I2(n10011), .I3(n10010), .O(n10013) );
  NAND_GATE U10679 ( .I1(n10014), .I2(n10013), .O(n10354) );
  NAND_GATE U10680 ( .I1(n10353), .I2(n10015), .O(n10199) );
  NAND_GATE U10681 ( .I1(n10193), .I2(n10199), .O(n10016) );
  NAND_GATE U10682 ( .I1(n10180), .I2(n10181), .O(n10017) );
  NAND_GATE U10683 ( .I1(n10187), .I2(n10017), .O(n10018) );
  NAND_GATE U10684 ( .I1(n10186), .I2(n10018), .O(n10166) );
  INV_GATE U10685 ( .I1(n10029), .O(n10021) );
  NAND_GATE U10686 ( .I1(n10022), .I2(n10021), .O(n10019) );
  NAND_GATE U10687 ( .I1(n10020), .I2(n10019), .O(n10027) );
  NAND_GATE U10688 ( .I1(n1203), .I2(n10029), .O(n10023) );
  NAND_GATE U10689 ( .I1(n10023), .I2(n10019), .O(n10024) );
  NAND_GATE U10690 ( .I1(n10025), .I2(n10024), .O(n10026) );
  NAND_GATE U10691 ( .I1(n10027), .I2(n10026), .O(n10032) );
  INV_GATE U10692 ( .I1(n10028), .O(n10030) );
  NAND_GATE U10693 ( .I1(n10030), .I2(n10029), .O(n10031) );
  NAND_GATE U10694 ( .I1(n10032), .I2(n10031), .O(n10167) );
  NAND_GATE U10695 ( .I1(n10166), .I2(n10167), .O(n10034) );
  NAND_GATE U10696 ( .I1(n10033), .I2(n10167), .O(n10170) );
  NAND3_GATE U10697 ( .I1(n10168), .I2(n10034), .I3(n10170), .O(n10165) );
  NAND_GATE U10698 ( .I1(n10653), .I2(n10163), .O(n10035) );
  NAND_GATE U10699 ( .I1(n10165), .I2(n10035), .O(n10036) );
  NAND_GATE U10700 ( .I1(n10037), .I2(n10036), .O(n10154) );
  NAND_GATE U10701 ( .I1(n1248), .I2(n10038), .O(n10045) );
  NAND3_GATE U10702 ( .I1(n10040), .I2(n755), .I3(n10039), .O(n10041) );
  NAND3_GATE U10703 ( .I1(n10043), .I2(n10042), .I3(n10041), .O(n10044) );
  NAND_GATE U10704 ( .I1(n10045), .I2(n10044), .O(n10155) );
  NAND_GATE U10705 ( .I1(n10154), .I2(n10155), .O(n10048) );
  NAND_GATE U10706 ( .I1(B[11]), .I2(A[17]), .O(n10158) );
  INV_GATE U10707 ( .I1(n10158), .O(n10151) );
  NAND_GATE U10708 ( .I1(n10154), .I2(n10151), .O(n10047) );
  NAND_GATE U10709 ( .I1(n10155), .I2(n10151), .O(n10046) );
  NAND3_GATE U10710 ( .I1(n10048), .I2(n10047), .I3(n10046), .O(n10383) );
  NAND_GATE U10711 ( .I1(n10380), .I2(n10387), .O(n10049) );
  NAND_GATE U10712 ( .I1(n10383), .I2(n10049), .O(n10050) );
  NAND_GATE U10713 ( .I1(n10382), .I2(n10050), .O(n10139) );
  INV_GATE U10714 ( .I1(n10053), .O(n10054) );
  NAND3_GATE U10715 ( .I1(n10055), .I2(n10054), .I3(n10052), .O(n10060) );
  NAND_GATE U10716 ( .I1(n672), .I2(n10053), .O(n10059) );
  NAND_GATE U10717 ( .I1(n10055), .I2(n10054), .O(n10056) );
  NAND_GATE U10718 ( .I1(n10057), .I2(n10056), .O(n10058) );
  NAND3_GATE U10719 ( .I1(n10060), .I2(n10059), .I3(n10058), .O(n10141) );
  NAND_GATE U10720 ( .I1(n10140), .I2(n10141), .O(n10146) );
  NAND_GATE U10721 ( .I1(n10139), .I2(n10146), .O(n10062) );
  NAND_GATE U10722 ( .I1(B[11]), .I2(A[19]), .O(n10142) );
  INV_GATE U10723 ( .I1(n10142), .O(n10147) );
  NAND_GATE U10724 ( .I1(n10146), .I2(n10147), .O(n10061) );
  NAND_GATE U10725 ( .I1(n10139), .I2(n10147), .O(n10145) );
  NAND3_GATE U10726 ( .I1(n10062), .I2(n10061), .I3(n10145), .O(n10395) );
  NAND_GATE U10727 ( .I1(n10394), .I2(n10615), .O(n10063) );
  NAND_GATE U10728 ( .I1(n10395), .I2(n10063), .O(n10064) );
  NAND_GATE U10729 ( .I1(n10391), .I2(n10064), .O(n10133) );
  NAND_GATE U10730 ( .I1(n10081), .I2(n10133), .O(n10129) );
  NAND_GATE U10731 ( .I1(n10069), .I2(n10068), .O(n10065) );
  NAND_GATE U10732 ( .I1(n10066), .I2(n10065), .O(n10074) );
  NAND_GATE U10733 ( .I1(n10067), .I2(n10072), .O(n10070) );
  NAND_GATE U10734 ( .I1(n10070), .I2(n10065), .O(n10077) );
  NAND_GATE U10735 ( .I1(n10074), .I2(n10079), .O(n10073) );
  NAND_GATE U10736 ( .I1(n10073), .I2(n10075), .O(n10132) );
  NAND_GATE U10737 ( .I1(n10133), .I2(n10132), .O(n10082) );
  INV_GATE U10738 ( .I1(n10074), .O(n10076) );
  NAND_GATE U10739 ( .I1(n10076), .I2(n10075), .O(n10080) );
  NAND_GATE U10740 ( .I1(n10078), .I2(n10077), .O(n10079) );
  NAND3_GATE U10741 ( .I1(n10081), .I2(n10080), .I3(n10079), .O(n10128) );
  NAND_GATE U10742 ( .I1(n10122), .I2(n10125), .O(n10083) );
  NAND_GATE U10743 ( .I1(n10124), .I2(n10083), .O(n10084) );
  NAND_GATE U10744 ( .I1(n10085), .I2(n10084), .O(n10416) );
  NAND_GATE U10745 ( .I1(n10413), .I2(n10593), .O(n10086) );
  NAND_GATE U10746 ( .I1(n10416), .I2(n10086), .O(n10087) );
  NAND_GATE U10747 ( .I1(n10088), .I2(n10087), .O(n10422) );
  NAND4_GATE U10748 ( .I1(n10091), .I2(n10090), .I3(n10568), .I4(n10089), .O(
        n10094) );
  NAND_GATE U10749 ( .I1(n10568), .I2(n10092), .O(n10093) );
  NAND3_GATE U10750 ( .I1(n10422), .I2(n10094), .I3(n10093), .O(n10095) );
  NAND_GATE U10751 ( .I1(n10545), .I2(n10115), .O(n10096) );
  NAND_GATE U10752 ( .I1(n10119), .I2(n10096), .O(n10097) );
  NAND3_GATE U10753 ( .I1(n10100), .I2(n10099), .I3(n10433), .O(n10101) );
  NAND_GATE U10754 ( .I1(n10102), .I2(n10101), .O(n10442) );
  NAND_GATE U10755 ( .I1(n10936), .I2(n10445), .O(n10103) );
  NAND_GATE U10756 ( .I1(n10442), .I2(n10103), .O(n10104) );
  NAND_GATE U10757 ( .I1(n10105), .I2(n10104), .O(n10453) );
  NAND_GATE U10758 ( .I1(n10456), .I2(n10457), .O(n10106) );
  NAND_GATE U10759 ( .I1(n10453), .I2(n10106), .O(n10107) );
  NAND_GATE U10760 ( .I1(n10450), .I2(n10107), .O(n10463) );
  NAND_GATE U10761 ( .I1(n10465), .I2(n10506), .O(n10108) );
  NAND_GATE U10762 ( .I1(n10477), .I2(n10480), .O(n10109) );
  NAND_GATE U10763 ( .I1(n10475), .I2(n10109), .O(n10110) );
  NAND_GATE U10764 ( .I1(n10490), .I2(n15336), .O(n10111) );
  NAND_GATE U10765 ( .I1(n10493), .I2(n10111), .O(n10112) );
  NAND_GATE U10766 ( .I1(n10492), .I2(n10112), .O(n10113) );
  AND_GATE U10767 ( .I1(n15334), .I2(n10114), .O(\A1[41] ) );
  NAND_GATE U10768 ( .I1(B[10]), .I2(A[31]), .O(n10503) );
  INV_GATE U10769 ( .I1(n10503), .O(n10485) );
  NAND_GATE U10770 ( .I1(B[10]), .I2(A[30]), .O(n10513) );
  INV_GATE U10771 ( .I1(n10513), .O(n10515) );
  NAND_GATE U10772 ( .I1(B[10]), .I2(A[29]), .O(n10981) );
  INV_GATE U10773 ( .I1(n10981), .O(n10461) );
  NAND_GATE U10774 ( .I1(B[10]), .I2(A[28]), .O(n10943) );
  INV_GATE U10775 ( .I1(n10943), .O(n10947) );
  NAND_GATE U10776 ( .I1(B[10]), .I2(A[27]), .O(n10535) );
  INV_GATE U10777 ( .I1(n10535), .O(n10538) );
  NAND_GATE U10778 ( .I1(B[10]), .I2(A[26]), .O(n10554) );
  INV_GATE U10779 ( .I1(n10554), .O(n10557) );
  NAND_GATE U10780 ( .I1(n10120), .I2(n10116), .O(n10546) );
  NAND_GATE U10781 ( .I1(n736), .I2(n10119), .O(n10117) );
  NAND_GATE U10782 ( .I1(n10115), .I2(n782), .O(n10116) );
  NAND_GATE U10783 ( .I1(n10117), .I2(n10116), .O(n10544) );
  NAND_GATE U10784 ( .I1(n10545), .I2(n10544), .O(n10118) );
  NAND_GATE U10785 ( .I1(n10546), .I2(n10118), .O(n10121) );
  NAND3_GATE U10786 ( .I1(n10120), .I2(n10119), .I3(n736), .O(n10547) );
  NAND_GATE U10787 ( .I1(n10121), .I2(n10547), .O(n10556) );
  NAND_GATE U10788 ( .I1(n10557), .I2(n10556), .O(n10430) );
  NAND_GATE U10789 ( .I1(B[10]), .I2(A[25]), .O(n10578) );
  INV_GATE U10790 ( .I1(n10578), .O(n10427) );
  NAND3_GATE U10791 ( .I1(n10122), .I2(n10124), .I3(n10123), .O(n10407) );
  NAND3_GATE U10792 ( .I1(n10122), .I2(n10125), .I3(n825), .O(n10406) );
  AND_GATE U10793 ( .I1(n10407), .I2(n10406), .O(n10127) );
  NAND3_GATE U10794 ( .I1(n10124), .I2(n10123), .I3(n10404), .O(n10409) );
  NAND_GATE U10795 ( .I1(n10125), .I2(n825), .O(n10403) );
  NAND3_GATE U10796 ( .I1(n10409), .I2(n10403), .I3(n10404), .O(n10126) );
  NAND_GATE U10797 ( .I1(B[10]), .I2(A[23]), .O(n10602) );
  INV_GATE U10798 ( .I1(n10602), .O(n10410) );
  NAND3_GATE U10799 ( .I1(n10127), .I2(n10126), .I3(n10410), .O(n10603) );
  OR_GATE U10800 ( .I1(n10128), .I2(n10133), .O(n10131) );
  OR_GATE U10801 ( .I1(n10132), .I2(n10129), .O(n10130) );
  AND_GATE U10802 ( .I1(n10131), .I2(n10130), .O(n10138) );
  NAND_GATE U10803 ( .I1(n955), .I2(n10132), .O(n10135) );
  NAND3_GATE U10804 ( .I1(n10136), .I2(n10135), .I3(n10134), .O(n10137) );
  NAND_GATE U10805 ( .I1(n10138), .I2(n10137), .O(n10914) );
  NAND_GATE U10806 ( .I1(B[10]), .I2(A[22]), .O(n11008) );
  INV_GATE U10807 ( .I1(n11008), .O(n10911) );
  NAND_GATE U10808 ( .I1(n244), .I2(n10911), .O(n10912) );
  NAND_GATE U10809 ( .I1(B[10]), .I2(A[21]), .O(n10621) );
  INV_GATE U10810 ( .I1(n10621), .O(n10399) );
  NAND_GATE U10811 ( .I1(B[10]), .I2(A[20]), .O(n10896) );
  INV_GATE U10812 ( .I1(n10896), .O(n10895) );
  NAND_GATE U10813 ( .I1(n743), .I2(n10146), .O(n10144) );
  NAND3_GATE U10814 ( .I1(n10141), .I2(n10140), .I3(n10139), .O(n10143) );
  NAND3_GATE U10815 ( .I1(n10144), .I2(n10143), .I3(n10142), .O(n10150) );
  OR_GATE U10816 ( .I1(n10145), .I2(n10146), .O(n10149) );
  NAND3_GATE U10817 ( .I1(n10147), .I2(n743), .I3(n10146), .O(n10148) );
  NAND3_GATE U10818 ( .I1(n10150), .I2(n10149), .I3(n10148), .O(n10897) );
  NAND_GATE U10819 ( .I1(n10895), .I2(n603), .O(n10901) );
  NAND_GATE U10820 ( .I1(B[10]), .I2(A[19]), .O(n10632) );
  INV_GATE U10821 ( .I1(n10632), .O(n10388) );
  NAND3_GATE U10822 ( .I1(n10151), .I2(n576), .I3(n10154), .O(n10152) );
  AND_GATE U10823 ( .I1(n10153), .I2(n10152), .O(n10160) );
  NAND_GATE U10824 ( .I1(n10154), .I2(n576), .O(n10157) );
  NAND_GATE U10825 ( .I1(n565), .I2(n10155), .O(n10156) );
  NAND3_GATE U10826 ( .I1(n10158), .I2(n10157), .I3(n10156), .O(n10159) );
  NAND_GATE U10827 ( .I1(B[10]), .I2(A[18]), .O(n10885) );
  INV_GATE U10828 ( .I1(n10885), .O(n10879) );
  NAND_GATE U10829 ( .I1(n505), .I2(n10879), .O(n10876) );
  NAND_GATE U10830 ( .I1(B[10]), .I2(A[17]), .O(n10649) );
  INV_GATE U10831 ( .I1(n10649), .O(n10375) );
  NAND_GATE U10832 ( .I1(n1328), .I2(n10165), .O(n10162) );
  NAND_GATE U10833 ( .I1(n10163), .I2(n567), .O(n10161) );
  NAND_GATE U10834 ( .I1(n10162), .I2(n10161), .O(n10652) );
  NAND3_GATE U10835 ( .I1(n10375), .I2(n10646), .I3(n10647), .O(n10656) );
  NAND_GATE U10836 ( .I1(B[10]), .I2(A[16]), .O(n11060) );
  INV_GATE U10837 ( .I1(n11060), .O(n10869) );
  INV_GATE U10838 ( .I1(n10167), .O(n10169) );
  INV_GATE U10839 ( .I1(n10166), .O(n10171) );
  NAND_GATE U10840 ( .I1(n10171), .I2(n10167), .O(n10174) );
  NAND3_GATE U10841 ( .I1(n10173), .I2(n10174), .I3(n10175), .O(n10172) );
  NAND_GATE U10842 ( .I1(n164), .I2(n10169), .O(n10177) );
  NAND3_GATE U10843 ( .I1(n10172), .I2(n10177), .I3(n10176), .O(n10867) );
  NAND_GATE U10844 ( .I1(n10869), .I2(n566), .O(n10374) );
  NAND4_GATE U10845 ( .I1(n10175), .I2(n11060), .I3(n10174), .I4(n10173), .O(
        n10372) );
  NAND_GATE U10846 ( .I1(B[10]), .I2(A[15]), .O(n10661) );
  INV_GATE U10847 ( .I1(n10661), .O(n10369) );
  NAND_GATE U10848 ( .I1(n10182), .I2(n10178), .O(n10179) );
  NAND_GATE U10849 ( .I1(n10180), .I2(n10179), .O(n10185) );
  NAND_GATE U10850 ( .I1(n10181), .I2(n857), .O(n10182) );
  NAND_GATE U10851 ( .I1(n10183), .I2(n10182), .O(n10184) );
  NAND_GATE U10852 ( .I1(n10185), .I2(n10184), .O(n10190) );
  INV_GATE U10853 ( .I1(n10186), .O(n10188) );
  NAND_GATE U10854 ( .I1(n10188), .I2(n10187), .O(n10189) );
  NAND_GATE U10855 ( .I1(n10190), .I2(n10189), .O(n10664) );
  NAND_GATE U10856 ( .I1(n10369), .I2(n10664), .O(n10666) );
  INV_GATE U10857 ( .I1(n10191), .O(n10192) );
  NAND_GATE U10858 ( .I1(n10194), .I2(n10192), .O(n10202) );
  NAND_GATE U10859 ( .I1(n10194), .I2(n10199), .O(n10196) );
  NAND3_GATE U10860 ( .I1(n10197), .I2(n10196), .I3(n10195), .O(n10201) );
  OR_GATE U10861 ( .I1(n10199), .I2(n10198), .O(n10200) );
  NAND3_GATE U10862 ( .I1(n10202), .I2(n10201), .I3(n10200), .O(n10674) );
  INV_GATE U10863 ( .I1(n10674), .O(n10676) );
  NAND_GATE U10864 ( .I1(B[10]), .I2(A[14]), .O(n10680) );
  INV_GATE U10865 ( .I1(n10680), .O(n10672) );
  NAND_GATE U10866 ( .I1(n10676), .I2(n10672), .O(n10671) );
  NAND_GATE U10867 ( .I1(B[10]), .I2(A[13]), .O(n10689) );
  INV_GATE U10868 ( .I1(n10689), .O(n10365) );
  OR_GATE U10869 ( .I1(n10203), .I2(n10208), .O(n10206) );
  OR_GATE U10870 ( .I1(n10207), .I2(n10204), .O(n10205) );
  NAND_GATE U10871 ( .I1(n969), .I2(n10207), .O(n10211) );
  NAND3_GATE U10872 ( .I1(n10211), .I2(n10210), .I3(n10209), .O(n10212) );
  NAND_GATE U10873 ( .I1(B[10]), .I2(A[12]), .O(n10852) );
  NAND_GATE U10874 ( .I1(n100), .I2(n695), .O(n10846) );
  NAND_GATE U10875 ( .I1(B[10]), .I2(A[11]), .O(n10700) );
  INV_GATE U10876 ( .I1(n10700), .O(n10349) );
  INV_GATE U10877 ( .I1(n10213), .O(n10214) );
  NAND_GATE U10878 ( .I1(n10214), .I2(n10218), .O(n10224) );
  INV_GATE U10879 ( .I1(n10218), .O(n10215) );
  NAND_GATE U10880 ( .I1(n10216), .I2(n10215), .O(n10219) );
  NAND_GATE U10881 ( .I1(n10217), .I2(n10219), .O(n10222) );
  NAND_GATE U10882 ( .I1(n10222), .I2(n10221), .O(n10223) );
  NAND_GATE U10883 ( .I1(n10224), .I2(n10223), .O(n10698) );
  NAND_GATE U10884 ( .I1(B[10]), .I2(A[10]), .O(n10713) );
  INV_GATE U10885 ( .I1(n10713), .O(n10707) );
  INV_GATE U10886 ( .I1(n10225), .O(n10226) );
  NAND_GATE U10887 ( .I1(n10226), .I2(n10230), .O(n10237) );
  INV_GATE U10888 ( .I1(n10230), .O(n10227) );
  NAND_GATE U10889 ( .I1(n10228), .I2(n10227), .O(n10232) );
  NAND_GATE U10890 ( .I1(n10229), .I2(n10232), .O(n10235) );
  NAND_GATE U10891 ( .I1(n10235), .I2(n10234), .O(n10236) );
  NAND_GATE U10892 ( .I1(n10237), .I2(n10236), .O(n10722) );
  OR_GATE U10893 ( .I1(n10238), .I2(n10243), .O(n10241) );
  OR_GATE U10894 ( .I1(n10239), .I2(n10242), .O(n10240) );
  AND_GATE U10895 ( .I1(n10241), .I2(n10240), .O(n10248) );
  NAND_GATE U10896 ( .I1(n10242), .I2(n997), .O(n10246) );
  NAND3_GATE U10897 ( .I1(n10246), .I2(n10245), .I3(n10244), .O(n10247) );
  NAND_GATE U10898 ( .I1(n10248), .I2(n10247), .O(n10731) );
  INV_GATE U10899 ( .I1(n10731), .O(n10734) );
  INV_GATE U10900 ( .I1(n10249), .O(n10250) );
  NAND_GATE U10901 ( .I1(n10255), .I2(n10250), .O(n10263) );
  INV_GATE U10902 ( .I1(n10255), .O(n10252) );
  NAND_GATE U10903 ( .I1(n10252), .I2(n10251), .O(n10257) );
  NAND_GATE U10904 ( .I1(n10253), .I2(n10257), .O(n10261) );
  NAND_GATE U10905 ( .I1(n10255), .I2(n10254), .O(n10256) );
  NAND_GATE U10906 ( .I1(n10257), .I2(n10256), .O(n10258) );
  NAND_GATE U10907 ( .I1(n10259), .I2(n10258), .O(n10260) );
  NAND_GATE U10908 ( .I1(n10261), .I2(n10260), .O(n10262) );
  NAND_GATE U10909 ( .I1(n10263), .I2(n10262), .O(n10747) );
  OR_GATE U10910 ( .I1(n10264), .I2(n10269), .O(n10267) );
  OR_GATE U10911 ( .I1(n10265), .I2(n10268), .O(n10266) );
  AND_GATE U10912 ( .I1(n10267), .I2(n10266), .O(n10274) );
  NAND_GATE U10913 ( .I1(n10268), .I2(n1103), .O(n10272) );
  NAND3_GATE U10914 ( .I1(n10272), .I2(n10271), .I3(n10270), .O(n10273) );
  NAND_GATE U10915 ( .I1(n10274), .I2(n10273), .O(n10756) );
  INV_GATE U10916 ( .I1(n10756), .O(n10759) );
  INV_GATE U10917 ( .I1(n10275), .O(n10276) );
  NAND_GATE U10918 ( .I1(n10281), .I2(n10276), .O(n10289) );
  INV_GATE U10919 ( .I1(n10281), .O(n10278) );
  NAND_GATE U10920 ( .I1(n10278), .I2(n10277), .O(n10283) );
  NAND_GATE U10921 ( .I1(n10279), .I2(n10283), .O(n10287) );
  NAND_GATE U10922 ( .I1(n10281), .I2(n10280), .O(n10282) );
  NAND_GATE U10923 ( .I1(n10283), .I2(n10282), .O(n10284) );
  NAND_GATE U10924 ( .I1(n10285), .I2(n10284), .O(n10286) );
  NAND_GATE U10925 ( .I1(n10287), .I2(n10286), .O(n10288) );
  NAND_GATE U10926 ( .I1(n10289), .I2(n10288), .O(n10772) );
  OR_GATE U10927 ( .I1(n10290), .I2(n10295), .O(n10293) );
  OR_GATE U10928 ( .I1(n10291), .I2(n10294), .O(n10292) );
  AND_GATE U10929 ( .I1(n10293), .I2(n10292), .O(n10300) );
  NAND_GATE U10930 ( .I1(n10294), .I2(n1171), .O(n10298) );
  NAND3_GATE U10931 ( .I1(n10298), .I2(n10297), .I3(n10296), .O(n10299) );
  NAND_GATE U10932 ( .I1(n10300), .I2(n10299), .O(n10781) );
  INV_GATE U10933 ( .I1(n10781), .O(n10784) );
  OR_GATE U10934 ( .I1(n10301), .I2(n10303), .O(n10314) );
  NAND_GATE U10935 ( .I1(n10303), .I2(n10302), .O(n10308) );
  NAND_GATE U10936 ( .I1(n10304), .I2(n10308), .O(n10312) );
  NAND_GATE U10937 ( .I1(n10306), .I2(n10305), .O(n10307) );
  NAND_GATE U10938 ( .I1(n10308), .I2(n10307), .O(n10309) );
  NAND_GATE U10939 ( .I1(n10310), .I2(n10309), .O(n10311) );
  NAND_GATE U10940 ( .I1(n10312), .I2(n10311), .O(n10313) );
  NAND_GATE U10941 ( .I1(n10314), .I2(n10313), .O(n10797) );
  NAND3_GATE U10942 ( .I1(B[10]), .I2(B[11]), .I3(n1196), .O(n10806) );
  INV_GATE U10943 ( .I1(n10806), .O(n10809) );
  NAND_GATE U10944 ( .I1(n1375), .I2(A[0]), .O(n10315) );
  NAND_GATE U10945 ( .I1(n14781), .I2(n10315), .O(n10316) );
  NAND_GATE U10946 ( .I1(B[12]), .I2(n10316), .O(n10320) );
  NAND_GATE U10947 ( .I1(n1376), .I2(A[1]), .O(n10317) );
  NAND_GATE U10948 ( .I1(n14784), .I2(n10317), .O(n10318) );
  NAND_GATE U10949 ( .I1(B[11]), .I2(n10318), .O(n10319) );
  NAND_GATE U10950 ( .I1(n10320), .I2(n10319), .O(n10808) );
  INV_GATE U10951 ( .I1(n10808), .O(n10805) );
  NAND_GATE U10952 ( .I1(B[10]), .I2(A[2]), .O(n10813) );
  NAND_GATE U10953 ( .I1(n10805), .I2(n10813), .O(n10321) );
  NAND_GATE U10954 ( .I1(n10809), .I2(n10321), .O(n10322) );
  INV_GATE U10955 ( .I1(n10813), .O(n10807) );
  NAND_GATE U10956 ( .I1(n10808), .I2(n10807), .O(n10804) );
  NAND_GATE U10957 ( .I1(n10322), .I2(n10804), .O(n10798) );
  NAND_GATE U10958 ( .I1(n10797), .I2(n10798), .O(n10324) );
  NAND_GATE U10959 ( .I1(B[10]), .I2(A[3]), .O(n10799) );
  INV_GATE U10960 ( .I1(n10799), .O(n10323) );
  NAND_GATE U10961 ( .I1(n10797), .I2(n10323), .O(n10794) );
  NAND_GATE U10962 ( .I1(n10798), .I2(n10323), .O(n10793) );
  NAND3_GATE U10963 ( .I1(n10324), .I2(n10794), .I3(n10793), .O(n10783) );
  INV_GATE U10964 ( .I1(n10783), .O(n10780) );
  NAND_GATE U10965 ( .I1(B[10]), .I2(A[4]), .O(n10788) );
  NAND_GATE U10966 ( .I1(n10780), .I2(n10788), .O(n10325) );
  NAND_GATE U10967 ( .I1(n10784), .I2(n10325), .O(n10326) );
  INV_GATE U10968 ( .I1(n10788), .O(n10782) );
  NAND_GATE U10969 ( .I1(n10783), .I2(n10782), .O(n10779) );
  NAND_GATE U10970 ( .I1(n10326), .I2(n10779), .O(n10773) );
  NAND_GATE U10971 ( .I1(n10772), .I2(n10773), .O(n10328) );
  NAND_GATE U10972 ( .I1(B[10]), .I2(A[5]), .O(n10774) );
  INV_GATE U10973 ( .I1(n10774), .O(n10327) );
  NAND_GATE U10974 ( .I1(n10772), .I2(n10327), .O(n10769) );
  NAND_GATE U10975 ( .I1(n10773), .I2(n10327), .O(n10768) );
  NAND3_GATE U10976 ( .I1(n10328), .I2(n10769), .I3(n10768), .O(n10758) );
  INV_GATE U10977 ( .I1(n10758), .O(n10755) );
  NAND_GATE U10978 ( .I1(B[10]), .I2(A[6]), .O(n10763) );
  NAND_GATE U10979 ( .I1(n10755), .I2(n10763), .O(n10329) );
  NAND_GATE U10980 ( .I1(n10759), .I2(n10329), .O(n10330) );
  INV_GATE U10981 ( .I1(n10763), .O(n10757) );
  NAND_GATE U10982 ( .I1(n10758), .I2(n10757), .O(n10754) );
  NAND_GATE U10983 ( .I1(n10330), .I2(n10754), .O(n10748) );
  NAND_GATE U10984 ( .I1(n10747), .I2(n10748), .O(n10332) );
  NAND_GATE U10985 ( .I1(B[10]), .I2(A[7]), .O(n10749) );
  INV_GATE U10986 ( .I1(n10749), .O(n10331) );
  NAND_GATE U10987 ( .I1(n10747), .I2(n10331), .O(n10744) );
  NAND_GATE U10988 ( .I1(n10748), .I2(n10331), .O(n10743) );
  NAND3_GATE U10989 ( .I1(n10332), .I2(n10744), .I3(n10743), .O(n10733) );
  INV_GATE U10990 ( .I1(n10733), .O(n10730) );
  NAND_GATE U10991 ( .I1(B[10]), .I2(A[8]), .O(n10738) );
  NAND_GATE U10992 ( .I1(n10730), .I2(n10738), .O(n10333) );
  NAND_GATE U10993 ( .I1(n10734), .I2(n10333), .O(n10334) );
  INV_GATE U10994 ( .I1(n10738), .O(n10732) );
  NAND_GATE U10995 ( .I1(n10733), .I2(n10732), .O(n10729) );
  NAND_GATE U10996 ( .I1(n10334), .I2(n10729), .O(n10723) );
  NAND_GATE U10997 ( .I1(n10722), .I2(n10723), .O(n10336) );
  NAND_GATE U10998 ( .I1(B[10]), .I2(A[9]), .O(n10724) );
  INV_GATE U10999 ( .I1(n10724), .O(n10335) );
  NAND_GATE U11000 ( .I1(n10722), .I2(n10335), .O(n10719) );
  NAND_GATE U11001 ( .I1(n10723), .I2(n10335), .O(n10718) );
  NAND3_GATE U11002 ( .I1(n10336), .I2(n10719), .I3(n10718), .O(n10709) );
  NAND_GATE U11003 ( .I1(n10707), .I2(n10709), .O(n10704) );
  OR_GATE U11004 ( .I1(n10337), .I2(n10342), .O(n10340) );
  OR_GATE U11005 ( .I1(n10341), .I2(n10338), .O(n10339) );
  NAND_GATE U11006 ( .I1(n945), .I2(n10341), .O(n10345) );
  NAND3_GATE U11007 ( .I1(n10345), .I2(n10344), .I3(n10343), .O(n10346) );
  INV_GATE U11008 ( .I1(n10705), .O(n10708) );
  INV_GATE U11009 ( .I1(n10709), .O(n10706) );
  NAND_GATE U11010 ( .I1(n10713), .I2(n10706), .O(n10347) );
  NAND_GATE U11011 ( .I1(n10708), .I2(n10347), .O(n10348) );
  NAND_GATE U11012 ( .I1(n10704), .I2(n10348), .O(n10699) );
  NAND_GATE U11013 ( .I1(n10698), .I2(n10699), .O(n10350) );
  NAND_GATE U11014 ( .I1(n10349), .I2(n10699), .O(n10694) );
  NAND3_GATE U11015 ( .I1(n10695), .I2(n10350), .I3(n10694), .O(n10850) );
  NAND_GATE U11016 ( .I1(n10849), .I2(n10852), .O(n10351) );
  NAND_GATE U11017 ( .I1(n10850), .I2(n10351), .O(n10352) );
  NAND_GATE U11018 ( .I1(n10846), .I2(n10352), .O(n10688) );
  NAND_GATE U11019 ( .I1(n10365), .I2(n10688), .O(n10684) );
  OR_GATE U11020 ( .I1(n10354), .I2(n10353), .O(n10364) );
  NAND_GATE U11021 ( .I1(n860), .I2(n10354), .O(n10358) );
  NAND_GATE U11022 ( .I1(n10355), .I2(n10358), .O(n10362) );
  NAND_GATE U11023 ( .I1(n10358), .I2(n10357), .O(n10359) );
  NAND_GATE U11024 ( .I1(n10360), .I2(n10359), .O(n10361) );
  NAND_GATE U11025 ( .I1(n10362), .I2(n10361), .O(n10363) );
  NAND_GATE U11026 ( .I1(n10364), .I2(n10363), .O(n10687) );
  NAND_GATE U11027 ( .I1(n10688), .I2(n10687), .O(n10366) );
  NAND3_GATE U11028 ( .I1(n10684), .I2(n10366), .I3(n10683), .O(n10675) );
  NAND_GATE U11029 ( .I1(n10674), .I2(n10680), .O(n10367) );
  NAND_GATE U11030 ( .I1(n10675), .I2(n10367), .O(n10368) );
  NAND_GATE U11031 ( .I1(n10664), .I2(n10667), .O(n10370) );
  NAND3_GATE U11032 ( .I1(n10666), .I2(n10370), .I3(n10665), .O(n10870) );
  NAND3_GATE U11033 ( .I1(n10372), .I2(n10371), .I3(n10870), .O(n10373) );
  NAND_GATE U11034 ( .I1(n10374), .I2(n10373), .O(n10657) );
  NAND3_GATE U11035 ( .I1(n10646), .I2(n10647), .I3(n10657), .O(n10376) );
  NAND_GATE U11036 ( .I1(n10375), .I2(n10657), .O(n10655) );
  NAND3_GATE U11037 ( .I1(n10656), .I2(n10376), .I3(n10655), .O(n10882) );
  NAND_GATE U11038 ( .I1(n10881), .I2(n10885), .O(n10377) );
  NAND_GATE U11039 ( .I1(n10882), .I2(n10377), .O(n10378) );
  NAND_GATE U11040 ( .I1(n10876), .I2(n10378), .O(n10641) );
  NAND_GATE U11041 ( .I1(n10388), .I2(n10641), .O(n10637) );
  INV_GATE U11042 ( .I1(n10383), .O(n10379) );
  NAND_GATE U11043 ( .I1(n10380), .I2(n10379), .O(n10385) );
  NAND_GATE U11044 ( .I1(n10381), .I2(n10385), .O(n10636) );
  NAND_GATE U11045 ( .I1(n741), .I2(n10383), .O(n10384) );
  NAND_GATE U11046 ( .I1(n10385), .I2(n10384), .O(n10386) );
  NAND_GATE U11047 ( .I1(n10387), .I2(n10386), .O(n10635) );
  NAND3_GATE U11048 ( .I1(n10641), .I2(n10631), .I3(n10635), .O(n10389) );
  NAND3_GATE U11049 ( .I1(n10388), .I2(n10631), .I3(n10635), .O(n10642) );
  NAND_GATE U11050 ( .I1(n10896), .I2(n10897), .O(n10390) );
  NAND_GATE U11051 ( .I1(n10902), .I2(n10390), .O(n10619) );
  NAND_GATE U11052 ( .I1(n10901), .I2(n10619), .O(n10617) );
  NAND_GATE U11053 ( .I1(n10399), .I2(n10617), .O(n10624) );
  NAND_GATE U11054 ( .I1(n10392), .I2(n10397), .O(n10611) );
  NAND_GATE U11055 ( .I1(n10394), .I2(n10393), .O(n10397) );
  NAND_GATE U11056 ( .I1(n670), .I2(n10395), .O(n10396) );
  NAND_GATE U11057 ( .I1(n10397), .I2(n10396), .O(n10614) );
  NAND_GATE U11058 ( .I1(n10611), .I2(n10618), .O(n10398) );
  NAND_GATE U11059 ( .I1(n10613), .I2(n10398), .O(n10625) );
  NAND_GATE U11060 ( .I1(n10617), .I2(n10625), .O(n10400) );
  NAND_GATE U11061 ( .I1(n10399), .I2(n10625), .O(n10610) );
  NAND_GATE U11062 ( .I1(n10914), .I2(n11008), .O(n10401) );
  NAND_GATE U11063 ( .I1(n669), .I2(n10401), .O(n10402) );
  NAND_GATE U11064 ( .I1(n10912), .I2(n10402), .O(n10604) );
  NAND_GATE U11065 ( .I1(n10404), .I2(n10403), .O(n10405) );
  NAND3_GATE U11066 ( .I1(n10407), .I2(n10406), .I3(n10405), .O(n10408) );
  NAND_GATE U11067 ( .I1(n10409), .I2(n10408), .O(n10605) );
  NAND_GATE U11068 ( .I1(n10604), .I2(n10605), .O(n10411) );
  NAND_GATE U11069 ( .I1(n10410), .I2(n10604), .O(n10606) );
  NAND3_GATE U11070 ( .I1(n10603), .I2(n10411), .I3(n10606), .O(n10588) );
  NAND_GATE U11071 ( .I1(n806), .I2(n10416), .O(n10412) );
  NAND_GATE U11072 ( .I1(n10414), .I2(n10412), .O(n10592) );
  NAND_GATE U11073 ( .I1(n10593), .I2(n10592), .O(n10417) );
  NAND_GATE U11074 ( .I1(n10415), .I2(n10414), .O(n10594) );
  NAND3_GATE U11075 ( .I1(n10416), .I2(n10415), .I3(n806), .O(n10598) );
  NAND3_GATE U11076 ( .I1(n10588), .I2(n10417), .I3(n10583), .O(n10419) );
  NAND_GATE U11077 ( .I1(B[10]), .I2(A[24]), .O(n10585) );
  INV_GATE U11078 ( .I1(n10585), .O(n10418) );
  NAND3_GATE U11079 ( .I1(n10418), .I2(n10417), .I3(n10583), .O(n10589) );
  NAND_GATE U11080 ( .I1(n10418), .I2(n10588), .O(n10595) );
  NAND3_GATE U11081 ( .I1(n10419), .I2(n10589), .I3(n10595), .O(n10575) );
  NAND_GATE U11082 ( .I1(n10427), .I2(n10575), .O(n10564) );
  NAND_GATE U11083 ( .I1(n10420), .I2(n10425), .O(n10563) );
  INV_GATE U11084 ( .I1(n10563), .O(n10570) );
  NAND_GATE U11085 ( .I1(n10423), .I2(n10422), .O(n10426) );
  NAND_GATE U11086 ( .I1(n10424), .I2(n15), .O(n10425) );
  NAND_GATE U11087 ( .I1(n10426), .I2(n10425), .O(n10567) );
  NAND3_GATE U11088 ( .I1(n10575), .I2(n10573), .I3(n10572), .O(n10428) );
  NAND3_GATE U11089 ( .I1(n10427), .I2(n10573), .I3(n10572), .O(n10562) );
  NAND3_GATE U11090 ( .I1(n10564), .I2(n10428), .I3(n10562), .O(n10550) );
  NAND_GATE U11091 ( .I1(n10556), .I2(n10550), .O(n10429) );
  NAND_GATE U11092 ( .I1(n10557), .I2(n10550), .O(n10555) );
  NAND3_GATE U11093 ( .I1(n10430), .I2(n10429), .I3(n10555), .O(n10532) );
  NAND_GATE U11094 ( .I1(n10538), .I2(n10532), .O(n10539) );
  NAND3_GATE U11095 ( .I1(n10432), .I2(n10433), .I3(n10434), .O(n10528) );
  NAND_GATE U11096 ( .I1(n10435), .I2(n569), .O(n10431) );
  NAND_GATE U11097 ( .I1(n10432), .I2(n10431), .O(n10527) );
  NAND_GATE U11098 ( .I1(n10434), .I2(n10433), .O(n10436) );
  NAND_GATE U11099 ( .I1(n10436), .I2(n10431), .O(n10529) );
  NAND_GATE U11100 ( .I1(n10527), .I2(n10533), .O(n10437) );
  NAND_GATE U11101 ( .I1(n10528), .I2(n10437), .O(n10540) );
  NAND_GATE U11102 ( .I1(n10538), .I2(n10540), .O(n10439) );
  NAND_GATE U11103 ( .I1(n10532), .I2(n10540), .O(n10438) );
  NAND3_GATE U11104 ( .I1(n10539), .I2(n10439), .I3(n10438), .O(n10938) );
  NAND_GATE U11105 ( .I1(n10947), .I2(n10938), .O(n10944) );
  NAND3_GATE U11106 ( .I1(n10441), .I2(n10442), .I3(n10443), .O(n10934) );
  INV_GATE U11107 ( .I1(n10442), .O(n10444) );
  NAND_GATE U11108 ( .I1(n10445), .I2(n10444), .O(n10440) );
  NAND_GATE U11109 ( .I1(n10441), .I2(n10440), .O(n10933) );
  NAND_GATE U11110 ( .I1(n10443), .I2(n10442), .O(n10446) );
  NAND_GATE U11111 ( .I1(n10446), .I2(n10440), .O(n10935) );
  NAND_GATE U11112 ( .I1(n10933), .I2(n10939), .O(n10447) );
  NAND_GATE U11113 ( .I1(n10934), .I2(n10447), .O(n10945) );
  NAND_GATE U11114 ( .I1(n10947), .I2(n10945), .O(n10449) );
  NAND_GATE U11115 ( .I1(n10938), .I2(n10945), .O(n10448) );
  NAND3_GATE U11116 ( .I1(n10944), .I2(n10449), .I3(n10448), .O(n10523) );
  NAND_GATE U11117 ( .I1(n10461), .I2(n10523), .O(n10521) );
  INV_GATE U11118 ( .I1(n10453), .O(n10455) );
  NAND_GATE U11119 ( .I1(n10456), .I2(n10455), .O(n10451) );
  NAND_GATE U11120 ( .I1(n10452), .I2(n10451), .O(n10458) );
  NAND_GATE U11121 ( .I1(n10460), .I2(n10459), .O(n10524) );
  NAND_GATE U11122 ( .I1(n10461), .I2(n10524), .O(n10522) );
  NAND_GATE U11123 ( .I1(n10523), .I2(n10524), .O(n10462) );
  NAND3_GATE U11124 ( .I1(n10521), .I2(n10522), .I3(n10462), .O(n10510) );
  NAND_GATE U11125 ( .I1(n10515), .I2(n10510), .O(n10516) );
  NAND_GATE U11126 ( .I1(n10465), .I2(n10464), .O(n10466) );
  NAND_GATE U11127 ( .I1(n10467), .I2(n10466), .O(n10505) );
  NAND_GATE U11128 ( .I1(n10504), .I2(n10468), .O(n10517) );
  NAND_GATE U11129 ( .I1(n10515), .I2(n10517), .O(n10470) );
  NAND_GATE U11130 ( .I1(n10510), .I2(n10517), .O(n10469) );
  NAND3_GATE U11131 ( .I1(n10516), .I2(n10470), .I3(n10469), .O(n10961) );
  NAND_GATE U11132 ( .I1(n10485), .I2(n10961), .O(n10959) );
  INV_GATE U11133 ( .I1(n10471), .O(n10472) );
  NAND_GATE U11134 ( .I1(n10472), .I2(n10475), .O(n10484) );
  NAND_GATE U11135 ( .I1(n10477), .I2(n1242), .O(n10473) );
  NAND_GATE U11136 ( .I1(n10474), .I2(n10473), .O(n10482) );
  NAND_GATE U11137 ( .I1(n10478), .I2(n10473), .O(n10479) );
  NAND_GATE U11138 ( .I1(n10480), .I2(n10479), .O(n10481) );
  NAND_GATE U11139 ( .I1(n10482), .I2(n10481), .O(n10483) );
  NAND_GATE U11140 ( .I1(n10484), .I2(n10483), .O(n10960) );
  NAND_GATE U11141 ( .I1(n10485), .I2(n10960), .O(n10962) );
  NAND_GATE U11142 ( .I1(n10961), .I2(n10960), .O(n10486) );
  NAND3_GATE U11143 ( .I1(n10959), .I2(n10962), .I3(n10486), .O(n15340) );
  NAND_GATE U11144 ( .I1(n10487), .I2(n10493), .O(n10489) );
  NAND_GATE U11145 ( .I1(n10490), .I2(n821), .O(n10488) );
  NAND_GATE U11146 ( .I1(n10489), .I2(n10488), .O(n15335) );
  NAND_GATE U11147 ( .I1(n10491), .I2(n10488), .O(n15337) );
  NAND_GATE U11148 ( .I1(n10495), .I2(n10496), .O(n10494) );
  OR_GATE U11149 ( .I1(n15340), .I2(n10494), .O(n10499) );
  NAND_GATE U11150 ( .I1(n10496), .I2(n10495), .O(n10497) );
  NAND_GATE U11151 ( .I1(n15340), .I2(n10497), .O(n10498) );
  NAND_GATE U11152 ( .I1(n10499), .I2(n10498), .O(\A1[40] ) );
  NAND_GATE U11153 ( .I1(n10961), .I2(n275), .O(n10502) );
  INV_GATE U11154 ( .I1(n10961), .O(n10500) );
  NAND_GATE U11155 ( .I1(n10500), .I2(n10960), .O(n10501) );
  NAND3_GATE U11156 ( .I1(n10503), .I2(n10502), .I3(n10501), .O(n10965) );
  NAND_GATE U11157 ( .I1(B[9]), .I2(A[31]), .O(n15343) );
  INV_GATE U11158 ( .I1(n15343), .O(n10973) );
  NAND_GATE U11159 ( .I1(n10504), .I2(n1252), .O(n10508) );
  NAND_GATE U11160 ( .I1(n10506), .I2(n10505), .O(n10507) );
  NAND3_GATE U11161 ( .I1(n10508), .I2(n10514), .I3(n10507), .O(n10512) );
  NAND_GATE U11162 ( .I1(n10508), .I2(n10507), .O(n10509) );
  NAND_GATE U11163 ( .I1(n10510), .I2(n10509), .O(n10511) );
  NAND3_GATE U11164 ( .I1(n10513), .I2(n10512), .I3(n10511), .O(n10520) );
  NAND3_GATE U11165 ( .I1(n10515), .I2(n10514), .I3(n10517), .O(n10519) );
  OR_GATE U11166 ( .I1(n10517), .I2(n10516), .O(n10518) );
  NAND3_GATE U11167 ( .I1(n10520), .I2(n10519), .I3(n10518), .O(n10971) );
  INV_GATE U11168 ( .I1(n10971), .O(n10974) );
  NAND_GATE U11169 ( .I1(n10973), .I2(n10974), .O(n10958) );
  INV_GATE U11170 ( .I1(n10523), .O(n10525) );
  NAND_GATE U11171 ( .I1(n10525), .I2(n10524), .O(n10979) );
  NAND3_GATE U11172 ( .I1(n10981), .I2(n10980), .I3(n10979), .O(n10526) );
  NAND3_GATE U11173 ( .I1(n10977), .I2(n10976), .I3(n10526), .O(n10982) );
  NAND_GATE U11174 ( .I1(B[9]), .I2(A[30]), .O(n10983) );
  NAND_GATE U11175 ( .I1(B[9]), .I2(A[28]), .O(n11417) );
  INV_GATE U11176 ( .I1(n11417), .O(n11355) );
  NAND_GATE U11177 ( .I1(n10530), .I2(n10529), .O(n10533) );
  NAND_GATE U11178 ( .I1(n10534), .I2(n10533), .O(n10531) );
  NAND_GATE U11179 ( .I1(n10532), .I2(n10531), .O(n10537) );
  NAND3_GATE U11180 ( .I1(n10534), .I2(n10533), .I3(n594), .O(n10536) );
  NAND3_GATE U11181 ( .I1(n10537), .I2(n10536), .I3(n10535), .O(n10543) );
  NAND3_GATE U11182 ( .I1(n10538), .I2(n594), .I3(n10540), .O(n10542) );
  OR_GATE U11183 ( .I1(n10540), .I2(n10539), .O(n10541) );
  NAND3_GATE U11184 ( .I1(n10543), .I2(n10542), .I3(n10541), .O(n11415) );
  NAND_GATE U11185 ( .I1(n11355), .I2(n621), .O(n10932) );
  NAND_GATE U11186 ( .I1(B[9]), .I2(A[27]), .O(n11440) );
  INV_GATE U11187 ( .I1(n11440), .O(n10990) );
  INV_GATE U11188 ( .I1(n10546), .O(n10548) );
  NAND_GATE U11189 ( .I1(n10548), .I2(n10547), .O(n10551) );
  NAND_GATE U11190 ( .I1(n10118), .I2(n10551), .O(n10549) );
  NAND_GATE U11191 ( .I1(n10550), .I2(n10549), .O(n10553) );
  INV_GATE U11192 ( .I1(n10550), .O(n10558) );
  NAND3_GATE U11193 ( .I1(n10551), .I2(n10558), .I3(n10118), .O(n10552) );
  NAND3_GATE U11194 ( .I1(n10554), .I2(n10553), .I3(n10552), .O(n10561) );
  OR_GATE U11195 ( .I1(n10555), .I2(n10556), .O(n10560) );
  NAND3_GATE U11196 ( .I1(n10558), .I2(n10557), .I3(n10556), .O(n10559) );
  NAND3_GATE U11197 ( .I1(n10561), .I2(n10560), .I3(n10559), .O(n11436) );
  NAND_GATE U11198 ( .I1(n10990), .I2(n738), .O(n10929) );
  NAND_GATE U11199 ( .I1(B[9]), .I2(A[26]), .O(n11458) );
  INV_GATE U11200 ( .I1(n11458), .O(n10993) );
  OR_GATE U11201 ( .I1(n10562), .I2(n10575), .O(n10581) );
  NAND_GATE U11202 ( .I1(n10563), .I2(n10572), .O(n10566) );
  INV_GATE U11203 ( .I1(n10564), .O(n10565) );
  NAND3_GATE U11204 ( .I1(n10566), .I2(n10565), .I3(n10569), .O(n10580) );
  NAND_GATE U11205 ( .I1(n10568), .I2(n10567), .O(n10572) );
  INV_GATE U11206 ( .I1(n10575), .O(n10571) );
  NAND_GATE U11207 ( .I1(n10570), .I2(n10569), .O(n10573) );
  NAND3_GATE U11208 ( .I1(n10572), .I2(n10571), .I3(n10573), .O(n10577) );
  NAND_GATE U11209 ( .I1(n10573), .I2(n10572), .O(n10574) );
  NAND_GATE U11210 ( .I1(n10575), .I2(n10574), .O(n10576) );
  NAND3_GATE U11211 ( .I1(n10578), .I2(n10577), .I3(n10576), .O(n10579) );
  NAND3_GATE U11212 ( .I1(n10581), .I2(n10580), .I3(n10579), .O(n10995) );
  NAND_GATE U11213 ( .I1(n10993), .I2(n10997), .O(n10926) );
  NAND_GATE U11214 ( .I1(B[9]), .I2(A[25]), .O(n11825) );
  INV_GATE U11215 ( .I1(n11825), .O(n11000) );
  NAND_GATE U11216 ( .I1(n10593), .I2(n10592), .O(n10582) );
  NAND_GATE U11217 ( .I1(n10583), .I2(n10582), .O(n10584) );
  NAND_GATE U11218 ( .I1(n10588), .I2(n10584), .O(n10587) );
  OR_GATE U11219 ( .I1(n10584), .I2(n10588), .O(n10586) );
  NAND3_GATE U11220 ( .I1(n10587), .I2(n10586), .I3(n10585), .O(n10591) );
  OR_GATE U11221 ( .I1(n10589), .I2(n10588), .O(n10590) );
  NAND_GATE U11222 ( .I1(n10594), .I2(n10417), .O(n10597) );
  INV_GATE U11223 ( .I1(n10595), .O(n10596) );
  NAND3_GATE U11224 ( .I1(n10598), .I2(n10597), .I3(n10596), .O(n10599) );
  INV_GATE U11225 ( .I1(n11003), .O(n11002) );
  NAND_GATE U11226 ( .I1(n11000), .I2(n11002), .O(n10923) );
  NAND_GATE U11227 ( .I1(B[9]), .I2(A[24]), .O(n11334) );
  INV_GATE U11228 ( .I1(n11334), .O(n11338) );
  NAND_GATE U11229 ( .I1(n242), .I2(n10605), .O(n10601) );
  NAND3_GATE U11230 ( .I1(n10602), .I2(n10601), .I3(n10600), .O(n10609) );
  OR_GATE U11231 ( .I1(n10604), .I2(n10603), .O(n10608) );
  OR_GATE U11232 ( .I1(n10606), .I2(n10605), .O(n10607) );
  NAND3_GATE U11233 ( .I1(n10609), .I2(n10608), .I3(n10607), .O(n11336) );
  NAND_GATE U11234 ( .I1(n11338), .I2(n243), .O(n11342) );
  NAND_GATE U11235 ( .I1(B[9]), .I2(A[23]), .O(n11019) );
  INV_GATE U11236 ( .I1(n11019), .O(n10915) );
  NAND_GATE U11237 ( .I1(B[9]), .I2(A[22]), .O(n11316) );
  INV_GATE U11238 ( .I1(n11316), .O(n11320) );
  OR_GATE U11239 ( .I1(n10610), .I2(n10617), .O(n10628) );
  INV_GATE U11240 ( .I1(n10611), .O(n10612) );
  NAND_GATE U11241 ( .I1(n10613), .I2(n10612), .O(n10620) );
  NAND_GATE U11242 ( .I1(n10615), .I2(n10614), .O(n10618) );
  NAND_GATE U11243 ( .I1(n10620), .I2(n10618), .O(n10616) );
  NAND_GATE U11244 ( .I1(n10617), .I2(n10616), .O(n10623) );
  NAND4_GATE U11245 ( .I1(n10620), .I2(n10619), .I3(n10901), .I4(n10618), .O(
        n10622) );
  NAND3_GATE U11246 ( .I1(n10623), .I2(n10622), .I3(n10621), .O(n10627) );
  OR_GATE U11247 ( .I1(n10625), .I2(n10624), .O(n10626) );
  NAND3_GATE U11248 ( .I1(n10628), .I2(n10627), .I3(n10626), .O(n11318) );
  INV_GATE U11249 ( .I1(n11318), .O(n11315) );
  NAND_GATE U11250 ( .I1(n11320), .I2(n11315), .O(n11324) );
  NAND_GATE U11251 ( .I1(B[9]), .I2(A[21]), .O(n11026) );
  INV_GATE U11252 ( .I1(n11026), .O(n10906) );
  NAND_GATE U11253 ( .I1(n10631), .I2(n10635), .O(n10629) );
  NAND_GATE U11254 ( .I1(n10641), .I2(n10629), .O(n10634) );
  INV_GATE U11255 ( .I1(n10641), .O(n10630) );
  NAND3_GATE U11256 ( .I1(n10631), .I2(n10635), .I3(n10630), .O(n10633) );
  NAND3_GATE U11257 ( .I1(n10634), .I2(n10633), .I3(n10632), .O(n10645) );
  NAND_GATE U11258 ( .I1(n10636), .I2(n10635), .O(n10639) );
  INV_GATE U11259 ( .I1(n10637), .O(n10638) );
  NAND3_GATE U11260 ( .I1(n10640), .I2(n10639), .I3(n10638), .O(n10644) );
  OR_GATE U11261 ( .I1(n10642), .I2(n10641), .O(n10643) );
  NAND3_GATE U11262 ( .I1(n10645), .I2(n10644), .I3(n10643), .O(n11307) );
  INV_GATE U11263 ( .I1(n11307), .O(n11304) );
  NAND_GATE U11264 ( .I1(B[9]), .I2(A[20]), .O(n11305) );
  INV_GATE U11265 ( .I1(n11305), .O(n11502) );
  NAND_GATE U11266 ( .I1(n11304), .I2(n11502), .O(n11308) );
  NAND_GATE U11267 ( .I1(B[9]), .I2(A[19]), .O(n11041) );
  INV_GATE U11268 ( .I1(n11041), .O(n11034) );
  NAND_GATE U11269 ( .I1(n10653), .I2(n10652), .O(n10646) );
  NAND_GATE U11270 ( .I1(n10647), .I2(n10646), .O(n10648) );
  OR_GATE U11271 ( .I1(n10648), .I2(n10657), .O(n10651) );
  NAND_GATE U11272 ( .I1(n10657), .I2(n10648), .O(n10650) );
  NAND3_GATE U11273 ( .I1(n10651), .I2(n10650), .I3(n10649), .O(n10660) );
  OR_GATE U11274 ( .I1(n10657), .I2(n10656), .O(n10658) );
  NAND3_GATE U11275 ( .I1(n10660), .I2(n10659), .I3(n10658), .O(n11048) );
  NAND_GATE U11276 ( .I1(B[9]), .I2(A[18]), .O(n11052) );
  INV_GATE U11277 ( .I1(n11052), .O(n11046) );
  NAND_GATE U11278 ( .I1(n1327), .I2(n11046), .O(n11055) );
  NAND_GATE U11279 ( .I1(B[9]), .I2(A[17]), .O(n11072) );
  INV_GATE U11280 ( .I1(n11072), .O(n10872) );
  NAND_GATE U11281 ( .I1(n10664), .I2(n170), .O(n10663) );
  NAND3_GATE U11282 ( .I1(n10663), .I2(n10662), .I3(n10661), .O(n10670) );
  OR_GATE U11283 ( .I1(n10665), .I2(n10664), .O(n10669) );
  OR_GATE U11284 ( .I1(n10667), .I2(n10666), .O(n10668) );
  NAND3_GATE U11285 ( .I1(n10670), .I2(n10669), .I3(n10668), .O(n11287) );
  INV_GATE U11286 ( .I1(n11287), .O(n11289) );
  NAND_GATE U11287 ( .I1(B[9]), .I2(A[16]), .O(n11291) );
  INV_GATE U11288 ( .I1(n11291), .O(n11285) );
  NAND_GATE U11289 ( .I1(n11289), .I2(n11285), .O(n11283) );
  NAND_GATE U11290 ( .I1(B[9]), .I2(A[15]), .O(n11087) );
  INV_GATE U11291 ( .I1(n11087), .O(n10861) );
  INV_GATE U11292 ( .I1(n10675), .O(n10673) );
  NAND_GATE U11293 ( .I1(n10672), .I2(n10678), .O(n10681) );
  NAND_GATE U11294 ( .I1(n10674), .I2(n10673), .O(n10678) );
  NAND_GATE U11295 ( .I1(n10676), .I2(n10675), .O(n10677) );
  NAND_GATE U11296 ( .I1(n10678), .I2(n10677), .O(n10679) );
  NAND_GATE U11297 ( .I1(n10861), .I2(n11081), .O(n11077) );
  NAND_GATE U11298 ( .I1(n10680), .I2(n10679), .O(n11083) );
  OR_GATE U11299 ( .I1(n10683), .I2(n10688), .O(n10686) );
  OR_GATE U11300 ( .I1(n10687), .I2(n10684), .O(n10685) );
  AND_GATE U11301 ( .I1(n10686), .I2(n10685), .O(n10693) );
  NAND_GATE U11302 ( .I1(n508), .I2(n10687), .O(n10691) );
  NAND3_GATE U11303 ( .I1(n10691), .I2(n10690), .I3(n10689), .O(n10692) );
  NAND_GATE U11304 ( .I1(n10693), .I2(n10692), .O(n11269) );
  INV_GATE U11305 ( .I1(n11269), .O(n11272) );
  NAND_GATE U11306 ( .I1(B[9]), .I2(A[14]), .O(n11274) );
  INV_GATE U11307 ( .I1(n11274), .O(n11270) );
  NAND_GATE U11308 ( .I1(n11272), .I2(n11270), .O(n11266) );
  NAND_GATE U11309 ( .I1(B[9]), .I2(A[13]), .O(n11097) );
  INV_GATE U11310 ( .I1(n11097), .O(n10857) );
  OR_GATE U11311 ( .I1(n10694), .I2(n10698), .O(n10697) );
  OR_GATE U11312 ( .I1(n10699), .I2(n10695), .O(n10696) );
  NAND_GATE U11313 ( .I1(n10698), .I2(n985), .O(n10702) );
  NAND3_GATE U11314 ( .I1(n10702), .I2(n10701), .I3(n10700), .O(n10703) );
  INV_GATE U11315 ( .I1(n11102), .O(n11105) );
  NAND_GATE U11316 ( .I1(B[9]), .I2(A[12]), .O(n11107) );
  INV_GATE U11317 ( .I1(n11107), .O(n11103) );
  NAND_GATE U11318 ( .I1(n11105), .I2(n11103), .O(n11101) );
  OR_GATE U11319 ( .I1(n10705), .I2(n10704), .O(n10717) );
  NAND_GATE U11320 ( .I1(n10706), .I2(n10705), .O(n10711) );
  NAND_GATE U11321 ( .I1(n10707), .I2(n10711), .O(n10715) );
  NAND_GATE U11322 ( .I1(n10709), .I2(n10708), .O(n10710) );
  NAND_GATE U11323 ( .I1(n10711), .I2(n10710), .O(n10712) );
  NAND_GATE U11324 ( .I1(n10713), .I2(n10712), .O(n10714) );
  NAND_GATE U11325 ( .I1(n10715), .I2(n10714), .O(n10716) );
  NAND_GATE U11326 ( .I1(n10717), .I2(n10716), .O(n11253) );
  OR_GATE U11327 ( .I1(n10718), .I2(n10722), .O(n10721) );
  OR_GATE U11328 ( .I1(n10719), .I2(n10723), .O(n10720) );
  AND_GATE U11329 ( .I1(n10721), .I2(n10720), .O(n10728) );
  NAND_GATE U11330 ( .I1(n10722), .I2(n975), .O(n10726) );
  NAND3_GATE U11331 ( .I1(n10726), .I2(n10725), .I3(n10724), .O(n10727) );
  NAND_GATE U11332 ( .I1(n10728), .I2(n10727), .O(n11114) );
  INV_GATE U11333 ( .I1(n11114), .O(n11117) );
  OR_GATE U11334 ( .I1(n10729), .I2(n10731), .O(n10742) );
  NAND_GATE U11335 ( .I1(n10731), .I2(n10730), .O(n10736) );
  NAND_GATE U11336 ( .I1(n10732), .I2(n10736), .O(n10740) );
  NAND_GATE U11337 ( .I1(n10734), .I2(n10733), .O(n10735) );
  NAND_GATE U11338 ( .I1(n10736), .I2(n10735), .O(n10737) );
  NAND_GATE U11339 ( .I1(n10738), .I2(n10737), .O(n10739) );
  NAND_GATE U11340 ( .I1(n10740), .I2(n10739), .O(n10741) );
  NAND_GATE U11341 ( .I1(n10742), .I2(n10741), .O(n11128) );
  OR_GATE U11342 ( .I1(n10743), .I2(n10747), .O(n10746) );
  OR_GATE U11343 ( .I1(n10744), .I2(n10748), .O(n10745) );
  AND_GATE U11344 ( .I1(n10746), .I2(n10745), .O(n10753) );
  NAND_GATE U11345 ( .I1(n10747), .I2(n1004), .O(n10751) );
  NAND3_GATE U11346 ( .I1(n10751), .I2(n10750), .I3(n10749), .O(n10752) );
  NAND_GATE U11347 ( .I1(n10753), .I2(n10752), .O(n11136) );
  INV_GATE U11348 ( .I1(n11136), .O(n11139) );
  OR_GATE U11349 ( .I1(n10754), .I2(n10756), .O(n10767) );
  NAND_GATE U11350 ( .I1(n10756), .I2(n10755), .O(n10761) );
  NAND_GATE U11351 ( .I1(n10757), .I2(n10761), .O(n10765) );
  NAND_GATE U11352 ( .I1(n10759), .I2(n10758), .O(n10760) );
  NAND_GATE U11353 ( .I1(n10761), .I2(n10760), .O(n10762) );
  NAND_GATE U11354 ( .I1(n10763), .I2(n10762), .O(n10764) );
  NAND_GATE U11355 ( .I1(n10765), .I2(n10764), .O(n10766) );
  NAND_GATE U11356 ( .I1(n10767), .I2(n10766), .O(n11152) );
  OR_GATE U11357 ( .I1(n10768), .I2(n10772), .O(n10771) );
  OR_GATE U11358 ( .I1(n10769), .I2(n10773), .O(n10770) );
  AND_GATE U11359 ( .I1(n10771), .I2(n10770), .O(n10778) );
  NAND_GATE U11360 ( .I1(n10772), .I2(n1013), .O(n10776) );
  NAND3_GATE U11361 ( .I1(n10776), .I2(n10775), .I3(n10774), .O(n10777) );
  NAND_GATE U11362 ( .I1(n10778), .I2(n10777), .O(n11161) );
  INV_GATE U11363 ( .I1(n11161), .O(n11164) );
  OR_GATE U11364 ( .I1(n10779), .I2(n10781), .O(n10792) );
  NAND_GATE U11365 ( .I1(n10781), .I2(n10780), .O(n10786) );
  NAND_GATE U11366 ( .I1(n10782), .I2(n10786), .O(n10790) );
  NAND_GATE U11367 ( .I1(n10784), .I2(n10783), .O(n10785) );
  NAND_GATE U11368 ( .I1(n10786), .I2(n10785), .O(n10787) );
  NAND_GATE U11369 ( .I1(n10788), .I2(n10787), .O(n10789) );
  NAND_GATE U11370 ( .I1(n10790), .I2(n10789), .O(n10791) );
  NAND_GATE U11371 ( .I1(n10792), .I2(n10791), .O(n11177) );
  OR_GATE U11372 ( .I1(n10793), .I2(n10797), .O(n10796) );
  OR_GATE U11373 ( .I1(n10794), .I2(n10798), .O(n10795) );
  AND_GATE U11374 ( .I1(n10796), .I2(n10795), .O(n10803) );
  NAND_GATE U11375 ( .I1(n10797), .I2(n1172), .O(n10801) );
  NAND3_GATE U11376 ( .I1(n10801), .I2(n10800), .I3(n10799), .O(n10802) );
  NAND_GATE U11377 ( .I1(n10803), .I2(n10802), .O(n11186) );
  INV_GATE U11378 ( .I1(n11186), .O(n11189) );
  OR_GATE U11379 ( .I1(n10804), .I2(n10806), .O(n10817) );
  NAND_GATE U11380 ( .I1(n10806), .I2(n10805), .O(n10811) );
  NAND_GATE U11381 ( .I1(n10807), .I2(n10811), .O(n10815) );
  NAND_GATE U11382 ( .I1(n10809), .I2(n10808), .O(n10810) );
  NAND_GATE U11383 ( .I1(n10811), .I2(n10810), .O(n10812) );
  NAND_GATE U11384 ( .I1(n10813), .I2(n10812), .O(n10814) );
  NAND_GATE U11385 ( .I1(n10815), .I2(n10814), .O(n10816) );
  NAND_GATE U11386 ( .I1(n10817), .I2(n10816), .O(n11202) );
  NAND_GATE U11387 ( .I1(n1374), .I2(A[0]), .O(n10818) );
  NAND_GATE U11388 ( .I1(n14781), .I2(n10818), .O(n10819) );
  NAND_GATE U11389 ( .I1(B[11]), .I2(n10819), .O(n10823) );
  NAND_GATE U11390 ( .I1(n1375), .I2(A[1]), .O(n10820) );
  NAND_GATE U11391 ( .I1(n14784), .I2(n10820), .O(n10821) );
  NAND_GATE U11392 ( .I1(B[10]), .I2(n10821), .O(n10822) );
  NAND_GATE U11393 ( .I1(n10823), .I2(n10822), .O(n11214) );
  NAND_GATE U11394 ( .I1(B[9]), .I2(A[2]), .O(n11218) );
  NAND3_GATE U11395 ( .I1(B[9]), .I2(B[10]), .I3(n1196), .O(n11211) );
  NAND_GATE U11396 ( .I1(n11218), .I2(n11211), .O(n10824) );
  NAND_GATE U11397 ( .I1(n11214), .I2(n10824), .O(n10825) );
  INV_GATE U11398 ( .I1(n11218), .O(n11212) );
  INV_GATE U11399 ( .I1(n11211), .O(n11213) );
  NAND_GATE U11400 ( .I1(n11212), .I2(n11213), .O(n11209) );
  NAND_GATE U11401 ( .I1(n10825), .I2(n11209), .O(n11203) );
  NAND_GATE U11402 ( .I1(n11202), .I2(n11203), .O(n10827) );
  NAND_GATE U11403 ( .I1(B[9]), .I2(A[3]), .O(n11204) );
  INV_GATE U11404 ( .I1(n11204), .O(n10826) );
  NAND_GATE U11405 ( .I1(n11202), .I2(n10826), .O(n11199) );
  NAND_GATE U11406 ( .I1(n11203), .I2(n10826), .O(n11198) );
  NAND3_GATE U11407 ( .I1(n10827), .I2(n11199), .I3(n11198), .O(n11188) );
  INV_GATE U11408 ( .I1(n11188), .O(n11185) );
  NAND_GATE U11409 ( .I1(B[9]), .I2(A[4]), .O(n11193) );
  NAND_GATE U11410 ( .I1(n11185), .I2(n11193), .O(n10828) );
  NAND_GATE U11411 ( .I1(n11189), .I2(n10828), .O(n10829) );
  INV_GATE U11412 ( .I1(n11193), .O(n11187) );
  NAND_GATE U11413 ( .I1(n11188), .I2(n11187), .O(n11184) );
  NAND_GATE U11414 ( .I1(n10829), .I2(n11184), .O(n11178) );
  NAND_GATE U11415 ( .I1(n11177), .I2(n11178), .O(n10831) );
  NAND_GATE U11416 ( .I1(B[9]), .I2(A[5]), .O(n11179) );
  INV_GATE U11417 ( .I1(n11179), .O(n10830) );
  NAND_GATE U11418 ( .I1(n11177), .I2(n10830), .O(n11174) );
  NAND_GATE U11419 ( .I1(n11178), .I2(n10830), .O(n11173) );
  NAND3_GATE U11420 ( .I1(n10831), .I2(n11174), .I3(n11173), .O(n11163) );
  INV_GATE U11421 ( .I1(n11163), .O(n11160) );
  NAND_GATE U11422 ( .I1(B[9]), .I2(A[6]), .O(n11168) );
  NAND_GATE U11423 ( .I1(n11160), .I2(n11168), .O(n10832) );
  NAND_GATE U11424 ( .I1(n11164), .I2(n10832), .O(n10833) );
  INV_GATE U11425 ( .I1(n11168), .O(n11162) );
  NAND_GATE U11426 ( .I1(n11163), .I2(n11162), .O(n11159) );
  NAND_GATE U11427 ( .I1(n10833), .I2(n11159), .O(n11153) );
  NAND_GATE U11428 ( .I1(n11152), .I2(n11153), .O(n10835) );
  NAND_GATE U11429 ( .I1(B[9]), .I2(A[7]), .O(n11154) );
  INV_GATE U11430 ( .I1(n11154), .O(n10834) );
  NAND_GATE U11431 ( .I1(n11152), .I2(n10834), .O(n11149) );
  NAND_GATE U11432 ( .I1(n11153), .I2(n10834), .O(n11148) );
  NAND3_GATE U11433 ( .I1(n10835), .I2(n11149), .I3(n11148), .O(n11138) );
  INV_GATE U11434 ( .I1(n11138), .O(n11135) );
  NAND_GATE U11435 ( .I1(B[9]), .I2(A[8]), .O(n11143) );
  NAND_GATE U11436 ( .I1(n11135), .I2(n11143), .O(n10836) );
  NAND_GATE U11437 ( .I1(n11139), .I2(n10836), .O(n10837) );
  INV_GATE U11438 ( .I1(n11143), .O(n11137) );
  NAND_GATE U11439 ( .I1(n11138), .I2(n11137), .O(n11134) );
  NAND_GATE U11440 ( .I1(n10837), .I2(n11134), .O(n11129) );
  NAND_GATE U11441 ( .I1(n11128), .I2(n11129), .O(n10839) );
  NAND_GATE U11442 ( .I1(B[9]), .I2(A[9]), .O(n11130) );
  INV_GATE U11443 ( .I1(n11130), .O(n10838) );
  NAND_GATE U11444 ( .I1(n11128), .I2(n10838), .O(n11125) );
  NAND_GATE U11445 ( .I1(n11129), .I2(n10838), .O(n11124) );
  NAND3_GATE U11446 ( .I1(n10839), .I2(n11125), .I3(n11124), .O(n11116) );
  INV_GATE U11447 ( .I1(n11116), .O(n11113) );
  NAND_GATE U11448 ( .I1(B[9]), .I2(A[10]), .O(n11121) );
  NAND_GATE U11449 ( .I1(n11113), .I2(n11121), .O(n10840) );
  NAND_GATE U11450 ( .I1(n11117), .I2(n10840), .O(n10841) );
  INV_GATE U11451 ( .I1(n11121), .O(n11115) );
  NAND_GATE U11452 ( .I1(n11116), .I2(n11115), .O(n11112) );
  NAND_GATE U11453 ( .I1(n10841), .I2(n11112), .O(n11254) );
  NAND_GATE U11454 ( .I1(n11253), .I2(n11254), .O(n10843) );
  NAND_GATE U11455 ( .I1(B[9]), .I2(A[11]), .O(n11255) );
  INV_GATE U11456 ( .I1(n11255), .O(n10842) );
  NAND_GATE U11457 ( .I1(n11254), .I2(n10842), .O(n11250) );
  NAND_GATE U11458 ( .I1(n11253), .I2(n10842), .O(n11249) );
  NAND_GATE U11459 ( .I1(n11102), .I2(n11107), .O(n10844) );
  NAND_GATE U11460 ( .I1(n11104), .I2(n10844), .O(n10845) );
  NAND_GATE U11461 ( .I1(n11101), .I2(n10845), .O(n11096) );
  NAND_GATE U11462 ( .I1(n10857), .I2(n11096), .O(n11092) );
  INV_GATE U11463 ( .I1(n10846), .O(n10847) );
  NAND_GATE U11464 ( .I1(n10847), .I2(n10850), .O(n10856) );
  INV_GATE U11465 ( .I1(n10850), .O(n10848) );
  NAND_GATE U11466 ( .I1(n10849), .I2(n10848), .O(n10851) );
  NAND_GATE U11467 ( .I1(n695), .I2(n10851), .O(n10854) );
  NAND_GATE U11468 ( .I1(n10854), .I2(n10853), .O(n10855) );
  NAND_GATE U11469 ( .I1(n10856), .I2(n10855), .O(n11095) );
  NAND_GATE U11470 ( .I1(n11096), .I2(n11095), .O(n10858) );
  NAND_GATE U11471 ( .I1(n10857), .I2(n11095), .O(n11091) );
  NAND3_GATE U11472 ( .I1(n11092), .I2(n10858), .I3(n11091), .O(n11271) );
  NAND_GATE U11473 ( .I1(n11269), .I2(n11274), .O(n10859) );
  NAND_GATE U11474 ( .I1(n11271), .I2(n10859), .O(n10860) );
  NAND_GATE U11475 ( .I1(n11266), .I2(n10860), .O(n11086) );
  NAND3_GATE U11476 ( .I1(n11083), .I2(n11084), .I3(n11086), .O(n10862) );
  NAND_GATE U11477 ( .I1(n10861), .I2(n11086), .O(n11078) );
  NAND3_GATE U11478 ( .I1(n11077), .I2(n10862), .I3(n11078), .O(n11288) );
  NAND_GATE U11479 ( .I1(n11287), .I2(n11291), .O(n10863) );
  NAND_GATE U11480 ( .I1(n11288), .I2(n10863), .O(n10864) );
  NAND_GATE U11481 ( .I1(n11283), .I2(n10864), .O(n11070) );
  NAND_GATE U11482 ( .I1(n10872), .I2(n11070), .O(n11063) );
  NAND_GATE U11483 ( .I1(n566), .I2(n10870), .O(n10865) );
  NAND_GATE U11484 ( .I1(n10865), .I2(n10868), .O(n11059) );
  NAND_GATE U11485 ( .I1(n10867), .I2(n10866), .O(n10868) );
  NAND_GATE U11486 ( .I1(n10869), .I2(n10868), .O(n11062) );
  NAND3_GATE U11487 ( .I1(n10870), .I2(n566), .I3(n10869), .O(n11071) );
  NAND3_GATE U11488 ( .I1(n11070), .I2(n11061), .I3(n10871), .O(n10873) );
  NAND3_GATE U11489 ( .I1(n10872), .I2(n11061), .I3(n10871), .O(n11064) );
  NAND3_GATE U11490 ( .I1(n11063), .I2(n10873), .I3(n11064), .O(n11056) );
  NAND_GATE U11491 ( .I1(n11048), .I2(n11052), .O(n10874) );
  NAND_GATE U11492 ( .I1(n11056), .I2(n10874), .O(n10875) );
  NAND_GATE U11493 ( .I1(n11055), .I2(n10875), .O(n11040) );
  NAND_GATE U11494 ( .I1(n11034), .I2(n11040), .O(n11035) );
  INV_GATE U11495 ( .I1(n10876), .O(n10877) );
  NAND_GATE U11496 ( .I1(n10877), .I2(n10882), .O(n10889) );
  INV_GATE U11497 ( .I1(n10882), .O(n10880) );
  NAND_GATE U11498 ( .I1(n10881), .I2(n10880), .O(n10878) );
  NAND_GATE U11499 ( .I1(n10879), .I2(n10878), .O(n10887) );
  NAND_GATE U11500 ( .I1(n505), .I2(n10882), .O(n10883) );
  NAND_GATE U11501 ( .I1(n10878), .I2(n10883), .O(n10884) );
  NAND_GATE U11502 ( .I1(n10885), .I2(n10884), .O(n10886) );
  NAND_GATE U11503 ( .I1(n10887), .I2(n10886), .O(n10888) );
  NAND_GATE U11504 ( .I1(n10889), .I2(n10888), .O(n11039) );
  NAND_GATE U11505 ( .I1(n11040), .I2(n11039), .O(n10891) );
  NAND_GATE U11506 ( .I1(n11034), .I2(n11039), .O(n10890) );
  NAND3_GATE U11507 ( .I1(n11035), .I2(n10891), .I3(n10890), .O(n11309) );
  NAND_GATE U11508 ( .I1(n11307), .I2(n11305), .O(n10892) );
  NAND_GATE U11509 ( .I1(n11309), .I2(n10892), .O(n10893) );
  NAND_GATE U11510 ( .I1(n11308), .I2(n10893), .O(n11027) );
  NAND_GATE U11511 ( .I1(n10906), .I2(n11027), .O(n11029) );
  NAND_GATE U11512 ( .I1(n10897), .I2(n1259), .O(n10894) );
  NAND_GATE U11513 ( .I1(n10895), .I2(n10894), .O(n10900) );
  NAND_GATE U11514 ( .I1(n603), .I2(n10902), .O(n10899) );
  NAND3_GATE U11515 ( .I1(n10897), .I2(n1259), .I3(n10896), .O(n10898) );
  NAND3_GATE U11516 ( .I1(n10900), .I2(n10899), .I3(n10898), .O(n10905) );
  INV_GATE U11517 ( .I1(n10901), .O(n10903) );
  NAND_GATE U11518 ( .I1(n10903), .I2(n10902), .O(n10904) );
  NAND_GATE U11519 ( .I1(n10905), .I2(n10904), .O(n11030) );
  NAND_GATE U11520 ( .I1(n11027), .I2(n11030), .O(n10907) );
  NAND_GATE U11521 ( .I1(n10906), .I2(n11030), .O(n11028) );
  NAND3_GATE U11522 ( .I1(n11029), .I2(n10907), .I3(n11028), .O(n11325) );
  NAND_GATE U11523 ( .I1(n11316), .I2(n11318), .O(n10908) );
  NAND_GATE U11524 ( .I1(n11325), .I2(n10908), .O(n10909) );
  NAND_GATE U11525 ( .I1(n11324), .I2(n10909), .O(n11016) );
  NAND_GATE U11526 ( .I1(n10915), .I2(n11016), .O(n11012) );
  NAND_GATE U11527 ( .I1(n10914), .I2(n678), .O(n10910) );
  NAND_GATE U11528 ( .I1(n10911), .I2(n10910), .O(n11009) );
  INV_GATE U11529 ( .I1(n11009), .O(n10913) );
  NAND_GATE U11530 ( .I1(n10913), .I2(n11011), .O(n10917) );
  NAND3_GATE U11531 ( .I1(n10915), .I2(n10917), .I3(n10916), .O(n11007) );
  NAND3_GATE U11532 ( .I1(n11016), .I2(n10917), .I3(n10916), .O(n10918) );
  NAND3_GATE U11533 ( .I1(n11012), .I2(n11007), .I3(n10918), .O(n11343) );
  NAND_GATE U11534 ( .I1(n11334), .I2(n11336), .O(n10919) );
  NAND_GATE U11535 ( .I1(n11343), .I2(n10919), .O(n10920) );
  NAND_GATE U11536 ( .I1(n11825), .I2(n11003), .O(n10921) );
  NAND_GATE U11537 ( .I1(n11001), .I2(n10921), .O(n10922) );
  NAND_GATE U11538 ( .I1(n10923), .I2(n10922), .O(n10996) );
  NAND_GATE U11539 ( .I1(n11458), .I2(n10995), .O(n10924) );
  NAND_GATE U11540 ( .I1(n10996), .I2(n10924), .O(n10925) );
  NAND_GATE U11541 ( .I1(n11440), .I2(n11436), .O(n10927) );
  NAND_GATE U11542 ( .I1(n11435), .I2(n10927), .O(n10928) );
  NAND_GATE U11543 ( .I1(n10929), .I2(n10928), .O(n11414) );
  NAND_GATE U11544 ( .I1(n11417), .I2(n11415), .O(n10930) );
  NAND_GATE U11545 ( .I1(n11414), .I2(n10930), .O(n10931) );
  NAND_GATE U11546 ( .I1(n10932), .I2(n10931), .O(n11361) );
  NAND_GATE U11547 ( .I1(n10936), .I2(n10935), .O(n10939) );
  NAND_GATE U11548 ( .I1(n10940), .I2(n10939), .O(n10937) );
  NAND_GATE U11549 ( .I1(n10938), .I2(n10937), .O(n10942) );
  NAND3_GATE U11550 ( .I1(n10946), .I2(n10940), .I3(n10939), .O(n10941) );
  NAND3_GATE U11551 ( .I1(n10943), .I2(n10942), .I3(n10941), .O(n10950) );
  OR_GATE U11552 ( .I1(n10945), .I2(n10944), .O(n10949) );
  NAND3_GATE U11553 ( .I1(n10947), .I2(n10946), .I3(n10945), .O(n10948) );
  AND_GATE U11554 ( .I1(n10949), .I2(n10948), .O(n10951) );
  NAND3_GATE U11555 ( .I1(n11361), .I2(n10950), .I3(n10951), .O(n10954) );
  NAND_GATE U11556 ( .I1(B[9]), .I2(A[29]), .O(n11396) );
  INV_GATE U11557 ( .I1(n11396), .O(n11392) );
  NAND_GATE U11558 ( .I1(n11392), .I2(n11361), .O(n10953) );
  NAND_GATE U11559 ( .I1(n10951), .I2(n10950), .O(n11363) );
  NAND_GATE U11560 ( .I1(n263), .I2(n10951), .O(n10952) );
  NAND3_GATE U11561 ( .I1(n10954), .I2(n10953), .I3(n10952), .O(n10984) );
  NAND_GATE U11562 ( .I1(n10982), .I2(n10983), .O(n10955) );
  NAND_GATE U11563 ( .I1(n15343), .I2(n10971), .O(n10956) );
  NAND_GATE U11564 ( .I1(n10975), .I2(n10956), .O(n10957) );
  NAND_GATE U11565 ( .I1(n10958), .I2(n10957), .O(n10967) );
  OR_GATE U11566 ( .I1(n10960), .I2(n10959), .O(n10964) );
  AND_GATE U11567 ( .I1(n10964), .I2(n10963), .O(n10966) );
  NAND3_GATE U11568 ( .I1(n10965), .I2(n10967), .I3(n10966), .O(n15341) );
  AND_GATE U11569 ( .I1(n10966), .I2(n10965), .O(n10968) );
  OR_GATE U11570 ( .I1(n10968), .I2(n10967), .O(n10969) );
  AND_GATE U11571 ( .I1(n15341), .I2(n10969), .O(\A1[39] ) );
  NAND_GATE U11572 ( .I1(n10970), .I2(n10972), .O(n15342) );
  NAND_GATE U11573 ( .I1(n10971), .I2(n1294), .O(n10972) );
  NAND3_GATE U11574 ( .I1(n10975), .I2(n10974), .I3(n10973), .O(n15347) );
  NAND_GATE U11575 ( .I1(n1251), .I2(n15347), .O(n11370) );
  NAND_GATE U11576 ( .I1(B[8]), .I2(A[31]), .O(n11377) );
  INV_GATE U11577 ( .I1(n11377), .O(n11378) );
  NAND_GATE U11578 ( .I1(n1356), .I2(n10984), .O(n10989) );
  NAND_GATE U11579 ( .I1(n10977), .I2(n10976), .O(n10978) );
  NAND3_GATE U11580 ( .I1(n10983), .I2(n973), .I3(n10982), .O(n10986) );
  NAND3_GATE U11581 ( .I1(n10987), .I2(n10986), .I3(n10985), .O(n10988) );
  NAND_GATE U11582 ( .I1(n10989), .I2(n10988), .O(n11381) );
  NAND_GATE U11583 ( .I1(n11378), .I2(n11381), .O(n11368) );
  NAND_GATE U11584 ( .I1(B[8]), .I2(A[30]), .O(n11404) );
  INV_GATE U11585 ( .I1(n11404), .O(n11386) );
  NAND_GATE U11586 ( .I1(B[8]), .I2(A[29]), .O(n11425) );
  INV_GATE U11587 ( .I1(n11425), .O(n11407) );
  NAND_GATE U11588 ( .I1(B[8]), .I2(A[28]), .O(n11446) );
  INV_GATE U11589 ( .I1(n11446), .O(n11430) );
  NAND3_GATE U11590 ( .I1(n10990), .I2(n11435), .I3(n738), .O(n11434) );
  NAND3_GATE U11591 ( .I1(n11436), .I2(n792), .I3(n11440), .O(n10991) );
  NAND_GATE U11592 ( .I1(n10990), .I2(n11437), .O(n11433) );
  NAND3_GATE U11593 ( .I1(n10991), .I2(n11438), .I3(n11433), .O(n10992) );
  NAND_GATE U11594 ( .I1(n11434), .I2(n10992), .O(n11429) );
  NAND_GATE U11595 ( .I1(n11430), .I2(n11429), .O(n11354) );
  NAND_GATE U11596 ( .I1(B[8]), .I2(A[27]), .O(n11452) );
  INV_GATE U11597 ( .I1(n11452), .O(n11456) );
  INV_GATE U11598 ( .I1(n10996), .O(n10994) );
  NAND_GATE U11599 ( .I1(n10993), .I2(n10999), .O(n11460) );
  NAND3_GATE U11600 ( .I1(n10996), .I2(n10997), .I3(n10993), .O(n11455) );
  NAND_GATE U11601 ( .I1(n10995), .I2(n10994), .O(n10999) );
  NAND_GATE U11602 ( .I1(n10997), .I2(n10996), .O(n10998) );
  NAND_GATE U11603 ( .I1(n10999), .I2(n10998), .O(n11457) );
  NAND3_GATE U11604 ( .I1(n11456), .I2(n11451), .I3(n11459), .O(n11464) );
  NAND_GATE U11605 ( .I1(B[8]), .I2(A[26]), .O(n11819) );
  INV_GATE U11606 ( .I1(n11819), .O(n11349) );
  NAND3_GATE U11607 ( .I1(n11001), .I2(n11002), .I3(n11000), .O(n11828) );
  NAND_GATE U11608 ( .I1(n826), .I2(n11828), .O(n11006) );
  NAND_GATE U11609 ( .I1(n11003), .I2(n154), .O(n11004) );
  NAND_GATE U11610 ( .I1(n11005), .I2(n11004), .O(n11824) );
  NAND3_GATE U11611 ( .I1(n11349), .I2(n11006), .I3(n11826), .O(n11822) );
  NAND_GATE U11612 ( .I1(B[8]), .I2(A[25]), .O(n11469) );
  INV_GATE U11613 ( .I1(n11469), .O(n11470) );
  NAND_GATE U11614 ( .I1(B[8]), .I2(A[24]), .O(n11476) );
  INV_GATE U11615 ( .I1(n11476), .O(n11483) );
  OR_GATE U11616 ( .I1(n11007), .I2(n11016), .O(n11014) );
  NAND_GATE U11617 ( .I1(n11011), .I2(n11010), .O(n11015) );
  OR_GATE U11618 ( .I1(n11015), .I2(n11012), .O(n11013) );
  AND_GATE U11619 ( .I1(n11014), .I2(n11013), .O(n11021) );
  NAND_GATE U11620 ( .I1(n954), .I2(n11015), .O(n11018) );
  NAND3_GATE U11621 ( .I1(n11019), .I2(n11018), .I3(n11017), .O(n11020) );
  NAND_GATE U11622 ( .I1(n11021), .I2(n11020), .O(n11478) );
  NAND_GATE U11623 ( .I1(n11483), .I2(n668), .O(n11333) );
  NAND_GATE U11624 ( .I1(B[8]), .I2(A[23]), .O(n11498) );
  INV_GATE U11625 ( .I1(n11498), .O(n11489) );
  NAND_GATE U11626 ( .I1(B[8]), .I2(A[22]), .O(n11800) );
  INV_GATE U11627 ( .I1(n11800), .O(n11796) );
  INV_GATE U11628 ( .I1(n11030), .O(n11022) );
  NAND_GATE U11629 ( .I1(n11027), .I2(n11022), .O(n11025) );
  INV_GATE U11630 ( .I1(n11027), .O(n11023) );
  NAND_GATE U11631 ( .I1(n11023), .I2(n11030), .O(n11024) );
  NAND3_GATE U11632 ( .I1(n11026), .I2(n11025), .I3(n11024), .O(n11033) );
  OR_GATE U11633 ( .I1(n11028), .I2(n11027), .O(n11032) );
  OR_GATE U11634 ( .I1(n11030), .I2(n11029), .O(n11031) );
  NAND3_GATE U11635 ( .I1(n11033), .I2(n11032), .I3(n11031), .O(n11799) );
  NAND_GATE U11636 ( .I1(n11796), .I2(n11797), .O(n11803) );
  NAND_GATE U11637 ( .I1(B[8]), .I2(A[21]), .O(n11508) );
  INV_GATE U11638 ( .I1(n11508), .O(n11311) );
  NAND_GATE U11639 ( .I1(B[8]), .I2(A[20]), .O(n11783) );
  INV_GATE U11640 ( .I1(n11783), .O(n11779) );
  INV_GATE U11641 ( .I1(n11040), .O(n11038) );
  NAND3_GATE U11642 ( .I1(n11034), .I2(n11038), .I3(n11039), .O(n11037) );
  OR_GATE U11643 ( .I1(n11039), .I2(n11035), .O(n11036) );
  AND_GATE U11644 ( .I1(n11037), .I2(n11036), .O(n11045) );
  NAND_GATE U11645 ( .I1(n11038), .I2(n11039), .O(n11043) );
  NAND3_GATE U11646 ( .I1(n11043), .I2(n11042), .I3(n11041), .O(n11044) );
  NAND_GATE U11647 ( .I1(n11045), .I2(n11044), .O(n11780) );
  NAND_GATE U11648 ( .I1(n11779), .I2(n1202), .O(n11786) );
  NAND_GATE U11649 ( .I1(B[8]), .I2(A[19]), .O(n11518) );
  INV_GATE U11650 ( .I1(n11518), .O(n11300) );
  INV_GATE U11651 ( .I1(n11056), .O(n11047) );
  NAND_GATE U11652 ( .I1(n11046), .I2(n11050), .O(n11054) );
  NAND_GATE U11653 ( .I1(n11048), .I2(n11047), .O(n11050) );
  NAND_GATE U11654 ( .I1(n1327), .I2(n11056), .O(n11049) );
  NAND_GATE U11655 ( .I1(n11050), .I2(n11049), .O(n11051) );
  NAND_GATE U11656 ( .I1(n11052), .I2(n11051), .O(n11053) );
  NAND_GATE U11657 ( .I1(n11054), .I2(n11053), .O(n11058) );
  NAND_GATE U11658 ( .I1(n11058), .I2(n11057), .O(n11521) );
  NAND_GATE U11659 ( .I1(n11300), .I2(n11521), .O(n11523) );
  NAND_GATE U11660 ( .I1(n11060), .I2(n11059), .O(n11061) );
  NAND_GATE U11661 ( .I1(n11062), .I2(n11061), .O(n11069) );
  NAND_GATE U11662 ( .I1(n11071), .I2(n11069), .O(n11067) );
  OR_GATE U11663 ( .I1(n11067), .I2(n11063), .O(n11066) );
  OR_GATE U11664 ( .I1(n11064), .I2(n11070), .O(n11065) );
  AND_GATE U11665 ( .I1(n11066), .I2(n11065), .O(n11076) );
  INV_GATE U11666 ( .I1(n11070), .O(n11068) );
  NAND_GATE U11667 ( .I1(n11068), .I2(n11067), .O(n11074) );
  NAND3_GATE U11668 ( .I1(n11071), .I2(n11070), .I3(n11069), .O(n11073) );
  NAND3_GATE U11669 ( .I1(n11074), .I2(n11073), .I3(n11072), .O(n11075) );
  NAND_GATE U11670 ( .I1(n11076), .I2(n11075), .O(n11767) );
  NAND_GATE U11671 ( .I1(B[8]), .I2(A[18]), .O(n11765) );
  INV_GATE U11672 ( .I1(n11765), .O(n11764) );
  NAND_GATE U11673 ( .I1(n233), .I2(n11764), .O(n11761) );
  NAND_GATE U11674 ( .I1(B[8]), .I2(A[17]), .O(n11534) );
  INV_GATE U11675 ( .I1(n11534), .O(n11296) );
  OR_GATE U11676 ( .I1(n11077), .I2(n11086), .O(n11080) );
  OR_GATE U11677 ( .I1(n11081), .I2(n11078), .O(n11079) );
  INV_GATE U11678 ( .I1(n11086), .O(n11082) );
  NAND_GATE U11679 ( .I1(n11082), .I2(n11081), .O(n11089) );
  NAND_GATE U11680 ( .I1(n11084), .I2(n11083), .O(n11085) );
  NAND_GATE U11681 ( .I1(n11086), .I2(n11085), .O(n11088) );
  NAND3_GATE U11682 ( .I1(n11089), .I2(n11088), .I3(n11087), .O(n11090) );
  INV_GATE U11683 ( .I1(n11541), .O(n11543) );
  NAND_GATE U11684 ( .I1(B[8]), .I2(A[16]), .O(n11547) );
  INV_GATE U11685 ( .I1(n11547), .O(n11540) );
  NAND_GATE U11686 ( .I1(B[8]), .I2(A[15]), .O(n11556) );
  INV_GATE U11687 ( .I1(n11556), .O(n11279) );
  OR_GATE U11688 ( .I1(n11091), .I2(n11096), .O(n11094) );
  OR_GATE U11689 ( .I1(n11095), .I2(n11092), .O(n11093) );
  NAND_GATE U11690 ( .I1(n965), .I2(n11095), .O(n11099) );
  NAND3_GATE U11691 ( .I1(n11099), .I2(n11098), .I3(n11097), .O(n11100) );
  NAND_GATE U11692 ( .I1(B[8]), .I2(A[14]), .O(n11567) );
  INV_GATE U11693 ( .I1(n11567), .O(n11564) );
  NAND_GATE U11694 ( .I1(n101), .I2(n11564), .O(n11560) );
  NAND_GATE U11695 ( .I1(n11102), .I2(n752), .O(n11106) );
  NAND_GATE U11696 ( .I1(n11103), .I2(n11106), .O(n11109) );
  NAND_GATE U11697 ( .I1(n11109), .I2(n11108), .O(n11110) );
  NAND_GATE U11698 ( .I1(n11111), .I2(n11110), .O(n11744) );
  OR_GATE U11699 ( .I1(n11112), .I2(n11114), .O(n11123) );
  NAND_GATE U11700 ( .I1(n11114), .I2(n11113), .O(n11119) );
  NAND_GATE U11701 ( .I1(n11115), .I2(n11119), .O(n11122) );
  NAND_GATE U11702 ( .I1(n11117), .I2(n11116), .O(n11118) );
  NAND_GATE U11703 ( .I1(n11119), .I2(n11118), .O(n11120) );
  OR_GATE U11704 ( .I1(n11124), .I2(n11128), .O(n11127) );
  OR_GATE U11705 ( .I1(n11125), .I2(n11129), .O(n11126) );
  NAND_GATE U11706 ( .I1(n11128), .I2(n998), .O(n11132) );
  NAND3_GATE U11707 ( .I1(n11132), .I2(n11131), .I3(n11130), .O(n11133) );
  INV_GATE U11708 ( .I1(n11586), .O(n11589) );
  OR_GATE U11709 ( .I1(n11134), .I2(n11136), .O(n11147) );
  NAND_GATE U11710 ( .I1(n11136), .I2(n11135), .O(n11141) );
  NAND_GATE U11711 ( .I1(n11137), .I2(n11141), .O(n11145) );
  NAND_GATE U11712 ( .I1(n11139), .I2(n11138), .O(n11140) );
  NAND_GATE U11713 ( .I1(n11141), .I2(n11140), .O(n11142) );
  NAND_GATE U11714 ( .I1(n11143), .I2(n11142), .O(n11144) );
  NAND_GATE U11715 ( .I1(n11145), .I2(n11144), .O(n11146) );
  NAND_GATE U11716 ( .I1(n11147), .I2(n11146), .O(n11602) );
  OR_GATE U11717 ( .I1(n11148), .I2(n11152), .O(n11151) );
  OR_GATE U11718 ( .I1(n11149), .I2(n11153), .O(n11150) );
  AND_GATE U11719 ( .I1(n11151), .I2(n11150), .O(n11158) );
  NAND_GATE U11720 ( .I1(n11152), .I2(n1009), .O(n11156) );
  NAND3_GATE U11721 ( .I1(n11156), .I2(n11155), .I3(n11154), .O(n11157) );
  NAND_GATE U11722 ( .I1(n11158), .I2(n11157), .O(n11611) );
  INV_GATE U11723 ( .I1(n11611), .O(n11614) );
  OR_GATE U11724 ( .I1(n11159), .I2(n11161), .O(n11172) );
  NAND_GATE U11725 ( .I1(n11161), .I2(n11160), .O(n11166) );
  NAND_GATE U11726 ( .I1(n11162), .I2(n11166), .O(n11170) );
  NAND_GATE U11727 ( .I1(n11164), .I2(n11163), .O(n11165) );
  NAND_GATE U11728 ( .I1(n11166), .I2(n11165), .O(n11167) );
  NAND_GATE U11729 ( .I1(n11168), .I2(n11167), .O(n11169) );
  NAND_GATE U11730 ( .I1(n11170), .I2(n11169), .O(n11171) );
  NAND_GATE U11731 ( .I1(n11172), .I2(n11171), .O(n11627) );
  OR_GATE U11732 ( .I1(n11173), .I2(n11177), .O(n11176) );
  OR_GATE U11733 ( .I1(n11174), .I2(n11178), .O(n11175) );
  AND_GATE U11734 ( .I1(n11176), .I2(n11175), .O(n11183) );
  NAND_GATE U11735 ( .I1(n11177), .I2(n1105), .O(n11181) );
  NAND3_GATE U11736 ( .I1(n11181), .I2(n11180), .I3(n11179), .O(n11182) );
  NAND_GATE U11737 ( .I1(n11183), .I2(n11182), .O(n11636) );
  INV_GATE U11738 ( .I1(n11636), .O(n11639) );
  OR_GATE U11739 ( .I1(n11184), .I2(n11186), .O(n11197) );
  NAND_GATE U11740 ( .I1(n11186), .I2(n11185), .O(n11191) );
  NAND_GATE U11741 ( .I1(n11187), .I2(n11191), .O(n11195) );
  NAND_GATE U11742 ( .I1(n11189), .I2(n11188), .O(n11190) );
  NAND_GATE U11743 ( .I1(n11191), .I2(n11190), .O(n11192) );
  NAND_GATE U11744 ( .I1(n11193), .I2(n11192), .O(n11194) );
  NAND_GATE U11745 ( .I1(n11195), .I2(n11194), .O(n11196) );
  NAND_GATE U11746 ( .I1(n11197), .I2(n11196), .O(n11652) );
  OR_GATE U11747 ( .I1(n11198), .I2(n11202), .O(n11201) );
  OR_GATE U11748 ( .I1(n11199), .I2(n11203), .O(n11200) );
  AND_GATE U11749 ( .I1(n11201), .I2(n11200), .O(n11208) );
  NAND_GATE U11750 ( .I1(n11202), .I2(n1183), .O(n11206) );
  NAND3_GATE U11751 ( .I1(n11206), .I2(n11205), .I3(n11204), .O(n11207) );
  NAND_GATE U11752 ( .I1(n11208), .I2(n11207), .O(n11661) );
  INV_GATE U11753 ( .I1(n11661), .O(n11664) );
  INV_GATE U11754 ( .I1(n11209), .O(n11210) );
  NAND_GATE U11755 ( .I1(n11214), .I2(n11210), .O(n11222) );
  NAND_GATE U11756 ( .I1(n11212), .I2(n11216), .O(n11220) );
  NAND_GATE U11757 ( .I1(n11214), .I2(n11213), .O(n11215) );
  NAND_GATE U11758 ( .I1(n11216), .I2(n11215), .O(n11217) );
  NAND_GATE U11759 ( .I1(n11218), .I2(n11217), .O(n11219) );
  NAND_GATE U11760 ( .I1(n11220), .I2(n11219), .O(n11221) );
  NAND_GATE U11761 ( .I1(n11222), .I2(n11221), .O(n11677) );
  NAND_GATE U11762 ( .I1(n1373), .I2(A[0]), .O(n11223) );
  NAND_GATE U11763 ( .I1(n14781), .I2(n11223), .O(n11224) );
  NAND_GATE U11764 ( .I1(B[10]), .I2(n11224), .O(n11228) );
  NAND_GATE U11765 ( .I1(n1374), .I2(A[1]), .O(n11225) );
  NAND_GATE U11766 ( .I1(n14784), .I2(n11225), .O(n11226) );
  NAND_GATE U11767 ( .I1(B[9]), .I2(n11226), .O(n11227) );
  NAND_GATE U11768 ( .I1(n11228), .I2(n11227), .O(n11689) );
  NAND_GATE U11769 ( .I1(B[8]), .I2(A[2]), .O(n11693) );
  NAND3_GATE U11770 ( .I1(B[8]), .I2(B[9]), .I3(n1196), .O(n11686) );
  NAND_GATE U11771 ( .I1(n11693), .I2(n11686), .O(n11229) );
  NAND_GATE U11772 ( .I1(n11689), .I2(n11229), .O(n11230) );
  INV_GATE U11773 ( .I1(n11693), .O(n11687) );
  INV_GATE U11774 ( .I1(n11686), .O(n11688) );
  NAND_GATE U11775 ( .I1(n11687), .I2(n11688), .O(n11684) );
  NAND_GATE U11776 ( .I1(n11230), .I2(n11684), .O(n11678) );
  NAND_GATE U11777 ( .I1(n11677), .I2(n11678), .O(n11232) );
  NAND_GATE U11778 ( .I1(B[8]), .I2(A[3]), .O(n11679) );
  INV_GATE U11779 ( .I1(n11679), .O(n11231) );
  NAND_GATE U11780 ( .I1(n11677), .I2(n11231), .O(n11674) );
  NAND_GATE U11781 ( .I1(n11678), .I2(n11231), .O(n11673) );
  NAND3_GATE U11782 ( .I1(n11232), .I2(n11674), .I3(n11673), .O(n11663) );
  INV_GATE U11783 ( .I1(n11663), .O(n11660) );
  NAND_GATE U11784 ( .I1(B[8]), .I2(A[4]), .O(n11668) );
  NAND_GATE U11785 ( .I1(n11660), .I2(n11668), .O(n11233) );
  NAND_GATE U11786 ( .I1(n11664), .I2(n11233), .O(n11234) );
  INV_GATE U11787 ( .I1(n11668), .O(n11662) );
  NAND_GATE U11788 ( .I1(n11663), .I2(n11662), .O(n11659) );
  NAND_GATE U11789 ( .I1(n11234), .I2(n11659), .O(n11653) );
  NAND_GATE U11790 ( .I1(n11652), .I2(n11653), .O(n11236) );
  NAND_GATE U11791 ( .I1(B[8]), .I2(A[5]), .O(n11654) );
  INV_GATE U11792 ( .I1(n11654), .O(n11235) );
  NAND_GATE U11793 ( .I1(n11652), .I2(n11235), .O(n11649) );
  NAND_GATE U11794 ( .I1(n11653), .I2(n11235), .O(n11648) );
  NAND3_GATE U11795 ( .I1(n11236), .I2(n11649), .I3(n11648), .O(n11638) );
  INV_GATE U11796 ( .I1(n11638), .O(n11635) );
  NAND_GATE U11797 ( .I1(B[8]), .I2(A[6]), .O(n11643) );
  NAND_GATE U11798 ( .I1(n11635), .I2(n11643), .O(n11237) );
  NAND_GATE U11799 ( .I1(n11639), .I2(n11237), .O(n11238) );
  INV_GATE U11800 ( .I1(n11643), .O(n11637) );
  NAND_GATE U11801 ( .I1(n11638), .I2(n11637), .O(n11634) );
  NAND_GATE U11802 ( .I1(n11238), .I2(n11634), .O(n11628) );
  NAND_GATE U11803 ( .I1(n11627), .I2(n11628), .O(n11240) );
  NAND_GATE U11804 ( .I1(B[8]), .I2(A[7]), .O(n11629) );
  INV_GATE U11805 ( .I1(n11629), .O(n11239) );
  NAND_GATE U11806 ( .I1(n11627), .I2(n11239), .O(n11624) );
  NAND_GATE U11807 ( .I1(n11628), .I2(n11239), .O(n11623) );
  NAND3_GATE U11808 ( .I1(n11240), .I2(n11624), .I3(n11623), .O(n11613) );
  INV_GATE U11809 ( .I1(n11613), .O(n11610) );
  NAND_GATE U11810 ( .I1(B[8]), .I2(A[8]), .O(n11618) );
  NAND_GATE U11811 ( .I1(n11610), .I2(n11618), .O(n11241) );
  NAND_GATE U11812 ( .I1(n11614), .I2(n11241), .O(n11242) );
  INV_GATE U11813 ( .I1(n11618), .O(n11612) );
  NAND_GATE U11814 ( .I1(n11613), .I2(n11612), .O(n11609) );
  NAND_GATE U11815 ( .I1(n11242), .I2(n11609), .O(n11603) );
  NAND_GATE U11816 ( .I1(n11602), .I2(n11603), .O(n11244) );
  NAND_GATE U11817 ( .I1(B[8]), .I2(A[9]), .O(n11604) );
  INV_GATE U11818 ( .I1(n11604), .O(n11243) );
  NAND_GATE U11819 ( .I1(n11602), .I2(n11243), .O(n11599) );
  NAND_GATE U11820 ( .I1(n11603), .I2(n11243), .O(n11598) );
  NAND3_GATE U11821 ( .I1(n11244), .I2(n11599), .I3(n11598), .O(n11588) );
  INV_GATE U11822 ( .I1(n11588), .O(n11585) );
  NAND_GATE U11823 ( .I1(B[8]), .I2(A[10]), .O(n11593) );
  NAND_GATE U11824 ( .I1(n11585), .I2(n11593), .O(n11245) );
  NAND_GATE U11825 ( .I1(n11589), .I2(n11245), .O(n11246) );
  INV_GATE U11826 ( .I1(n11593), .O(n11587) );
  NAND_GATE U11827 ( .I1(n11588), .I2(n11587), .O(n11584) );
  NAND_GATE U11828 ( .I1(n11246), .I2(n11584), .O(n11729) );
  NAND_GATE U11829 ( .I1(n11728), .I2(n11729), .O(n11248) );
  NAND_GATE U11830 ( .I1(B[8]), .I2(A[11]), .O(n11730) );
  INV_GATE U11831 ( .I1(n11730), .O(n11247) );
  NAND_GATE U11832 ( .I1(n11729), .I2(n11247), .O(n11725) );
  NAND_GATE U11833 ( .I1(n11728), .I2(n11247), .O(n11724) );
  NAND3_GATE U11834 ( .I1(n11248), .I2(n11725), .I3(n11724), .O(n11577) );
  NAND_GATE U11835 ( .I1(B[8]), .I2(A[12]), .O(n11579) );
  OR_GATE U11836 ( .I1(n11249), .I2(n11254), .O(n11252) );
  OR_GATE U11837 ( .I1(n11250), .I2(n11253), .O(n11251) );
  AND_GATE U11838 ( .I1(n11252), .I2(n11251), .O(n11259) );
  NAND_GATE U11839 ( .I1(n11253), .I2(n938), .O(n11257) );
  NAND3_GATE U11840 ( .I1(n11257), .I2(n11256), .I3(n11255), .O(n11258) );
  NAND_GATE U11841 ( .I1(n11259), .I2(n11258), .O(n11573) );
  NAND_GATE U11842 ( .I1(n11579), .I2(n11573), .O(n11260) );
  NAND_GATE U11843 ( .I1(n11577), .I2(n11260), .O(n11261) );
  INV_GATE U11844 ( .I1(n11579), .O(n11575) );
  INV_GATE U11845 ( .I1(n11573), .O(n11576) );
  NAND_GATE U11846 ( .I1(n11575), .I2(n11576), .O(n11572) );
  NAND_GATE U11847 ( .I1(n11261), .I2(n11572), .O(n11745) );
  NAND_GATE U11848 ( .I1(n11744), .I2(n11745), .O(n11263) );
  NAND_GATE U11849 ( .I1(B[8]), .I2(A[13]), .O(n11746) );
  INV_GATE U11850 ( .I1(n11746), .O(n11262) );
  NAND_GATE U11851 ( .I1(n11745), .I2(n11262), .O(n11740) );
  NAND_GATE U11852 ( .I1(n11744), .I2(n11262), .O(n11739) );
  NAND3_GATE U11853 ( .I1(n11263), .I2(n11740), .I3(n11739), .O(n11565) );
  NAND_GATE U11854 ( .I1(n11563), .I2(n11567), .O(n11264) );
  NAND_GATE U11855 ( .I1(n11565), .I2(n11264), .O(n11265) );
  NAND_GATE U11856 ( .I1(n11560), .I2(n11265), .O(n11555) );
  NAND_GATE U11857 ( .I1(n11279), .I2(n11555), .O(n11551) );
  INV_GATE U11858 ( .I1(n11266), .O(n11267) );
  NAND_GATE U11859 ( .I1(n11267), .I2(n11271), .O(n11278) );
  INV_GATE U11860 ( .I1(n11271), .O(n11268) );
  NAND_GATE U11861 ( .I1(n11269), .I2(n11268), .O(n11273) );
  NAND_GATE U11862 ( .I1(n11270), .I2(n11273), .O(n11276) );
  NAND_GATE U11863 ( .I1(n11276), .I2(n11275), .O(n11277) );
  NAND_GATE U11864 ( .I1(n11278), .I2(n11277), .O(n11554) );
  NAND_GATE U11865 ( .I1(n11555), .I2(n11554), .O(n11280) );
  NAND_GATE U11866 ( .I1(n11279), .I2(n11554), .O(n11550) );
  NAND_GATE U11867 ( .I1(n11541), .I2(n11547), .O(n11281) );
  NAND_GATE U11868 ( .I1(n11542), .I2(n11281), .O(n11282) );
  NAND_GATE U11869 ( .I1(n11539), .I2(n11282), .O(n11533) );
  NAND_GATE U11870 ( .I1(n11296), .I2(n11533), .O(n11529) );
  INV_GATE U11871 ( .I1(n11283), .O(n11284) );
  NAND_GATE U11872 ( .I1(n11284), .I2(n11288), .O(n11295) );
  INV_GATE U11873 ( .I1(n11288), .O(n11286) );
  NAND_GATE U11874 ( .I1(n11285), .I2(n11290), .O(n11293) );
  NAND_GATE U11875 ( .I1(n11287), .I2(n11286), .O(n11290) );
  NAND_GATE U11876 ( .I1(n11293), .I2(n11292), .O(n11294) );
  NAND_GATE U11877 ( .I1(n11295), .I2(n11294), .O(n11532) );
  NAND_GATE U11878 ( .I1(n11533), .I2(n11532), .O(n11297) );
  NAND_GATE U11879 ( .I1(n11296), .I2(n11532), .O(n11528) );
  NAND3_GATE U11880 ( .I1(n11529), .I2(n11297), .I3(n11528), .O(n11768) );
  NAND_GATE U11881 ( .I1(n11767), .I2(n11765), .O(n11298) );
  NAND_GATE U11882 ( .I1(n11768), .I2(n11298), .O(n11299) );
  NAND_GATE U11883 ( .I1(n11761), .I2(n11299), .O(n11524) );
  NAND_GATE U11884 ( .I1(n11521), .I2(n11524), .O(n11301) );
  NAND_GATE U11885 ( .I1(n11300), .I2(n11524), .O(n11522) );
  NAND3_GATE U11886 ( .I1(n11523), .I2(n11301), .I3(n11522), .O(n11787) );
  NAND_GATE U11887 ( .I1(n11783), .I2(n11780), .O(n11302) );
  NAND_GATE U11888 ( .I1(n11787), .I2(n11302), .O(n11303) );
  NAND_GATE U11889 ( .I1(n11786), .I2(n11303), .O(n11511) );
  NAND_GATE U11890 ( .I1(n11311), .I2(n11511), .O(n11513) );
  NAND3_GATE U11891 ( .I1(n11304), .I2(n11309), .I3(n11305), .O(n11503) );
  INV_GATE U11892 ( .I1(n11309), .O(n11306) );
  NAND3_GATE U11893 ( .I1(n11307), .I2(n11306), .I3(n11305), .O(n11505) );
  NAND_GATE U11894 ( .I1(n11307), .I2(n11306), .O(n11501) );
  NAND3_GATE U11895 ( .I1(n11502), .I2(n11501), .I3(n11507), .O(n11310) );
  NAND3_GATE U11896 ( .I1(n11511), .I2(n947), .I3(n11310), .O(n11312) );
  NAND3_GATE U11897 ( .I1(n11311), .I2(n947), .I3(n11310), .O(n11512) );
  NAND3_GATE U11898 ( .I1(n11513), .I2(n11312), .I3(n11512), .O(n11804) );
  NAND_GATE U11899 ( .I1(n11800), .I2(n11799), .O(n11313) );
  NAND_GATE U11900 ( .I1(n11804), .I2(n11313), .O(n11314) );
  NAND_GATE U11901 ( .I1(n11315), .I2(n11325), .O(n11323) );
  INV_GATE U11902 ( .I1(n11325), .O(n11317) );
  NAND3_GATE U11903 ( .I1(n11318), .I2(n11317), .I3(n11316), .O(n11322) );
  NAND_GATE U11904 ( .I1(n11318), .I2(n11317), .O(n11319) );
  NAND_GATE U11905 ( .I1(n11320), .I2(n11319), .O(n11321) );
  NAND3_GATE U11906 ( .I1(n11323), .I2(n11322), .I3(n11321), .O(n11328) );
  INV_GATE U11907 ( .I1(n11324), .O(n11326) );
  NAND_GATE U11908 ( .I1(n11326), .I2(n11325), .O(n11327) );
  NAND_GATE U11909 ( .I1(n11328), .I2(n11327), .O(n11494) );
  NAND_GATE U11910 ( .I1(n11495), .I2(n11494), .O(n11330) );
  NAND_GATE U11911 ( .I1(n11489), .I2(n11494), .O(n11329) );
  NAND3_GATE U11912 ( .I1(n11490), .I2(n11330), .I3(n11329), .O(n11479) );
  NAND_GATE U11913 ( .I1(n11476), .I2(n11478), .O(n11331) );
  NAND_GATE U11914 ( .I1(n11479), .I2(n11331), .O(n11332) );
  NAND_GATE U11915 ( .I1(n11333), .I2(n11332), .O(n11466) );
  NAND_GATE U11916 ( .I1(n11470), .I2(n11466), .O(n11471) );
  INV_GATE U11917 ( .I1(n11343), .O(n11335) );
  NAND3_GATE U11918 ( .I1(n11336), .I2(n11335), .I3(n11334), .O(n11341) );
  NAND_GATE U11919 ( .I1(n243), .I2(n11343), .O(n11340) );
  NAND_GATE U11920 ( .I1(n11336), .I2(n11335), .O(n11337) );
  NAND_GATE U11921 ( .I1(n11338), .I2(n11337), .O(n11339) );
  NAND3_GATE U11922 ( .I1(n11341), .I2(n11340), .I3(n11339), .O(n11346) );
  INV_GATE U11923 ( .I1(n11342), .O(n11344) );
  NAND_GATE U11924 ( .I1(n11344), .I2(n11343), .O(n11345) );
  NAND_GATE U11925 ( .I1(n11346), .I2(n11345), .O(n11472) );
  NAND_GATE U11926 ( .I1(n11470), .I2(n11472), .O(n11348) );
  NAND_GATE U11927 ( .I1(n11466), .I2(n11472), .O(n11347) );
  NAND3_GATE U11928 ( .I1(n11471), .I2(n11348), .I3(n11347), .O(n11823) );
  NAND3_GATE U11929 ( .I1(n11006), .I2(n11823), .I3(n11826), .O(n11350) );
  NAND_GATE U11930 ( .I1(n11349), .I2(n11823), .O(n11827) );
  NAND3_GATE U11931 ( .I1(n11822), .I2(n11350), .I3(n11827), .O(n11461) );
  NAND_GATE U11932 ( .I1(n11456), .I2(n11461), .O(n11352) );
  NAND3_GATE U11933 ( .I1(n11451), .I2(n11459), .I3(n11461), .O(n11351) );
  NAND3_GATE U11934 ( .I1(n11464), .I2(n11352), .I3(n11351), .O(n11442) );
  NAND_GATE U11935 ( .I1(n11442), .I2(n11429), .O(n11353) );
  NAND_GATE U11936 ( .I1(n11430), .I2(n11442), .O(n11428) );
  NAND3_GATE U11937 ( .I1(n11354), .I2(n11353), .I3(n11428), .O(n11422) );
  NAND_GATE U11938 ( .I1(n11407), .I2(n11422), .O(n11408) );
  NAND3_GATE U11939 ( .I1(n11355), .I2(n11414), .I3(n621), .O(n11413) );
  NAND3_GATE U11940 ( .I1(n11415), .I2(n585), .I3(n11417), .O(n11357) );
  NAND_GATE U11941 ( .I1(n621), .I2(n11414), .O(n11356) );
  NAND_GATE U11942 ( .I1(n11355), .I2(n11416), .O(n11412) );
  NAND3_GATE U11943 ( .I1(n11357), .I2(n11356), .I3(n11412), .O(n11358) );
  NAND_GATE U11944 ( .I1(n11413), .I2(n11358), .O(n11409) );
  NAND_GATE U11945 ( .I1(n11407), .I2(n11409), .O(n11360) );
  NAND_GATE U11946 ( .I1(n11422), .I2(n11409), .O(n11359) );
  NAND3_GATE U11947 ( .I1(n11408), .I2(n11360), .I3(n11359), .O(n11401) );
  NAND_GATE U11948 ( .I1(n11386), .I2(n11401), .O(n11388) );
  NAND3_GATE U11949 ( .I1(n11392), .I2(n11361), .I3(n1221), .O(n11393) );
  NAND_GATE U11950 ( .I1(n11363), .I2(n11362), .O(n11394) );
  NAND_GATE U11951 ( .I1(n11392), .I2(n11394), .O(n11385) );
  NAND_GATE U11952 ( .I1(n1221), .I2(n11361), .O(n11364) );
  NAND_GATE U11953 ( .I1(n11364), .I2(n11394), .O(n11395) );
  NAND3_GATE U11954 ( .I1(n11388), .I2(n11366), .I3(n11365), .O(n11374) );
  NAND_GATE U11955 ( .I1(n11374), .I2(n11381), .O(n11367) );
  NAND_GATE U11956 ( .I1(n11378), .I2(n11374), .O(n11380) );
  NAND3_GATE U11957 ( .I1(n11368), .I2(n11367), .I3(n11380), .O(n15349) );
  INV_GATE U11958 ( .I1(n15349), .O(n11369) );
  NAND3_GATE U11959 ( .I1(n15344), .I2(n11370), .I3(n11369), .O(n11373) );
  NAND_GATE U11960 ( .I1(n11370), .I2(n15344), .O(n11371) );
  NAND_GATE U11961 ( .I1(n15349), .I2(n11371), .O(n11372) );
  NAND_GATE U11962 ( .I1(n11373), .I2(n11372), .O(\A1[38] ) );
  NAND_GATE U11963 ( .I1(n11379), .I2(n11381), .O(n11376) );
  NAND3_GATE U11964 ( .I1(n11377), .I2(n11376), .I3(n11375), .O(n11384) );
  NAND3_GATE U11965 ( .I1(n11379), .I2(n11381), .I3(n11378), .O(n11383) );
  OR_GATE U11966 ( .I1(n11381), .I2(n11380), .O(n11382) );
  NAND3_GATE U11967 ( .I1(n11384), .I2(n11383), .I3(n11382), .O(n11849) );
  NAND_GATE U11968 ( .I1(B[7]), .I2(A[31]), .O(n15351) );
  INV_GATE U11969 ( .I1(n11401), .O(n11397) );
  NAND4_GATE U11970 ( .I1(n11386), .I2(n11397), .I3(n11387), .I4(n11398), .O(
        n11391) );
  AND_GATE U11971 ( .I1(n11387), .I2(n11398), .O(n11389) );
  OR_GATE U11972 ( .I1(n11389), .I2(n11388), .O(n11390) );
  AND_GATE U11973 ( .I1(n11391), .I2(n11390), .O(n11406) );
  NAND3_GATE U11974 ( .I1(n11394), .I2(n11393), .I3(n11392), .O(n11399) );
  NAND_GATE U11975 ( .I1(n11396), .I2(n11395), .O(n11398) );
  NAND3_GATE U11976 ( .I1(n11399), .I2(n11398), .I3(n11397), .O(n11403) );
  NAND_GATE U11977 ( .I1(n11399), .I2(n11398), .O(n11400) );
  NAND_GATE U11978 ( .I1(n11401), .I2(n11400), .O(n11402) );
  NAND3_GATE U11979 ( .I1(n11404), .I2(n11403), .I3(n11402), .O(n11405) );
  NAND_GATE U11980 ( .I1(n11406), .I2(n11405), .O(n11852) );
  INV_GATE U11981 ( .I1(n11852), .O(n11853) );
  NAND_GATE U11982 ( .I1(n1220), .I2(n11853), .O(n11848) );
  NAND_GATE U11983 ( .I1(B[7]), .I2(A[30]), .O(n12271) );
  INV_GATE U11984 ( .I1(n12271), .O(n12250) );
  NAND3_GATE U11985 ( .I1(n11407), .I2(n11418), .I3(n11409), .O(n11411) );
  OR_GATE U11986 ( .I1(n11409), .I2(n11408), .O(n11410) );
  AND_GATE U11987 ( .I1(n11411), .I2(n11410), .O(n11427) );
  NAND3_GATE U11988 ( .I1(n11420), .I2(n11418), .I3(n11419), .O(n11424) );
  NAND_GATE U11989 ( .I1(n11420), .I2(n11419), .O(n11421) );
  NAND_GATE U11990 ( .I1(n11422), .I2(n11421), .O(n11423) );
  NAND3_GATE U11991 ( .I1(n11425), .I2(n11424), .I3(n11423), .O(n11426) );
  NAND_GATE U11992 ( .I1(n11427), .I2(n11426), .O(n12268) );
  NAND_GATE U11993 ( .I1(n12250), .I2(n623), .O(n11845) );
  NAND_GATE U11994 ( .I1(B[7]), .I2(A[29]), .O(n12238) );
  INV_GATE U11995 ( .I1(n12238), .O(n12235) );
  OR_GATE U11996 ( .I1(n11429), .I2(n11428), .O(n11432) );
  INV_GATE U11997 ( .I1(n11442), .O(n11443) );
  NAND3_GATE U11998 ( .I1(n11430), .I2(n11443), .I3(n11429), .O(n11431) );
  NAND_GATE U11999 ( .I1(n11432), .I2(n11431), .O(n12232) );
  NAND_GATE U12000 ( .I1(n738), .I2(n11435), .O(n11438) );
  NAND_GATE U12001 ( .I1(n11436), .I2(n792), .O(n11437) );
  NAND_GATE U12002 ( .I1(n11438), .I2(n11437), .O(n11439) );
  NAND_GATE U12003 ( .I1(n11440), .I2(n11439), .O(n11444) );
  NAND_GATE U12004 ( .I1(n11445), .I2(n11444), .O(n11441) );
  NAND_GATE U12005 ( .I1(n11442), .I2(n11441), .O(n11448) );
  NAND3_GATE U12006 ( .I1(n11445), .I2(n11444), .I3(n11443), .O(n11447) );
  NAND3_GATE U12007 ( .I1(n11448), .I2(n11447), .I3(n11446), .O(n12231) );
  NAND_GATE U12008 ( .I1(n11449), .I2(n12231), .O(n12236) );
  NAND_GATE U12009 ( .I1(n11451), .I2(n11459), .O(n11450) );
  NAND_GATE U12010 ( .I1(n11461), .I2(n11450), .O(n11454) );
  INV_GATE U12011 ( .I1(n11461), .O(n11465) );
  NAND3_GATE U12012 ( .I1(n11451), .I2(n11459), .I3(n11465), .O(n11453) );
  NAND3_GATE U12013 ( .I1(n11454), .I2(n11453), .I3(n11452), .O(n11855) );
  NAND_GATE U12014 ( .I1(B[7]), .I2(A[28]), .O(n12292) );
  INV_GATE U12015 ( .I1(n12292), .O(n11856) );
  AND_GATE U12016 ( .I1(n11456), .I2(n11455), .O(n11463) );
  NAND_GATE U12017 ( .I1(n11458), .I2(n11457), .O(n11459) );
  NAND_GATE U12018 ( .I1(n11460), .I2(n11459), .O(n11462) );
  NAND3_GATE U12019 ( .I1(n11463), .I2(n11462), .I3(n11461), .O(n11838) );
  NAND3_GATE U12020 ( .I1(n11855), .I2(n11856), .I3(n915), .O(n11857) );
  NAND_GATE U12021 ( .I1(B[7]), .I2(A[26]), .O(n12332) );
  INV_GATE U12022 ( .I1(n12332), .O(n11873) );
  NAND_GATE U12023 ( .I1(n765), .I2(n11472), .O(n11468) );
  NAND_GATE U12024 ( .I1(n11466), .I2(n602), .O(n11467) );
  NAND3_GATE U12025 ( .I1(n11469), .I2(n11468), .I3(n11467), .O(n11475) );
  NAND3_GATE U12026 ( .I1(n765), .I2(n11472), .I3(n11470), .O(n11474) );
  OR_GATE U12027 ( .I1(n11472), .I2(n11471), .O(n11473) );
  NAND3_GATE U12028 ( .I1(n11475), .I2(n11474), .I3(n11473), .O(n11874) );
  INV_GATE U12029 ( .I1(n11874), .O(n11876) );
  NAND_GATE U12030 ( .I1(n11873), .I2(n11876), .O(n11816) );
  NAND3_GATE U12031 ( .I1(n11476), .I2(n11479), .I3(n668), .O(n11486) );
  NAND3_GATE U12032 ( .I1(n11478), .I2(n11477), .I3(n11476), .O(n11485) );
  AND_GATE U12033 ( .I1(n11486), .I2(n11485), .O(n11481) );
  NAND_GATE U12034 ( .I1(n11478), .I2(n11477), .O(n11482) );
  NAND3_GATE U12035 ( .I1(n11479), .I2(n668), .I3(n11483), .O(n11488) );
  NAND3_GATE U12036 ( .I1(n11482), .I2(n11488), .I3(n11483), .O(n11480) );
  NAND_GATE U12037 ( .I1(B[7]), .I2(A[25]), .O(n11888) );
  INV_GATE U12038 ( .I1(n11888), .O(n11812) );
  NAND3_GATE U12039 ( .I1(n11481), .I2(n11480), .I3(n11812), .O(n11879) );
  NAND_GATE U12040 ( .I1(n11483), .I2(n11482), .O(n11484) );
  NAND3_GATE U12041 ( .I1(n11486), .I2(n11485), .I3(n11484), .O(n11487) );
  NAND_GATE U12042 ( .I1(n11488), .I2(n11487), .O(n11885) );
  NAND_GATE U12043 ( .I1(B[7]), .I2(A[24]), .O(n11894) );
  INV_GATE U12044 ( .I1(n11894), .O(n11892) );
  NAND3_GATE U12045 ( .I1(n11493), .I2(n11489), .I3(n11494), .O(n11492) );
  OR_GATE U12046 ( .I1(n11494), .I2(n11490), .O(n11491) );
  AND_GATE U12047 ( .I1(n11492), .I2(n11491), .O(n11500) );
  NAND_GATE U12048 ( .I1(n11493), .I2(n11494), .O(n11497) );
  NAND3_GATE U12049 ( .I1(n11498), .I2(n11497), .I3(n11496), .O(n11499) );
  NAND_GATE U12050 ( .I1(n11500), .I2(n11499), .O(n11895) );
  INV_GATE U12051 ( .I1(n11895), .O(n11893) );
  NAND_GATE U12052 ( .I1(B[7]), .I2(A[23]), .O(n11905) );
  INV_GATE U12053 ( .I1(n11905), .O(n11808) );
  NAND_GATE U12054 ( .I1(n11502), .I2(n11501), .O(n11504) );
  NAND3_GATE U12055 ( .I1(n11505), .I2(n11504), .I3(n11503), .O(n11506) );
  NAND_GATE U12056 ( .I1(n11507), .I2(n11506), .O(n11514) );
  NAND_GATE U12057 ( .I1(n957), .I2(n11514), .O(n11510) );
  NAND3_GATE U12058 ( .I1(n11510), .I2(n11509), .I3(n11508), .O(n11517) );
  OR_GATE U12059 ( .I1(n11512), .I2(n11511), .O(n11516) );
  OR_GATE U12060 ( .I1(n11514), .I2(n11513), .O(n11515) );
  NAND3_GATE U12061 ( .I1(n11517), .I2(n11516), .I3(n11515), .O(n12208) );
  NAND_GATE U12062 ( .I1(B[7]), .I2(A[22]), .O(n12211) );
  INV_GATE U12063 ( .I1(n12211), .O(n12206) );
  NAND_GATE U12064 ( .I1(n12210), .I2(n12206), .O(n12203) );
  NAND_GATE U12065 ( .I1(B[7]), .I2(A[21]), .O(n11921) );
  INV_GATE U12066 ( .I1(n11921), .O(n11791) );
  NAND_GATE U12067 ( .I1(n11521), .I2(n234), .O(n11520) );
  NAND_GATE U12068 ( .I1(n1340), .I2(n11524), .O(n11519) );
  NAND3_GATE U12069 ( .I1(n11520), .I2(n11519), .I3(n11518), .O(n11527) );
  OR_GATE U12070 ( .I1(n11522), .I2(n11521), .O(n11526) );
  OR_GATE U12071 ( .I1(n11524), .I2(n11523), .O(n11525) );
  NAND3_GATE U12072 ( .I1(n11527), .I2(n11526), .I3(n11525), .O(n12189) );
  NAND_GATE U12073 ( .I1(B[7]), .I2(A[20]), .O(n12194) );
  INV_GATE U12074 ( .I1(n12194), .O(n12187) );
  NAND_GATE U12075 ( .I1(n1326), .I2(n12187), .O(n12186) );
  NAND_GATE U12076 ( .I1(B[7]), .I2(A[19]), .O(n11929) );
  INV_GATE U12077 ( .I1(n11929), .O(n11774) );
  OR_GATE U12078 ( .I1(n11532), .I2(n11529), .O(n11530) );
  AND_GATE U12079 ( .I1(n11531), .I2(n11530), .O(n11538) );
  NAND_GATE U12080 ( .I1(n928), .I2(n11532), .O(n11536) );
  NAND3_GATE U12081 ( .I1(n11536), .I2(n11535), .I3(n11534), .O(n11537) );
  NAND_GATE U12082 ( .I1(n11538), .I2(n11537), .O(n12172) );
  NAND_GATE U12083 ( .I1(B[7]), .I2(A[18]), .O(n12177) );
  INV_GATE U12084 ( .I1(n12177), .O(n12171) );
  NAND_GATE U12085 ( .I1(n605), .I2(n12171), .O(n12169) );
  NAND_GATE U12086 ( .I1(B[7]), .I2(A[17]), .O(n11943) );
  INV_GATE U12087 ( .I1(n11943), .O(n11757) );
  NAND_GATE U12088 ( .I1(n11540), .I2(n11545), .O(n11548) );
  NAND_GATE U12089 ( .I1(n11541), .I2(n719), .O(n11545) );
  NAND_GATE U12090 ( .I1(n11543), .I2(n11542), .O(n11544) );
  NAND_GATE U12091 ( .I1(n11545), .I2(n11544), .O(n11546) );
  NAND_GATE U12092 ( .I1(n11757), .I2(n11938), .O(n11934) );
  NAND_GATE U12093 ( .I1(n11547), .I2(n11546), .O(n11939) );
  OR_GATE U12094 ( .I1(n11550), .I2(n11555), .O(n11553) );
  OR_GATE U12095 ( .I1(n11554), .I2(n11551), .O(n11552) );
  NAND_GATE U12096 ( .I1(n933), .I2(n11554), .O(n11558) );
  NAND3_GATE U12097 ( .I1(n11558), .I2(n11557), .I3(n11556), .O(n11559) );
  INV_GATE U12098 ( .I1(n11950), .O(n11953) );
  NAND_GATE U12099 ( .I1(B[7]), .I2(A[16]), .O(n11955) );
  INV_GATE U12100 ( .I1(n11955), .O(n11951) );
  NAND_GATE U12101 ( .I1(n11953), .I2(n11951), .O(n11948) );
  INV_GATE U12102 ( .I1(n11560), .O(n11561) );
  NAND_GATE U12103 ( .I1(n11561), .I2(n11565), .O(n11571) );
  INV_GATE U12104 ( .I1(n11565), .O(n11562) );
  NAND_GATE U12105 ( .I1(n11563), .I2(n11562), .O(n11566) );
  NAND_GATE U12106 ( .I1(n11564), .I2(n11566), .O(n11569) );
  NAND_GATE U12107 ( .I1(n11569), .I2(n11568), .O(n11570) );
  NAND_GATE U12108 ( .I1(n11571), .I2(n11570), .O(n12156) );
  INV_GATE U12109 ( .I1(n11577), .O(n11574) );
  NAND_GATE U12110 ( .I1(n11574), .I2(n11573), .O(n11578) );
  NAND_GATE U12111 ( .I1(n11575), .I2(n11578), .O(n11581) );
  NAND_GATE U12112 ( .I1(n11581), .I2(n11580), .O(n11582) );
  NAND_GATE U12113 ( .I1(n11583), .I2(n11582), .O(n12141) );
  OR_GATE U12114 ( .I1(n11584), .I2(n11586), .O(n11597) );
  NAND_GATE U12115 ( .I1(n11586), .I2(n11585), .O(n11591) );
  NAND_GATE U12116 ( .I1(n11587), .I2(n11591), .O(n11595) );
  NAND_GATE U12117 ( .I1(n11589), .I2(n11588), .O(n11590) );
  NAND_GATE U12118 ( .I1(n11591), .I2(n11590), .O(n11592) );
  NAND_GATE U12119 ( .I1(n11593), .I2(n11592), .O(n11594) );
  NAND_GATE U12120 ( .I1(n11595), .I2(n11594), .O(n11596) );
  NAND_GATE U12121 ( .I1(n11597), .I2(n11596), .O(n12127) );
  OR_GATE U12122 ( .I1(n11598), .I2(n11602), .O(n11601) );
  OR_GATE U12123 ( .I1(n11599), .I2(n11603), .O(n11600) );
  AND_GATE U12124 ( .I1(n11601), .I2(n11600), .O(n11608) );
  NAND_GATE U12125 ( .I1(n11602), .I2(n1005), .O(n11606) );
  NAND3_GATE U12126 ( .I1(n11606), .I2(n11605), .I3(n11604), .O(n11607) );
  NAND_GATE U12127 ( .I1(n11608), .I2(n11607), .O(n11985) );
  INV_GATE U12128 ( .I1(n11985), .O(n11988) );
  OR_GATE U12129 ( .I1(n11609), .I2(n11611), .O(n11622) );
  NAND_GATE U12130 ( .I1(n11611), .I2(n11610), .O(n11616) );
  NAND_GATE U12131 ( .I1(n11612), .I2(n11616), .O(n11620) );
  NAND_GATE U12132 ( .I1(n11614), .I2(n11613), .O(n11615) );
  NAND_GATE U12133 ( .I1(n11616), .I2(n11615), .O(n11617) );
  NAND_GATE U12134 ( .I1(n11618), .I2(n11617), .O(n11619) );
  NAND_GATE U12135 ( .I1(n11620), .I2(n11619), .O(n11621) );
  NAND_GATE U12136 ( .I1(n11622), .I2(n11621), .O(n12001) );
  OR_GATE U12137 ( .I1(n11623), .I2(n11627), .O(n11626) );
  OR_GATE U12138 ( .I1(n11624), .I2(n11628), .O(n11625) );
  AND_GATE U12139 ( .I1(n11626), .I2(n11625), .O(n11633) );
  NAND_GATE U12140 ( .I1(n11627), .I2(n1014), .O(n11631) );
  NAND3_GATE U12141 ( .I1(n11631), .I2(n11630), .I3(n11629), .O(n11632) );
  NAND_GATE U12142 ( .I1(n11633), .I2(n11632), .O(n12010) );
  INV_GATE U12143 ( .I1(n12010), .O(n12013) );
  OR_GATE U12144 ( .I1(n11634), .I2(n11636), .O(n11647) );
  NAND_GATE U12145 ( .I1(n11636), .I2(n11635), .O(n11641) );
  NAND_GATE U12146 ( .I1(n11637), .I2(n11641), .O(n11645) );
  NAND_GATE U12147 ( .I1(n11639), .I2(n11638), .O(n11640) );
  NAND_GATE U12148 ( .I1(n11641), .I2(n11640), .O(n11642) );
  NAND_GATE U12149 ( .I1(n11643), .I2(n11642), .O(n11644) );
  NAND_GATE U12150 ( .I1(n11645), .I2(n11644), .O(n11646) );
  NAND_GATE U12151 ( .I1(n11647), .I2(n11646), .O(n12026) );
  OR_GATE U12152 ( .I1(n11648), .I2(n11652), .O(n11651) );
  OR_GATE U12153 ( .I1(n11649), .I2(n11653), .O(n11650) );
  AND_GATE U12154 ( .I1(n11651), .I2(n11650), .O(n11658) );
  NAND_GATE U12155 ( .I1(n11652), .I2(n1109), .O(n11656) );
  NAND3_GATE U12156 ( .I1(n11656), .I2(n11655), .I3(n11654), .O(n11657) );
  NAND_GATE U12157 ( .I1(n11658), .I2(n11657), .O(n12035) );
  INV_GATE U12158 ( .I1(n12035), .O(n12038) );
  OR_GATE U12159 ( .I1(n11659), .I2(n11661), .O(n11672) );
  NAND_GATE U12160 ( .I1(n11661), .I2(n11660), .O(n11666) );
  NAND_GATE U12161 ( .I1(n11662), .I2(n11666), .O(n11670) );
  NAND_GATE U12162 ( .I1(n11664), .I2(n11663), .O(n11665) );
  NAND_GATE U12163 ( .I1(n11666), .I2(n11665), .O(n11667) );
  NAND_GATE U12164 ( .I1(n11668), .I2(n11667), .O(n11669) );
  NAND_GATE U12165 ( .I1(n11670), .I2(n11669), .O(n11671) );
  NAND_GATE U12166 ( .I1(n11672), .I2(n11671), .O(n12051) );
  OR_GATE U12167 ( .I1(n11673), .I2(n11677), .O(n11676) );
  OR_GATE U12168 ( .I1(n11674), .I2(n11678), .O(n11675) );
  AND_GATE U12169 ( .I1(n11676), .I2(n11675), .O(n11683) );
  NAND_GATE U12170 ( .I1(n11677), .I2(n1184), .O(n11681) );
  NAND3_GATE U12171 ( .I1(n11681), .I2(n11680), .I3(n11679), .O(n11682) );
  NAND_GATE U12172 ( .I1(n11683), .I2(n11682), .O(n12060) );
  INV_GATE U12173 ( .I1(n12060), .O(n12063) );
  INV_GATE U12174 ( .I1(n11684), .O(n11685) );
  NAND_GATE U12175 ( .I1(n11689), .I2(n11685), .O(n11697) );
  NAND_GATE U12176 ( .I1(n11687), .I2(n11691), .O(n11695) );
  NAND_GATE U12177 ( .I1(n11689), .I2(n11688), .O(n11690) );
  NAND_GATE U12178 ( .I1(n11691), .I2(n11690), .O(n11692) );
  NAND_GATE U12179 ( .I1(n11693), .I2(n11692), .O(n11694) );
  NAND_GATE U12180 ( .I1(n11695), .I2(n11694), .O(n11696) );
  NAND_GATE U12181 ( .I1(n11697), .I2(n11696), .O(n12076) );
  NAND_GATE U12182 ( .I1(n1372), .I2(A[0]), .O(n11698) );
  NAND_GATE U12183 ( .I1(n14781), .I2(n11698), .O(n11699) );
  NAND_GATE U12184 ( .I1(B[9]), .I2(n11699), .O(n11703) );
  NAND_GATE U12185 ( .I1(n1373), .I2(A[1]), .O(n11700) );
  NAND_GATE U12186 ( .I1(n14784), .I2(n11700), .O(n11701) );
  NAND_GATE U12187 ( .I1(B[8]), .I2(n11701), .O(n11702) );
  NAND_GATE U12188 ( .I1(n11703), .I2(n11702), .O(n12088) );
  NAND_GATE U12189 ( .I1(B[7]), .I2(A[2]), .O(n12092) );
  NAND3_GATE U12190 ( .I1(B[7]), .I2(B[8]), .I3(n1196), .O(n12085) );
  NAND_GATE U12191 ( .I1(n12092), .I2(n12085), .O(n11704) );
  NAND_GATE U12192 ( .I1(n12088), .I2(n11704), .O(n11705) );
  INV_GATE U12193 ( .I1(n12092), .O(n12086) );
  INV_GATE U12194 ( .I1(n12085), .O(n12087) );
  NAND_GATE U12195 ( .I1(n12086), .I2(n12087), .O(n12083) );
  NAND_GATE U12196 ( .I1(n11705), .I2(n12083), .O(n12077) );
  NAND_GATE U12197 ( .I1(n12076), .I2(n12077), .O(n11707) );
  NAND_GATE U12198 ( .I1(B[7]), .I2(A[3]), .O(n12078) );
  INV_GATE U12199 ( .I1(n12078), .O(n11706) );
  NAND_GATE U12200 ( .I1(n12076), .I2(n11706), .O(n12073) );
  NAND_GATE U12201 ( .I1(n12077), .I2(n11706), .O(n12072) );
  NAND3_GATE U12202 ( .I1(n11707), .I2(n12073), .I3(n12072), .O(n12062) );
  INV_GATE U12203 ( .I1(n12062), .O(n12059) );
  NAND_GATE U12204 ( .I1(B[7]), .I2(A[4]), .O(n12067) );
  NAND_GATE U12205 ( .I1(n12059), .I2(n12067), .O(n11708) );
  NAND_GATE U12206 ( .I1(n12063), .I2(n11708), .O(n11709) );
  INV_GATE U12207 ( .I1(n12067), .O(n12061) );
  NAND_GATE U12208 ( .I1(n12062), .I2(n12061), .O(n12058) );
  NAND_GATE U12209 ( .I1(n11709), .I2(n12058), .O(n12052) );
  NAND_GATE U12210 ( .I1(n12051), .I2(n12052), .O(n11711) );
  NAND_GATE U12211 ( .I1(B[7]), .I2(A[5]), .O(n12053) );
  INV_GATE U12212 ( .I1(n12053), .O(n11710) );
  NAND_GATE U12213 ( .I1(n12051), .I2(n11710), .O(n12048) );
  NAND_GATE U12214 ( .I1(n12052), .I2(n11710), .O(n12047) );
  NAND3_GATE U12215 ( .I1(n11711), .I2(n12048), .I3(n12047), .O(n12037) );
  INV_GATE U12216 ( .I1(n12037), .O(n12034) );
  NAND_GATE U12217 ( .I1(B[7]), .I2(A[6]), .O(n12042) );
  NAND_GATE U12218 ( .I1(n12034), .I2(n12042), .O(n11712) );
  NAND_GATE U12219 ( .I1(n12038), .I2(n11712), .O(n11713) );
  INV_GATE U12220 ( .I1(n12042), .O(n12036) );
  NAND_GATE U12221 ( .I1(n12037), .I2(n12036), .O(n12033) );
  NAND_GATE U12222 ( .I1(n11713), .I2(n12033), .O(n12027) );
  NAND_GATE U12223 ( .I1(n12026), .I2(n12027), .O(n11715) );
  NAND_GATE U12224 ( .I1(B[7]), .I2(A[7]), .O(n12028) );
  INV_GATE U12225 ( .I1(n12028), .O(n11714) );
  NAND_GATE U12226 ( .I1(n12026), .I2(n11714), .O(n12023) );
  NAND_GATE U12227 ( .I1(n12027), .I2(n11714), .O(n12022) );
  NAND3_GATE U12228 ( .I1(n11715), .I2(n12023), .I3(n12022), .O(n12012) );
  INV_GATE U12229 ( .I1(n12012), .O(n12009) );
  NAND_GATE U12230 ( .I1(B[7]), .I2(A[8]), .O(n12017) );
  NAND_GATE U12231 ( .I1(n12009), .I2(n12017), .O(n11716) );
  NAND_GATE U12232 ( .I1(n12013), .I2(n11716), .O(n11717) );
  INV_GATE U12233 ( .I1(n12017), .O(n12011) );
  NAND_GATE U12234 ( .I1(n12012), .I2(n12011), .O(n12008) );
  NAND_GATE U12235 ( .I1(n11717), .I2(n12008), .O(n12002) );
  NAND_GATE U12236 ( .I1(n12001), .I2(n12002), .O(n11719) );
  NAND_GATE U12237 ( .I1(B[7]), .I2(A[9]), .O(n12003) );
  INV_GATE U12238 ( .I1(n12003), .O(n11718) );
  NAND_GATE U12239 ( .I1(n12001), .I2(n11718), .O(n11998) );
  NAND_GATE U12240 ( .I1(n12002), .I2(n11718), .O(n11997) );
  NAND3_GATE U12241 ( .I1(n11719), .I2(n11998), .I3(n11997), .O(n11987) );
  INV_GATE U12242 ( .I1(n11987), .O(n11984) );
  NAND_GATE U12243 ( .I1(B[7]), .I2(A[10]), .O(n11992) );
  NAND_GATE U12244 ( .I1(n11984), .I2(n11992), .O(n11720) );
  NAND_GATE U12245 ( .I1(n11988), .I2(n11720), .O(n11721) );
  INV_GATE U12246 ( .I1(n11992), .O(n11986) );
  NAND_GATE U12247 ( .I1(n11987), .I2(n11986), .O(n11983) );
  NAND_GATE U12248 ( .I1(n11721), .I2(n11983), .O(n12128) );
  NAND_GATE U12249 ( .I1(n12127), .I2(n12128), .O(n11723) );
  NAND_GATE U12250 ( .I1(B[7]), .I2(A[11]), .O(n12129) );
  INV_GATE U12251 ( .I1(n12129), .O(n11722) );
  NAND_GATE U12252 ( .I1(n12128), .I2(n11722), .O(n12124) );
  NAND_GATE U12253 ( .I1(n12127), .I2(n11722), .O(n12123) );
  NAND3_GATE U12254 ( .I1(n11723), .I2(n12124), .I3(n12123), .O(n11976) );
  NAND_GATE U12255 ( .I1(B[7]), .I2(A[12]), .O(n11978) );
  OR_GATE U12256 ( .I1(n11724), .I2(n11729), .O(n11727) );
  OR_GATE U12257 ( .I1(n11725), .I2(n11728), .O(n11726) );
  AND_GATE U12258 ( .I1(n11727), .I2(n11726), .O(n11734) );
  NAND_GATE U12259 ( .I1(n11728), .I2(n968), .O(n11732) );
  NAND3_GATE U12260 ( .I1(n11732), .I2(n11731), .I3(n11730), .O(n11733) );
  NAND_GATE U12261 ( .I1(n11734), .I2(n11733), .O(n11973) );
  NAND_GATE U12262 ( .I1(n11978), .I2(n11973), .O(n11735) );
  NAND_GATE U12263 ( .I1(n11976), .I2(n11735), .O(n11736) );
  INV_GATE U12264 ( .I1(n11978), .O(n11975) );
  NAND_GATE U12265 ( .I1(n11975), .I2(n40), .O(n11971) );
  NAND_GATE U12266 ( .I1(n11736), .I2(n11971), .O(n12142) );
  NAND_GATE U12267 ( .I1(n12141), .I2(n12142), .O(n11738) );
  NAND_GATE U12268 ( .I1(B[7]), .I2(A[13]), .O(n12143) );
  INV_GATE U12269 ( .I1(n12143), .O(n11737) );
  NAND_GATE U12270 ( .I1(n12142), .I2(n11737), .O(n12138) );
  NAND_GATE U12271 ( .I1(n12141), .I2(n11737), .O(n12137) );
  NAND3_GATE U12272 ( .I1(n11738), .I2(n12138), .I3(n12137), .O(n11964) );
  NAND_GATE U12273 ( .I1(B[7]), .I2(A[14]), .O(n11966) );
  OR_GATE U12274 ( .I1(n11740), .I2(n11744), .O(n11741) );
  AND_GATE U12275 ( .I1(n11742), .I2(n11741), .O(n11750) );
  INV_GATE U12276 ( .I1(n11745), .O(n11743) );
  NAND_GATE U12277 ( .I1(n11744), .I2(n11743), .O(n11748) );
  NAND_GATE U12278 ( .I1(n1286), .I2(n11745), .O(n11747) );
  NAND3_GATE U12279 ( .I1(n11748), .I2(n11747), .I3(n11746), .O(n11749) );
  NAND_GATE U12280 ( .I1(n11750), .I2(n11749), .O(n11961) );
  NAND_GATE U12281 ( .I1(n11966), .I2(n11961), .O(n11751) );
  NAND_GATE U12282 ( .I1(n11964), .I2(n11751), .O(n11752) );
  INV_GATE U12283 ( .I1(n11966), .O(n11962) );
  INV_GATE U12284 ( .I1(n11961), .O(n11963) );
  NAND_GATE U12285 ( .I1(n11962), .I2(n11963), .O(n11960) );
  NAND_GATE U12286 ( .I1(n11752), .I2(n11960), .O(n12157) );
  NAND_GATE U12287 ( .I1(n12156), .I2(n12157), .O(n11754) );
  NAND_GATE U12288 ( .I1(B[7]), .I2(A[15]), .O(n12158) );
  INV_GATE U12289 ( .I1(n12158), .O(n11753) );
  NAND_GATE U12290 ( .I1(n12157), .I2(n11753), .O(n12153) );
  NAND_GATE U12291 ( .I1(n11950), .I2(n11955), .O(n11755) );
  NAND_GATE U12292 ( .I1(n11952), .I2(n11755), .O(n11756) );
  NAND_GATE U12293 ( .I1(n11948), .I2(n11756), .O(n11942) );
  NAND3_GATE U12294 ( .I1(n11939), .I2(n11940), .I3(n11942), .O(n11758) );
  NAND_GATE U12295 ( .I1(n11757), .I2(n11942), .O(n11935) );
  NAND3_GATE U12296 ( .I1(n11934), .I2(n11758), .I3(n11935), .O(n12173) );
  NAND_GATE U12297 ( .I1(n12172), .I2(n12177), .O(n11759) );
  NAND_GATE U12298 ( .I1(n12173), .I2(n11759), .O(n11760) );
  NAND_GATE U12299 ( .I1(n12169), .I2(n11760), .O(n11928) );
  NAND_GATE U12300 ( .I1(n11774), .I2(n11928), .O(n11924) );
  INV_GATE U12301 ( .I1(n11761), .O(n11762) );
  NAND_GATE U12302 ( .I1(n11762), .I2(n11768), .O(n11773) );
  NAND_GATE U12303 ( .I1(n11767), .I2(n11766), .O(n11763) );
  NAND_GATE U12304 ( .I1(n11764), .I2(n11763), .O(n11771) );
  NAND3_GATE U12305 ( .I1(n11767), .I2(n11766), .I3(n11765), .O(n11770) );
  NAND_GATE U12306 ( .I1(n233), .I2(n11768), .O(n11769) );
  NAND3_GATE U12307 ( .I1(n11771), .I2(n11770), .I3(n11769), .O(n11772) );
  NAND_GATE U12308 ( .I1(n11773), .I2(n11772), .O(n11927) );
  NAND_GATE U12309 ( .I1(n11928), .I2(n11927), .O(n11775) );
  NAND_GATE U12310 ( .I1(n11774), .I2(n11927), .O(n11923) );
  NAND3_GATE U12311 ( .I1(n11924), .I2(n11775), .I3(n11923), .O(n12190) );
  NAND_GATE U12312 ( .I1(n12189), .I2(n12194), .O(n11776) );
  NAND_GATE U12313 ( .I1(n12190), .I2(n11776), .O(n11777) );
  NAND_GATE U12314 ( .I1(n12186), .I2(n11777), .O(n11918) );
  NAND_GATE U12315 ( .I1(n11791), .I2(n11918), .O(n11914) );
  NAND_GATE U12316 ( .I1(n11779), .I2(n11778), .O(n11785) );
  NAND_GATE U12317 ( .I1(n1202), .I2(n11787), .O(n11781) );
  NAND_GATE U12318 ( .I1(n11778), .I2(n11781), .O(n11782) );
  NAND_GATE U12319 ( .I1(n11783), .I2(n11782), .O(n11784) );
  NAND_GATE U12320 ( .I1(n11785), .I2(n11784), .O(n11790) );
  INV_GATE U12321 ( .I1(n11786), .O(n11788) );
  NAND_GATE U12322 ( .I1(n11788), .I2(n11787), .O(n11789) );
  NAND_GATE U12323 ( .I1(n11790), .I2(n11789), .O(n11917) );
  NAND_GATE U12324 ( .I1(n11918), .I2(n11917), .O(n11792) );
  NAND_GATE U12325 ( .I1(n11791), .I2(n11917), .O(n11913) );
  NAND3_GATE U12326 ( .I1(n11914), .I2(n11792), .I3(n11913), .O(n12209) );
  NAND_GATE U12327 ( .I1(n12208), .I2(n12211), .O(n11793) );
  NAND_GATE U12328 ( .I1(n12209), .I2(n11793), .O(n11794) );
  NAND_GATE U12329 ( .I1(n12203), .I2(n11794), .O(n11906) );
  NAND_GATE U12330 ( .I1(n11808), .I2(n11906), .O(n11908) );
  INV_GATE U12331 ( .I1(n11804), .O(n11798) );
  NAND_GATE U12332 ( .I1(n11799), .I2(n11798), .O(n11795) );
  NAND_GATE U12333 ( .I1(n11796), .I2(n11795), .O(n11802) );
  NAND_GATE U12334 ( .I1(n11802), .I2(n11801), .O(n11807) );
  INV_GATE U12335 ( .I1(n11803), .O(n11805) );
  NAND_GATE U12336 ( .I1(n11805), .I2(n11804), .O(n11806) );
  NAND_GATE U12337 ( .I1(n11807), .I2(n11806), .O(n11909) );
  NAND_GATE U12338 ( .I1(n11906), .I2(n11909), .O(n11809) );
  NAND_GATE U12339 ( .I1(n11808), .I2(n11909), .O(n11907) );
  NAND3_GATE U12340 ( .I1(n11908), .I2(n11809), .I3(n11907), .O(n11900) );
  NAND_GATE U12341 ( .I1(n11894), .I2(n11895), .O(n11810) );
  NAND_GATE U12342 ( .I1(n11900), .I2(n11810), .O(n11811) );
  NAND_GATE U12343 ( .I1(n11899), .I2(n11811), .O(n11883) );
  NAND_GATE U12344 ( .I1(n11885), .I2(n11883), .O(n11813) );
  NAND_GATE U12345 ( .I1(n11812), .I2(n11883), .O(n11880) );
  NAND_GATE U12346 ( .I1(n12332), .I2(n11874), .O(n11814) );
  NAND_GATE U12347 ( .I1(n11875), .I2(n11814), .O(n11815) );
  NAND_GATE U12348 ( .I1(n11816), .I2(n11815), .O(n11869) );
  NAND_GATE U12349 ( .I1(n11006), .I2(n11826), .O(n11817) );
  NAND_GATE U12350 ( .I1(n11823), .I2(n11817), .O(n11821) );
  INV_GATE U12351 ( .I1(n11823), .O(n11818) );
  NAND3_GATE U12352 ( .I1(n11006), .I2(n11818), .I3(n11826), .O(n11820) );
  NAND3_GATE U12353 ( .I1(n11821), .I2(n11820), .I3(n11819), .O(n11833) );
  OR_GATE U12354 ( .I1(n11823), .I2(n11822), .O(n11832) );
  NAND_GATE U12355 ( .I1(n11825), .I2(n11824), .O(n11826) );
  NAND_GATE U12356 ( .I1(n241), .I2(n11826), .O(n11830) );
  INV_GATE U12357 ( .I1(n11827), .O(n11829) );
  NAND3_GATE U12358 ( .I1(n11830), .I2(n11829), .I3(n11828), .O(n11831) );
  AND_GATE U12359 ( .I1(n11832), .I2(n11831), .O(n11834) );
  NAND3_GATE U12360 ( .I1(n11869), .I2(n11833), .I3(n11834), .O(n11836) );
  NAND_GATE U12361 ( .I1(B[7]), .I2(A[27]), .O(n11861) );
  INV_GATE U12362 ( .I1(n11861), .O(n11864) );
  NAND_GATE U12363 ( .I1(n11864), .I2(n11869), .O(n11835) );
  NAND3_GATE U12364 ( .I1(n11836), .I2(n11835), .I3(n11868), .O(n12296) );
  NAND4_GATE U12365 ( .I1(n11838), .I2(n11837), .I3(n12296), .I4(n11855), .O(
        n11840) );
  NAND_GATE U12366 ( .I1(n11856), .I2(n12296), .O(n11839) );
  NAND3_GATE U12367 ( .I1(n11857), .I2(n11840), .I3(n11839), .O(n12243) );
  NAND_GATE U12368 ( .I1(n12238), .I2(n12236), .O(n11841) );
  NAND_GATE U12369 ( .I1(n12243), .I2(n11841), .O(n11842) );
  NAND_GATE U12370 ( .I1(n12242), .I2(n11842), .O(n12267) );
  NAND_GATE U12371 ( .I1(n12271), .I2(n12268), .O(n11843) );
  NAND_GATE U12372 ( .I1(n12267), .I2(n11843), .O(n11844) );
  NAND_GATE U12373 ( .I1(n11845), .I2(n11844), .O(n11854) );
  NAND_GATE U12374 ( .I1(n15351), .I2(n11852), .O(n11846) );
  NAND_GATE U12375 ( .I1(n11854), .I2(n11846), .O(n11847) );
  NAND_GATE U12376 ( .I1(n11849), .I2(n479), .O(n11850) );
  AND_GATE U12377 ( .I1(n11851), .I2(n11850), .O(\A1[37] ) );
  NAND_GATE U12378 ( .I1(n11852), .I2(n622), .O(n15350) );
  NAND3_GATE U12379 ( .I1(n15350), .I2(n15354), .I3(n1220), .O(n12256) );
  NAND_GATE U12380 ( .I1(B[6]), .I2(A[31]), .O(n12279) );
  INV_GATE U12381 ( .I1(n12279), .O(n12260) );
  NAND_GATE U12382 ( .I1(B[6]), .I2(A[30]), .O(n12285) );
  INV_GATE U12383 ( .I1(n12285), .O(n12286) );
  NAND_GATE U12384 ( .I1(B[6]), .I2(A[29]), .O(n12315) );
  INV_GATE U12385 ( .I1(n12315), .O(n12302) );
  NAND_GATE U12386 ( .I1(n915), .I2(n11855), .O(n12294) );
  NAND_GATE U12387 ( .I1(n11856), .I2(n11858), .O(n12297) );
  INV_GATE U12388 ( .I1(n12294), .O(n12295) );
  NAND_GATE U12389 ( .I1(n12296), .I2(n12295), .O(n11859) );
  NAND_GATE U12390 ( .I1(n12293), .I2(n12294), .O(n11858) );
  NAND_GATE U12391 ( .I1(n11859), .I2(n11858), .O(n11860) );
  NAND_GATE U12392 ( .I1(n12292), .I2(n11860), .O(n12307) );
  NAND_GATE U12393 ( .I1(n918), .I2(n12307), .O(n12230) );
  NAND_GATE U12394 ( .I1(n1300), .I2(n11869), .O(n11867) );
  NAND3_GATE U12395 ( .I1(n11861), .I2(n11862), .I3(n666), .O(n11866) );
  NAND_GATE U12396 ( .I1(n666), .I2(n11862), .O(n11863) );
  NAND_GATE U12397 ( .I1(n11864), .I2(n11863), .O(n11865) );
  NAND3_GATE U12398 ( .I1(n11867), .I2(n11866), .I3(n11865), .O(n11872) );
  INV_GATE U12399 ( .I1(n11868), .O(n11870) );
  NAND_GATE U12400 ( .I1(n11870), .I2(n11869), .O(n11871) );
  NAND_GATE U12401 ( .I1(n11872), .I2(n11871), .O(n12321) );
  NAND_GATE U12402 ( .I1(B[6]), .I2(A[27]), .O(n12701) );
  INV_GATE U12403 ( .I1(n12701), .O(n12223) );
  NAND_GATE U12404 ( .I1(n11873), .I2(n11878), .O(n12327) );
  INV_GATE U12405 ( .I1(n12327), .O(n12330) );
  NAND3_GATE U12406 ( .I1(n11873), .I2(n11875), .I3(n11876), .O(n12329) );
  NAND_GATE U12407 ( .I1(n11874), .I2(n187), .O(n11878) );
  NAND_GATE U12408 ( .I1(n11876), .I2(n11875), .O(n11877) );
  NAND_GATE U12409 ( .I1(n11878), .I2(n11877), .O(n12331) );
  NAND3_GATE U12410 ( .I1(n12223), .I2(n12335), .I3(n12326), .O(n12325) );
  OR_GATE U12411 ( .I1(n11883), .I2(n11879), .O(n11882) );
  OR_GATE U12412 ( .I1(n11880), .I2(n11885), .O(n11881) );
  AND_GATE U12413 ( .I1(n11882), .I2(n11881), .O(n11890) );
  NAND_GATE U12414 ( .I1(n1239), .I2(n11883), .O(n11887) );
  INV_GATE U12415 ( .I1(n11883), .O(n11884) );
  NAND_GATE U12416 ( .I1(n11885), .I2(n11884), .O(n11886) );
  NAND3_GATE U12417 ( .I1(n11888), .I2(n11887), .I3(n11886), .O(n11889) );
  NAND_GATE U12418 ( .I1(n11890), .I2(n11889), .O(n12342) );
  INV_GATE U12419 ( .I1(n12342), .O(n12340) );
  NAND_GATE U12420 ( .I1(B[6]), .I2(A[26]), .O(n12338) );
  INV_GATE U12421 ( .I1(n12338), .O(n12344) );
  NAND_GATE U12422 ( .I1(n12340), .I2(n12344), .O(n12337) );
  NAND_GATE U12423 ( .I1(n11895), .I2(n591), .O(n11891) );
  NAND_GATE U12424 ( .I1(n11892), .I2(n11891), .O(n11898) );
  NAND_GATE U12425 ( .I1(n11893), .I2(n11900), .O(n11897) );
  NAND3_GATE U12426 ( .I1(n11895), .I2(n591), .I3(n11894), .O(n11896) );
  NAND3_GATE U12427 ( .I1(n11898), .I2(n11897), .I3(n11896), .O(n11902) );
  NAND_GATE U12428 ( .I1(n190), .I2(n11900), .O(n11901) );
  NAND_GATE U12429 ( .I1(n11902), .I2(n11901), .O(n12354) );
  NAND_GATE U12430 ( .I1(n922), .I2(n11909), .O(n11904) );
  NAND3_GATE U12431 ( .I1(n11905), .I2(n11904), .I3(n11903), .O(n11912) );
  OR_GATE U12432 ( .I1(n11907), .I2(n11906), .O(n11911) );
  OR_GATE U12433 ( .I1(n11909), .I2(n11908), .O(n11910) );
  NAND3_GATE U12434 ( .I1(n11912), .I2(n11911), .I3(n11910), .O(n12366) );
  INV_GATE U12435 ( .I1(n12366), .O(n12362) );
  NAND_GATE U12436 ( .I1(B[6]), .I2(A[24]), .O(n12365) );
  INV_GATE U12437 ( .I1(n12365), .O(n12360) );
  NAND_GATE U12438 ( .I1(n12362), .I2(n12360), .O(n12358) );
  NAND_GATE U12439 ( .I1(B[6]), .I2(A[23]), .O(n12375) );
  INV_GATE U12440 ( .I1(n12375), .O(n12368) );
  NAND_GATE U12441 ( .I1(B[6]), .I2(A[22]), .O(n12681) );
  OR_GATE U12442 ( .I1(n11913), .I2(n11918), .O(n11916) );
  OR_GATE U12443 ( .I1(n11917), .I2(n11914), .O(n11915) );
  NAND_GATE U12444 ( .I1(n232), .I2(n11917), .O(n11920) );
  NAND3_GATE U12445 ( .I1(n11921), .I2(n11920), .I3(n11919), .O(n11922) );
  INV_GATE U12446 ( .I1(n12680), .O(n12678) );
  NAND_GATE U12447 ( .I1(n339), .I2(n12678), .O(n12684) );
  NAND_GATE U12448 ( .I1(B[6]), .I2(A[21]), .O(n12388) );
  INV_GATE U12449 ( .I1(n12388), .O(n12199) );
  OR_GATE U12450 ( .I1(n11923), .I2(n11928), .O(n11926) );
  OR_GATE U12451 ( .I1(n11927), .I2(n11924), .O(n11925) );
  AND_GATE U12452 ( .I1(n11926), .I2(n11925), .O(n11933) );
  NAND_GATE U12453 ( .I1(n956), .I2(n11927), .O(n11931) );
  NAND3_GATE U12454 ( .I1(n11931), .I2(n11930), .I3(n11929), .O(n11932) );
  NAND_GATE U12455 ( .I1(n11933), .I2(n11932), .O(n12664) );
  NAND_GATE U12456 ( .I1(B[6]), .I2(A[20]), .O(n12669) );
  INV_GATE U12457 ( .I1(n12669), .O(n12663) );
  NAND_GATE U12458 ( .I1(n625), .I2(n12663), .O(n12661) );
  NAND_GATE U12459 ( .I1(B[6]), .I2(A[19]), .O(n12399) );
  INV_GATE U12460 ( .I1(n12399), .O(n12182) );
  OR_GATE U12461 ( .I1(n11934), .I2(n11942), .O(n11937) );
  OR_GATE U12462 ( .I1(n11938), .I2(n11935), .O(n11936) );
  AND_GATE U12463 ( .I1(n11937), .I2(n11936), .O(n11947) );
  NAND_GATE U12464 ( .I1(n113), .I2(n11938), .O(n11945) );
  NAND_GATE U12465 ( .I1(n11940), .I2(n11939), .O(n11941) );
  NAND_GATE U12466 ( .I1(n11942), .I2(n11941), .O(n11944) );
  NAND3_GATE U12467 ( .I1(n11945), .I2(n11944), .I3(n11943), .O(n11946) );
  NAND_GATE U12468 ( .I1(B[6]), .I2(A[18]), .O(n12411) );
  INV_GATE U12469 ( .I1(n12411), .O(n12407) );
  NAND_GATE U12470 ( .I1(n629), .I2(n12407), .O(n12404) );
  INV_GATE U12471 ( .I1(n11948), .O(n11949) );
  NAND_GATE U12472 ( .I1(n11949), .I2(n11952), .O(n11959) );
  NAND_GATE U12473 ( .I1(n11950), .I2(n686), .O(n11954) );
  NAND_GATE U12474 ( .I1(n11951), .I2(n11954), .O(n11957) );
  NAND_GATE U12475 ( .I1(n11957), .I2(n11956), .O(n11958) );
  NAND_GATE U12476 ( .I1(n11959), .I2(n11958), .O(n12648) );
  NAND_GATE U12477 ( .I1(n11962), .I2(n11965), .O(n11968) );
  NAND_GATE U12478 ( .I1(n11968), .I2(n11967), .O(n11969) );
  NAND_GATE U12479 ( .I1(n11970), .I2(n11969), .O(n12633) );
  INV_GATE U12480 ( .I1(n11971), .O(n11972) );
  NAND_GATE U12481 ( .I1(n11976), .I2(n11972), .O(n11982) );
  INV_GATE U12482 ( .I1(n11976), .O(n11974) );
  NAND_GATE U12483 ( .I1(n11974), .I2(n11973), .O(n11977) );
  NAND_GATE U12484 ( .I1(n11975), .I2(n11977), .O(n11980) );
  NAND_GATE U12485 ( .I1(n11980), .I2(n11979), .O(n11981) );
  NAND_GATE U12486 ( .I1(n11982), .I2(n11981), .O(n12617) );
  OR_GATE U12487 ( .I1(n11983), .I2(n11985), .O(n11996) );
  NAND_GATE U12488 ( .I1(n11985), .I2(n11984), .O(n11990) );
  NAND_GATE U12489 ( .I1(n11986), .I2(n11990), .O(n11994) );
  NAND_GATE U12490 ( .I1(n11988), .I2(n11987), .O(n11989) );
  NAND_GATE U12491 ( .I1(n11990), .I2(n11989), .O(n11991) );
  NAND_GATE U12492 ( .I1(n11992), .I2(n11991), .O(n11993) );
  NAND_GATE U12493 ( .I1(n11994), .I2(n11993), .O(n11995) );
  NAND_GATE U12494 ( .I1(n11996), .I2(n11995), .O(n12602) );
  OR_GATE U12495 ( .I1(n11997), .I2(n12001), .O(n12000) );
  OR_GATE U12496 ( .I1(n11998), .I2(n12002), .O(n11999) );
  AND_GATE U12497 ( .I1(n12000), .I2(n11999), .O(n12007) );
  NAND_GATE U12498 ( .I1(n12001), .I2(n1010), .O(n12005) );
  NAND3_GATE U12499 ( .I1(n12005), .I2(n12004), .I3(n12003), .O(n12006) );
  NAND_GATE U12500 ( .I1(n12007), .I2(n12006), .O(n12460) );
  INV_GATE U12501 ( .I1(n12460), .O(n12463) );
  OR_GATE U12502 ( .I1(n12008), .I2(n12010), .O(n12021) );
  NAND_GATE U12503 ( .I1(n12010), .I2(n12009), .O(n12015) );
  NAND_GATE U12504 ( .I1(n12011), .I2(n12015), .O(n12019) );
  NAND_GATE U12505 ( .I1(n12013), .I2(n12012), .O(n12014) );
  NAND_GATE U12506 ( .I1(n12015), .I2(n12014), .O(n12016) );
  NAND_GATE U12507 ( .I1(n12017), .I2(n12016), .O(n12018) );
  NAND_GATE U12508 ( .I1(n12019), .I2(n12018), .O(n12020) );
  NAND_GATE U12509 ( .I1(n12021), .I2(n12020), .O(n12476) );
  OR_GATE U12510 ( .I1(n12022), .I2(n12026), .O(n12025) );
  OR_GATE U12511 ( .I1(n12023), .I2(n12027), .O(n12024) );
  AND_GATE U12512 ( .I1(n12025), .I2(n12024), .O(n12032) );
  NAND_GATE U12513 ( .I1(n12026), .I2(n1018), .O(n12030) );
  NAND3_GATE U12514 ( .I1(n12030), .I2(n12029), .I3(n12028), .O(n12031) );
  NAND_GATE U12515 ( .I1(n12032), .I2(n12031), .O(n12485) );
  INV_GATE U12516 ( .I1(n12485), .O(n12488) );
  OR_GATE U12517 ( .I1(n12033), .I2(n12035), .O(n12046) );
  NAND_GATE U12518 ( .I1(n12035), .I2(n12034), .O(n12040) );
  NAND_GATE U12519 ( .I1(n12036), .I2(n12040), .O(n12044) );
  NAND_GATE U12520 ( .I1(n12038), .I2(n12037), .O(n12039) );
  NAND_GATE U12521 ( .I1(n12040), .I2(n12039), .O(n12041) );
  NAND_GATE U12522 ( .I1(n12042), .I2(n12041), .O(n12043) );
  NAND_GATE U12523 ( .I1(n12044), .I2(n12043), .O(n12045) );
  NAND_GATE U12524 ( .I1(n12046), .I2(n12045), .O(n12501) );
  OR_GATE U12525 ( .I1(n12047), .I2(n12051), .O(n12050) );
  OR_GATE U12526 ( .I1(n12048), .I2(n12052), .O(n12049) );
  AND_GATE U12527 ( .I1(n12050), .I2(n12049), .O(n12057) );
  NAND_GATE U12528 ( .I1(n12051), .I2(n1113), .O(n12055) );
  NAND3_GATE U12529 ( .I1(n12055), .I2(n12054), .I3(n12053), .O(n12056) );
  NAND_GATE U12530 ( .I1(n12057), .I2(n12056), .O(n12510) );
  INV_GATE U12531 ( .I1(n12510), .O(n12513) );
  OR_GATE U12532 ( .I1(n12058), .I2(n12060), .O(n12071) );
  NAND_GATE U12533 ( .I1(n12060), .I2(n12059), .O(n12065) );
  NAND_GATE U12534 ( .I1(n12061), .I2(n12065), .O(n12069) );
  NAND_GATE U12535 ( .I1(n12063), .I2(n12062), .O(n12064) );
  NAND_GATE U12536 ( .I1(n12065), .I2(n12064), .O(n12066) );
  NAND_GATE U12537 ( .I1(n12067), .I2(n12066), .O(n12068) );
  NAND_GATE U12538 ( .I1(n12069), .I2(n12068), .O(n12070) );
  NAND_GATE U12539 ( .I1(n12071), .I2(n12070), .O(n12526) );
  OR_GATE U12540 ( .I1(n12072), .I2(n12076), .O(n12075) );
  OR_GATE U12541 ( .I1(n12073), .I2(n12077), .O(n12074) );
  AND_GATE U12542 ( .I1(n12075), .I2(n12074), .O(n12082) );
  NAND_GATE U12543 ( .I1(n12076), .I2(n1185), .O(n12080) );
  NAND3_GATE U12544 ( .I1(n12080), .I2(n12079), .I3(n12078), .O(n12081) );
  NAND_GATE U12545 ( .I1(n12082), .I2(n12081), .O(n12535) );
  INV_GATE U12546 ( .I1(n12535), .O(n12538) );
  INV_GATE U12547 ( .I1(n12083), .O(n12084) );
  NAND_GATE U12548 ( .I1(n12088), .I2(n12084), .O(n12096) );
  NAND_GATE U12549 ( .I1(n12086), .I2(n12090), .O(n12094) );
  NAND_GATE U12550 ( .I1(n12088), .I2(n12087), .O(n12089) );
  NAND_GATE U12551 ( .I1(n12090), .I2(n12089), .O(n12091) );
  NAND_GATE U12552 ( .I1(n12092), .I2(n12091), .O(n12093) );
  NAND_GATE U12553 ( .I1(n12094), .I2(n12093), .O(n12095) );
  NAND_GATE U12554 ( .I1(n12096), .I2(n12095), .O(n12551) );
  NAND_GATE U12555 ( .I1(n1371), .I2(A[0]), .O(n12097) );
  NAND_GATE U12556 ( .I1(n14781), .I2(n12097), .O(n12098) );
  NAND_GATE U12557 ( .I1(B[8]), .I2(n12098), .O(n12102) );
  NAND_GATE U12558 ( .I1(n1372), .I2(A[1]), .O(n12099) );
  NAND_GATE U12559 ( .I1(n14784), .I2(n12099), .O(n12100) );
  NAND_GATE U12560 ( .I1(B[7]), .I2(n12100), .O(n12101) );
  NAND_GATE U12561 ( .I1(n12102), .I2(n12101), .O(n12563) );
  NAND_GATE U12562 ( .I1(B[6]), .I2(A[2]), .O(n12567) );
  NAND3_GATE U12563 ( .I1(B[6]), .I2(B[7]), .I3(n1196), .O(n12560) );
  NAND_GATE U12564 ( .I1(n12567), .I2(n12560), .O(n12103) );
  NAND_GATE U12565 ( .I1(n12563), .I2(n12103), .O(n12104) );
  INV_GATE U12566 ( .I1(n12567), .O(n12561) );
  INV_GATE U12567 ( .I1(n12560), .O(n12562) );
  NAND_GATE U12568 ( .I1(n12561), .I2(n12562), .O(n12558) );
  NAND_GATE U12569 ( .I1(n12104), .I2(n12558), .O(n12552) );
  NAND_GATE U12570 ( .I1(n12551), .I2(n12552), .O(n12106) );
  NAND_GATE U12571 ( .I1(B[6]), .I2(A[3]), .O(n12553) );
  INV_GATE U12572 ( .I1(n12553), .O(n12105) );
  NAND_GATE U12573 ( .I1(n12551), .I2(n12105), .O(n12548) );
  NAND_GATE U12574 ( .I1(n12552), .I2(n12105), .O(n12547) );
  NAND3_GATE U12575 ( .I1(n12106), .I2(n12548), .I3(n12547), .O(n12537) );
  INV_GATE U12576 ( .I1(n12537), .O(n12534) );
  NAND_GATE U12577 ( .I1(B[6]), .I2(A[4]), .O(n12542) );
  NAND_GATE U12578 ( .I1(n12534), .I2(n12542), .O(n12107) );
  NAND_GATE U12579 ( .I1(n12538), .I2(n12107), .O(n12108) );
  INV_GATE U12580 ( .I1(n12542), .O(n12536) );
  NAND_GATE U12581 ( .I1(n12537), .I2(n12536), .O(n12533) );
  NAND_GATE U12582 ( .I1(n12108), .I2(n12533), .O(n12527) );
  NAND_GATE U12583 ( .I1(n12526), .I2(n12527), .O(n12110) );
  NAND_GATE U12584 ( .I1(B[6]), .I2(A[5]), .O(n12528) );
  INV_GATE U12585 ( .I1(n12528), .O(n12109) );
  NAND_GATE U12586 ( .I1(n12526), .I2(n12109), .O(n12523) );
  NAND_GATE U12587 ( .I1(n12527), .I2(n12109), .O(n12522) );
  NAND3_GATE U12588 ( .I1(n12110), .I2(n12523), .I3(n12522), .O(n12512) );
  INV_GATE U12589 ( .I1(n12512), .O(n12509) );
  NAND_GATE U12590 ( .I1(B[6]), .I2(A[6]), .O(n12517) );
  NAND_GATE U12591 ( .I1(n12509), .I2(n12517), .O(n12111) );
  NAND_GATE U12592 ( .I1(n12513), .I2(n12111), .O(n12112) );
  INV_GATE U12593 ( .I1(n12517), .O(n12511) );
  NAND_GATE U12594 ( .I1(n12512), .I2(n12511), .O(n12508) );
  NAND_GATE U12595 ( .I1(n12112), .I2(n12508), .O(n12502) );
  NAND_GATE U12596 ( .I1(n12501), .I2(n12502), .O(n12114) );
  NAND_GATE U12597 ( .I1(B[6]), .I2(A[7]), .O(n12503) );
  INV_GATE U12598 ( .I1(n12503), .O(n12113) );
  NAND_GATE U12599 ( .I1(n12501), .I2(n12113), .O(n12498) );
  NAND_GATE U12600 ( .I1(n12502), .I2(n12113), .O(n12497) );
  NAND3_GATE U12601 ( .I1(n12114), .I2(n12498), .I3(n12497), .O(n12487) );
  INV_GATE U12602 ( .I1(n12487), .O(n12484) );
  NAND_GATE U12603 ( .I1(B[6]), .I2(A[8]), .O(n12492) );
  NAND_GATE U12604 ( .I1(n12484), .I2(n12492), .O(n12115) );
  NAND_GATE U12605 ( .I1(n12488), .I2(n12115), .O(n12116) );
  INV_GATE U12606 ( .I1(n12492), .O(n12486) );
  NAND_GATE U12607 ( .I1(n12487), .I2(n12486), .O(n12483) );
  NAND_GATE U12608 ( .I1(n12116), .I2(n12483), .O(n12477) );
  NAND_GATE U12609 ( .I1(n12476), .I2(n12477), .O(n12118) );
  NAND_GATE U12610 ( .I1(B[6]), .I2(A[9]), .O(n12478) );
  INV_GATE U12611 ( .I1(n12478), .O(n12117) );
  NAND_GATE U12612 ( .I1(n12476), .I2(n12117), .O(n12473) );
  NAND_GATE U12613 ( .I1(n12477), .I2(n12117), .O(n12472) );
  NAND3_GATE U12614 ( .I1(n12118), .I2(n12473), .I3(n12472), .O(n12462) );
  INV_GATE U12615 ( .I1(n12462), .O(n12459) );
  NAND_GATE U12616 ( .I1(B[6]), .I2(A[10]), .O(n12467) );
  NAND_GATE U12617 ( .I1(n12459), .I2(n12467), .O(n12119) );
  NAND_GATE U12618 ( .I1(n12463), .I2(n12119), .O(n12120) );
  INV_GATE U12619 ( .I1(n12467), .O(n12461) );
  NAND_GATE U12620 ( .I1(n12462), .I2(n12461), .O(n12458) );
  NAND_GATE U12621 ( .I1(n12120), .I2(n12458), .O(n12603) );
  NAND_GATE U12622 ( .I1(n12602), .I2(n12603), .O(n12122) );
  NAND_GATE U12623 ( .I1(B[6]), .I2(A[11]), .O(n12604) );
  INV_GATE U12624 ( .I1(n12604), .O(n12121) );
  NAND_GATE U12625 ( .I1(n12603), .I2(n12121), .O(n12599) );
  NAND_GATE U12626 ( .I1(n12602), .I2(n12121), .O(n12598) );
  NAND3_GATE U12627 ( .I1(n12122), .I2(n12599), .I3(n12598), .O(n12449) );
  NAND_GATE U12628 ( .I1(B[6]), .I2(A[12]), .O(n12453) );
  OR_GATE U12629 ( .I1(n12123), .I2(n12128), .O(n12126) );
  OR_GATE U12630 ( .I1(n12124), .I2(n12127), .O(n12125) );
  NAND_GATE U12631 ( .I1(n12127), .I2(n996), .O(n12131) );
  NAND3_GATE U12632 ( .I1(n12131), .I2(n12130), .I3(n12129), .O(n12132) );
  NAND_GATE U12633 ( .I1(n12453), .I2(n12445), .O(n12133) );
  NAND_GATE U12634 ( .I1(n12449), .I2(n12133), .O(n12134) );
  INV_GATE U12635 ( .I1(n12453), .O(n12447) );
  INV_GATE U12636 ( .I1(n12445), .O(n12448) );
  NAND_GATE U12637 ( .I1(n12447), .I2(n12448), .O(n12443) );
  NAND_GATE U12638 ( .I1(n12134), .I2(n12443), .O(n12618) );
  NAND_GATE U12639 ( .I1(n12617), .I2(n12618), .O(n12136) );
  NAND_GATE U12640 ( .I1(B[6]), .I2(A[13]), .O(n12619) );
  INV_GATE U12641 ( .I1(n12619), .O(n12135) );
  NAND_GATE U12642 ( .I1(n12618), .I2(n12135), .O(n12614) );
  NAND_GATE U12643 ( .I1(n12617), .I2(n12135), .O(n12613) );
  NAND3_GATE U12644 ( .I1(n12136), .I2(n12614), .I3(n12613), .O(n12434) );
  NAND_GATE U12645 ( .I1(B[6]), .I2(A[14]), .O(n12438) );
  OR_GATE U12646 ( .I1(n12137), .I2(n12142), .O(n12140) );
  OR_GATE U12647 ( .I1(n12138), .I2(n12141), .O(n12139) );
  AND_GATE U12648 ( .I1(n12140), .I2(n12139), .O(n12147) );
  NAND_GATE U12649 ( .I1(n12141), .I2(n935), .O(n12145) );
  NAND3_GATE U12650 ( .I1(n12145), .I2(n12144), .I3(n12143), .O(n12146) );
  NAND_GATE U12651 ( .I1(n12147), .I2(n12146), .O(n12430) );
  NAND_GATE U12652 ( .I1(n12438), .I2(n12430), .O(n12148) );
  NAND_GATE U12653 ( .I1(n12434), .I2(n12148), .O(n12149) );
  INV_GATE U12654 ( .I1(n12438), .O(n12432) );
  INV_GATE U12655 ( .I1(n12430), .O(n12433) );
  NAND_GATE U12656 ( .I1(n12432), .I2(n12433), .O(n12428) );
  NAND_GATE U12657 ( .I1(n12149), .I2(n12428), .O(n12634) );
  NAND_GATE U12658 ( .I1(n12633), .I2(n12634), .O(n12151) );
  NAND_GATE U12659 ( .I1(B[6]), .I2(A[15]), .O(n12635) );
  INV_GATE U12660 ( .I1(n12635), .O(n12150) );
  NAND_GATE U12661 ( .I1(n12634), .I2(n12150), .O(n12629) );
  NAND_GATE U12662 ( .I1(n12633), .I2(n12150), .O(n12628) );
  NAND3_GATE U12663 ( .I1(n12151), .I2(n12629), .I3(n12628), .O(n12421) );
  NAND_GATE U12664 ( .I1(B[6]), .I2(A[16]), .O(n12423) );
  OR_GATE U12665 ( .I1(n12152), .I2(n12157), .O(n12155) );
  OR_GATE U12666 ( .I1(n12153), .I2(n12156), .O(n12154) );
  AND_GATE U12667 ( .I1(n12155), .I2(n12154), .O(n12162) );
  NAND_GATE U12668 ( .I1(n12156), .I2(n961), .O(n12160) );
  NAND3_GATE U12669 ( .I1(n12160), .I2(n12159), .I3(n12158), .O(n12161) );
  NAND_GATE U12670 ( .I1(n12162), .I2(n12161), .O(n12418) );
  NAND_GATE U12671 ( .I1(n12423), .I2(n12418), .O(n12163) );
  NAND_GATE U12672 ( .I1(n12421), .I2(n12163), .O(n12164) );
  INV_GATE U12673 ( .I1(n12423), .O(n12420) );
  NAND_GATE U12674 ( .I1(n12420), .I2(n522), .O(n12416) );
  NAND_GATE U12675 ( .I1(n12164), .I2(n12416), .O(n12649) );
  NAND_GATE U12676 ( .I1(n12648), .I2(n12649), .O(n12166) );
  NAND_GATE U12677 ( .I1(B[6]), .I2(A[17]), .O(n12650) );
  INV_GATE U12678 ( .I1(n12650), .O(n12165) );
  NAND_GATE U12679 ( .I1(n12649), .I2(n12165), .O(n12645) );
  NAND_GATE U12680 ( .I1(n12648), .I2(n12165), .O(n12644) );
  NAND3_GATE U12681 ( .I1(n12166), .I2(n12645), .I3(n12644), .O(n12410) );
  NAND_GATE U12682 ( .I1(n12409), .I2(n12411), .O(n12167) );
  NAND_GATE U12683 ( .I1(n12410), .I2(n12167), .O(n12168) );
  NAND_GATE U12684 ( .I1(n12404), .I2(n12168), .O(n12398) );
  NAND_GATE U12685 ( .I1(n12182), .I2(n12398), .O(n12394) );
  INV_GATE U12686 ( .I1(n12169), .O(n12170) );
  NAND_GATE U12687 ( .I1(n12170), .I2(n12173), .O(n12181) );
  NAND_GATE U12688 ( .I1(n12171), .I2(n12175), .O(n12179) );
  NAND_GATE U12689 ( .I1(n12172), .I2(n627), .O(n12175) );
  NAND_GATE U12690 ( .I1(n605), .I2(n12173), .O(n12174) );
  NAND_GATE U12691 ( .I1(n12175), .I2(n12174), .O(n12176) );
  NAND_GATE U12692 ( .I1(n12177), .I2(n12176), .O(n12178) );
  NAND_GATE U12693 ( .I1(n12179), .I2(n12178), .O(n12180) );
  NAND_GATE U12694 ( .I1(n12181), .I2(n12180), .O(n12397) );
  NAND_GATE U12695 ( .I1(n12398), .I2(n12397), .O(n12183) );
  NAND_GATE U12696 ( .I1(n12182), .I2(n12397), .O(n12393) );
  NAND3_GATE U12697 ( .I1(n12394), .I2(n12183), .I3(n12393), .O(n12665) );
  NAND_GATE U12698 ( .I1(n12664), .I2(n12669), .O(n12184) );
  NAND_GATE U12699 ( .I1(n12665), .I2(n12184), .O(n12185) );
  NAND_GATE U12700 ( .I1(n12661), .I2(n12185), .O(n12387) );
  NAND_GATE U12701 ( .I1(n12199), .I2(n12387), .O(n12381) );
  NAND_GATE U12702 ( .I1(n12187), .I2(n12192), .O(n12196) );
  NAND_GATE U12703 ( .I1(n12189), .I2(n12188), .O(n12192) );
  NAND_GATE U12704 ( .I1(n1326), .I2(n12190), .O(n12191) );
  NAND_GATE U12705 ( .I1(n12192), .I2(n12191), .O(n12193) );
  NAND_GATE U12706 ( .I1(n12194), .I2(n12193), .O(n12195) );
  NAND_GATE U12707 ( .I1(n12196), .I2(n12195), .O(n12197) );
  NAND_GATE U12708 ( .I1(n12198), .I2(n12197), .O(n12385) );
  NAND_GATE U12709 ( .I1(n12387), .I2(n12385), .O(n12200) );
  NAND3_GATE U12710 ( .I1(n12381), .I2(n12200), .I3(n12380), .O(n12685) );
  NAND_GATE U12711 ( .I1(n12681), .I2(n12680), .O(n12201) );
  NAND_GATE U12712 ( .I1(n12685), .I2(n12201), .O(n12202) );
  NAND_GATE U12713 ( .I1(n12684), .I2(n12202), .O(n12374) );
  NAND_GATE U12714 ( .I1(n12368), .I2(n12374), .O(n12369) );
  INV_GATE U12715 ( .I1(n12203), .O(n12204) );
  NAND_GATE U12716 ( .I1(n12204), .I2(n12209), .O(n12215) );
  NAND_GATE U12717 ( .I1(n12208), .I2(n12207), .O(n12205) );
  NAND_GATE U12718 ( .I1(n12206), .I2(n12205), .O(n12213) );
  NAND_GATE U12719 ( .I1(n12213), .I2(n12212), .O(n12214) );
  NAND_GATE U12720 ( .I1(n12215), .I2(n12214), .O(n12373) );
  NAND_GATE U12721 ( .I1(n12374), .I2(n12373), .O(n12217) );
  NAND_GATE U12722 ( .I1(n12368), .I2(n12373), .O(n12216) );
  NAND_GATE U12723 ( .I1(n12366), .I2(n12365), .O(n12218) );
  NAND_GATE U12724 ( .I1(n12361), .I2(n12218), .O(n12219) );
  NAND_GATE U12725 ( .I1(n12358), .I2(n12219), .O(n12348) );
  NAND_GATE U12726 ( .I1(n12354), .I2(n12348), .O(n12221) );
  NAND_GATE U12727 ( .I1(B[6]), .I2(A[25]), .O(n12351) );
  INV_GATE U12728 ( .I1(n12351), .O(n12353) );
  NAND_GATE U12729 ( .I1(n12354), .I2(n12353), .O(n12220) );
  NAND_GATE U12730 ( .I1(n12348), .I2(n12353), .O(n12352) );
  NAND3_GATE U12731 ( .I1(n12221), .I2(n12220), .I3(n12352), .O(n12339) );
  NAND_GATE U12732 ( .I1(n12223), .I2(n12334), .O(n12328) );
  NAND3_GATE U12733 ( .I1(n12335), .I2(n12334), .I3(n12326), .O(n12224) );
  NAND3_GATE U12734 ( .I1(n12325), .I2(n12328), .I3(n12224), .O(n12319) );
  NAND_GATE U12735 ( .I1(n12321), .I2(n12319), .O(n12226) );
  NAND_GATE U12736 ( .I1(B[6]), .I2(A[28]), .O(n12316) );
  INV_GATE U12737 ( .I1(n12316), .O(n12320) );
  NAND_GATE U12738 ( .I1(n12320), .I2(n12319), .O(n12301) );
  NAND_GATE U12739 ( .I1(n12320), .I2(n12321), .O(n12225) );
  NAND3_GATE U12740 ( .I1(n12226), .I2(n12301), .I3(n12225), .O(n12308) );
  NAND_GATE U12741 ( .I1(n12302), .I2(n12308), .O(n12229) );
  NAND3_GATE U12742 ( .I1(n12227), .I2(n12308), .I3(n12307), .O(n12228) );
  NAND3_GATE U12743 ( .I1(n12230), .I2(n12229), .I3(n12228), .O(n12282) );
  NAND_GATE U12744 ( .I1(n12286), .I2(n12282), .O(n12287) );
  OR_GATE U12745 ( .I1(n12243), .I2(n12231), .O(n12234) );
  INV_GATE U12746 ( .I1(n12243), .O(n12237) );
  NAND_GATE U12747 ( .I1(n12232), .I2(n12237), .O(n12233) );
  NAND3_GATE U12748 ( .I1(n12235), .I2(n12234), .I3(n12233), .O(n12241) );
  NAND_GATE U12749 ( .I1(n589), .I2(n12243), .O(n12240) );
  NAND3_GATE U12750 ( .I1(n12238), .I2(n12237), .I3(n12236), .O(n12239) );
  NAND3_GATE U12751 ( .I1(n12241), .I2(n12240), .I3(n12239), .O(n12246) );
  INV_GATE U12752 ( .I1(n12242), .O(n12244) );
  NAND_GATE U12753 ( .I1(n12244), .I2(n12243), .O(n12245) );
  NAND_GATE U12754 ( .I1(n12246), .I2(n12245), .O(n12288) );
  NAND_GATE U12755 ( .I1(n12282), .I2(n12288), .O(n12248) );
  NAND_GATE U12756 ( .I1(n12286), .I2(n12288), .O(n12247) );
  NAND3_GATE U12757 ( .I1(n12287), .I2(n12248), .I3(n12247), .O(n12276) );
  NAND_GATE U12758 ( .I1(n12260), .I2(n12276), .O(n12261) );
  NAND3_GATE U12759 ( .I1(n12250), .I2(n12267), .I3(n623), .O(n12266) );
  NAND3_GATE U12760 ( .I1(n12268), .I2(n593), .I3(n12271), .O(n12251) );
  NAND_GATE U12761 ( .I1(n12268), .I2(n593), .O(n12249) );
  NAND3_GATE U12762 ( .I1(n12251), .I2(n12269), .I3(n12265), .O(n12252) );
  NAND_GATE U12763 ( .I1(n12266), .I2(n12252), .O(n12262) );
  NAND_GATE U12764 ( .I1(n12260), .I2(n12262), .O(n12254) );
  NAND_GATE U12765 ( .I1(n12276), .I2(n12262), .O(n12253) );
  NAND3_GATE U12766 ( .I1(n12261), .I2(n12254), .I3(n12253), .O(n15355) );
  NAND_GATE U12767 ( .I1(n12256), .I2(n12255), .O(n12257) );
  NAND_GATE U12768 ( .I1(n15355), .I2(n12257), .O(n12258) );
  NAND_GATE U12769 ( .I1(n12259), .I2(n12258), .O(\A1[36] ) );
  INV_GATE U12770 ( .I1(n12276), .O(n12272) );
  NAND3_GATE U12771 ( .I1(n12260), .I2(n12272), .I3(n12262), .O(n12264) );
  OR_GATE U12772 ( .I1(n12262), .I2(n12261), .O(n12263) );
  AND_GATE U12773 ( .I1(n12264), .I2(n12263), .O(n12281) );
  NAND_GATE U12774 ( .I1(n623), .I2(n12267), .O(n12269) );
  NAND_GATE U12775 ( .I1(n12269), .I2(n12249), .O(n12270) );
  NAND_GATE U12776 ( .I1(n12271), .I2(n12270), .O(n12273) );
  NAND3_GATE U12777 ( .I1(n12274), .I2(n12272), .I3(n12273), .O(n12278) );
  NAND_GATE U12778 ( .I1(n12274), .I2(n12273), .O(n12275) );
  NAND_GATE U12779 ( .I1(n12276), .I2(n12275), .O(n12277) );
  NAND3_GATE U12780 ( .I1(n12279), .I2(n12278), .I3(n12277), .O(n12280) );
  NAND_GATE U12781 ( .I1(n12282), .I2(n739), .O(n12284) );
  NAND_GATE U12782 ( .I1(n408), .I2(n12288), .O(n12283) );
  NAND3_GATE U12783 ( .I1(n12285), .I2(n12284), .I3(n12283), .O(n12291) );
  NAND3_GATE U12784 ( .I1(n408), .I2(n12288), .I3(n12286), .O(n12290) );
  OR_GATE U12785 ( .I1(n12288), .I2(n12287), .O(n12289) );
  NAND3_GATE U12786 ( .I1(n12291), .I2(n12290), .I3(n12289), .O(n12719) );
  NAND_GATE U12787 ( .I1(B[5]), .I2(A[31]), .O(n12717) );
  INV_GATE U12788 ( .I1(n12717), .O(n12721) );
  NAND_GATE U12789 ( .I1(B[5]), .I2(A[30]), .O(n12736) );
  INV_GATE U12790 ( .I1(n12736), .O(n12733) );
  NAND3_GATE U12791 ( .I1(n12294), .I2(n12293), .I3(n12292), .O(n12298) );
  NAND3_GATE U12792 ( .I1(n12298), .I2(n11859), .I3(n12297), .O(n12299) );
  NAND_GATE U12793 ( .I1(n12300), .I2(n12299), .O(n12309) );
  OR_GATE U12794 ( .I1(n12301), .I2(n12315), .O(n12305) );
  NAND3_GATE U12795 ( .I1(n12320), .I2(n12302), .I3(n12321), .O(n12304) );
  NAND3_GATE U12796 ( .I1(n12321), .I2(n12302), .I3(n12319), .O(n12303) );
  NAND3_GATE U12797 ( .I1(n12305), .I2(n12304), .I3(n12303), .O(n12306) );
  INV_GATE U12798 ( .I1(n12308), .O(n12310) );
  NAND3_GATE U12799 ( .I1(n12307), .I2(n12310), .I3(n918), .O(n12311) );
  NAND_GATE U12800 ( .I1(n12312), .I2(n12311), .O(n12730) );
  INV_GATE U12801 ( .I1(n12730), .O(n12735) );
  NAND_GATE U12802 ( .I1(n12310), .I2(n12309), .O(n12313) );
  NAND3_GATE U12803 ( .I1(n12314), .I2(n12313), .I3(n12315), .O(n12734) );
  NAND3_GATE U12804 ( .I1(n12733), .I2(n12735), .I3(n12734), .O(n12741) );
  NAND_GATE U12805 ( .I1(n12736), .I2(n12730), .O(n12711) );
  NAND4_GATE U12806 ( .I1(n12315), .I2(n12314), .I3(n12736), .I4(n12313), .O(
        n12710) );
  INV_GATE U12807 ( .I1(n12319), .O(n12322) );
  NAND_GATE U12808 ( .I1(n12321), .I2(n12322), .O(n12318) );
  NAND_GATE U12809 ( .I1(n677), .I2(n12319), .O(n12317) );
  NAND3_GATE U12810 ( .I1(n12318), .I2(n12317), .I3(n12316), .O(n12745) );
  NAND_GATE U12811 ( .I1(B[5]), .I2(A[29]), .O(n13163) );
  NAND3_GATE U12812 ( .I1(n12319), .I2(n677), .I3(n12320), .O(n12324) );
  NAND3_GATE U12813 ( .I1(n12322), .I2(n12321), .I3(n12320), .O(n12323) );
  AND_GATE U12814 ( .I1(n12324), .I2(n12323), .O(n12746) );
  NAND3_GATE U12815 ( .I1(n12745), .I2(n462), .I3(n12746), .O(n12709) );
  NAND_GATE U12816 ( .I1(B[5]), .I2(A[28]), .O(n13187) );
  INV_GATE U12817 ( .I1(n13187), .O(n13178) );
  NAND_GATE U12818 ( .I1(n12332), .I2(n12331), .O(n12326) );
  NAND_GATE U12819 ( .I1(n12330), .I2(n12329), .O(n12335) );
  NAND_GATE U12820 ( .I1(n12335), .I2(n12326), .O(n12333) );
  NAND_GATE U12821 ( .I1(n12334), .I2(n12333), .O(n12700) );
  NAND3_GATE U12822 ( .I1(n12326), .I2(n12335), .I3(n742), .O(n12699) );
  NAND3_GATE U12823 ( .I1(n12700), .I2(n12699), .I3(n12701), .O(n12752) );
  NAND3_GATE U12824 ( .I1(n742), .I2(n13187), .I3(n12336), .O(n12704) );
  NAND_GATE U12825 ( .I1(n13187), .I2(n1291), .O(n12703) );
  NAND_GATE U12826 ( .I1(B[5]), .I2(A[27]), .O(n13135) );
  INV_GATE U12827 ( .I1(n13135), .O(n12760) );
  NAND3_GATE U12828 ( .I1(n12338), .I2(n12341), .I3(n12342), .O(n12347) );
  NAND_GATE U12829 ( .I1(n12340), .I2(n12339), .O(n12346) );
  NAND_GATE U12830 ( .I1(n12342), .I2(n12341), .O(n12343) );
  NAND_GATE U12831 ( .I1(n12344), .I2(n12343), .O(n12345) );
  NAND3_GATE U12832 ( .I1(n12347), .I2(n12346), .I3(n12345), .O(n12757) );
  NAND_GATE U12833 ( .I1(n12756), .I2(n12757), .O(n13133) );
  NAND_GATE U12834 ( .I1(n12760), .I2(n13133), .O(n12698) );
  NAND_GATE U12835 ( .I1(B[5]), .I2(A[26]), .O(n12765) );
  INV_GATE U12836 ( .I1(n12765), .O(n12768) );
  NAND_GATE U12837 ( .I1(n12354), .I2(n525), .O(n12350) );
  NAND3_GATE U12838 ( .I1(n12351), .I2(n12350), .I3(n12349), .O(n12357) );
  OR_GATE U12839 ( .I1(n12352), .I2(n12354), .O(n12356) );
  NAND3_GATE U12840 ( .I1(n525), .I2(n12354), .I3(n12353), .O(n12355) );
  NAND3_GATE U12841 ( .I1(n12357), .I2(n12356), .I3(n12355), .O(n12766) );
  INV_GATE U12842 ( .I1(n12766), .O(n12764) );
  NAND_GATE U12843 ( .I1(B[5]), .I2(A[25]), .O(n12786) );
  INV_GATE U12844 ( .I1(n12786), .O(n12778) );
  NAND_GATE U12845 ( .I1(n12366), .I2(n1266), .O(n12359) );
  NAND_GATE U12846 ( .I1(n12360), .I2(n12359), .O(n12364) );
  NAND_GATE U12847 ( .I1(n12362), .I2(n12361), .O(n12363) );
  AND_GATE U12848 ( .I1(n12364), .I2(n12363), .O(n12787) );
  NAND3_GATE U12849 ( .I1(n12366), .I2(n1266), .I3(n12365), .O(n12785) );
  NAND_GATE U12850 ( .I1(n167), .I2(n12364), .O(n12367) );
  NAND_GATE U12851 ( .I1(n12782), .I2(n12367), .O(n12792) );
  NAND_GATE U12852 ( .I1(B[5]), .I2(A[24]), .O(n13117) );
  INV_GATE U12853 ( .I1(n13117), .O(n13116) );
  INV_GATE U12854 ( .I1(n12374), .O(n12372) );
  NAND3_GATE U12855 ( .I1(n12372), .I2(n12368), .I3(n12373), .O(n12371) );
  OR_GATE U12856 ( .I1(n12373), .I2(n12369), .O(n12370) );
  AND_GATE U12857 ( .I1(n12371), .I2(n12370), .O(n12379) );
  NAND_GATE U12858 ( .I1(n12372), .I2(n12373), .O(n12377) );
  NAND3_GATE U12859 ( .I1(n12377), .I2(n12376), .I3(n12375), .O(n12378) );
  NAND_GATE U12860 ( .I1(n12379), .I2(n12378), .O(n13119) );
  NAND_GATE U12861 ( .I1(n13116), .I2(n231), .O(n13123) );
  NAND_GATE U12862 ( .I1(B[5]), .I2(A[23]), .O(n13109) );
  INV_GATE U12863 ( .I1(n13109), .O(n13103) );
  OR_GATE U12864 ( .I1(n12380), .I2(n12387), .O(n12383) );
  OR_GATE U12865 ( .I1(n12385), .I2(n12381), .O(n12382) );
  AND_GATE U12866 ( .I1(n12383), .I2(n12382), .O(n12392) );
  INV_GATE U12867 ( .I1(n12387), .O(n12384) );
  NAND_GATE U12868 ( .I1(n12384), .I2(n12385), .O(n12390) );
  INV_GATE U12869 ( .I1(n12385), .O(n12386) );
  NAND_GATE U12870 ( .I1(n12387), .I2(n12386), .O(n12389) );
  NAND3_GATE U12871 ( .I1(n12390), .I2(n12389), .I3(n12388), .O(n12391) );
  NAND_GATE U12872 ( .I1(n12392), .I2(n12391), .O(n13091) );
  NAND_GATE U12873 ( .I1(B[5]), .I2(A[22]), .O(n13096) );
  INV_GATE U12874 ( .I1(n13096), .O(n13089) );
  NAND_GATE U12875 ( .I1(n328), .I2(n12391), .O(n13088) );
  NAND_GATE U12876 ( .I1(B[5]), .I2(A[21]), .O(n12802) );
  INV_GATE U12877 ( .I1(n12802), .O(n12674) );
  OR_GATE U12878 ( .I1(n12397), .I2(n12394), .O(n12395) );
  AND_GATE U12879 ( .I1(n12396), .I2(n12395), .O(n12403) );
  NAND_GATE U12880 ( .I1(n924), .I2(n12397), .O(n12401) );
  NAND3_GATE U12881 ( .I1(n12401), .I2(n12400), .I3(n12399), .O(n12402) );
  NAND_GATE U12882 ( .I1(n12403), .I2(n12402), .O(n12810) );
  INV_GATE U12883 ( .I1(n12810), .O(n12812) );
  NAND_GATE U12884 ( .I1(B[5]), .I2(A[20]), .O(n12814) );
  INV_GATE U12885 ( .I1(n12814), .O(n12809) );
  NAND_GATE U12886 ( .I1(n12812), .I2(n12809), .O(n12807) );
  INV_GATE U12887 ( .I1(n12404), .O(n12405) );
  NAND_GATE U12888 ( .I1(n12405), .I2(n12410), .O(n12415) );
  INV_GATE U12889 ( .I1(n12410), .O(n12408) );
  NAND_GATE U12890 ( .I1(n12409), .I2(n12408), .O(n12406) );
  NAND_GATE U12891 ( .I1(n12407), .I2(n12406), .O(n12413) );
  NAND_GATE U12892 ( .I1(n12413), .I2(n12412), .O(n12414) );
  NAND_GATE U12893 ( .I1(n12415), .I2(n12414), .O(n13076) );
  INV_GATE U12894 ( .I1(n12416), .O(n12417) );
  NAND_GATE U12895 ( .I1(n12421), .I2(n12417), .O(n12427) );
  INV_GATE U12896 ( .I1(n12421), .O(n12419) );
  NAND_GATE U12897 ( .I1(n12419), .I2(n12418), .O(n12422) );
  NAND_GATE U12898 ( .I1(n12420), .I2(n12422), .O(n12425) );
  NAND_GATE U12899 ( .I1(n12425), .I2(n12424), .O(n12426) );
  NAND_GATE U12900 ( .I1(n12427), .I2(n12426), .O(n13061) );
  INV_GATE U12901 ( .I1(n12428), .O(n12429) );
  NAND_GATE U12902 ( .I1(n12434), .I2(n12429), .O(n12442) );
  INV_GATE U12903 ( .I1(n12434), .O(n12431) );
  NAND_GATE U12904 ( .I1(n12431), .I2(n12430), .O(n12436) );
  NAND_GATE U12905 ( .I1(n12432), .I2(n12436), .O(n12440) );
  NAND_GATE U12906 ( .I1(n12434), .I2(n12433), .O(n12435) );
  NAND_GATE U12907 ( .I1(n12436), .I2(n12435), .O(n12437) );
  NAND_GATE U12908 ( .I1(n12438), .I2(n12437), .O(n12439) );
  NAND_GATE U12909 ( .I1(n12440), .I2(n12439), .O(n12441) );
  NAND_GATE U12910 ( .I1(n12442), .I2(n12441), .O(n13047) );
  INV_GATE U12911 ( .I1(n12443), .O(n12444) );
  NAND_GATE U12912 ( .I1(n12449), .I2(n12444), .O(n12457) );
  INV_GATE U12913 ( .I1(n12449), .O(n12446) );
  NAND_GATE U12914 ( .I1(n12446), .I2(n12445), .O(n12451) );
  NAND_GATE U12915 ( .I1(n12447), .I2(n12451), .O(n12455) );
  NAND_GATE U12916 ( .I1(n12449), .I2(n12448), .O(n12450) );
  NAND_GATE U12917 ( .I1(n12451), .I2(n12450), .O(n12452) );
  NAND_GATE U12918 ( .I1(n12453), .I2(n12452), .O(n12454) );
  NAND_GATE U12919 ( .I1(n12455), .I2(n12454), .O(n12456) );
  NAND_GATE U12920 ( .I1(n12457), .I2(n12456), .O(n13032) );
  OR_GATE U12921 ( .I1(n12458), .I2(n12460), .O(n12471) );
  NAND_GATE U12922 ( .I1(n12460), .I2(n12459), .O(n12465) );
  NAND_GATE U12923 ( .I1(n12461), .I2(n12465), .O(n12469) );
  NAND_GATE U12924 ( .I1(n12463), .I2(n12462), .O(n12464) );
  NAND_GATE U12925 ( .I1(n12465), .I2(n12464), .O(n12466) );
  NAND_GATE U12926 ( .I1(n12467), .I2(n12466), .O(n12468) );
  NAND_GATE U12927 ( .I1(n12469), .I2(n12468), .O(n12470) );
  NAND_GATE U12928 ( .I1(n12471), .I2(n12470), .O(n13017) );
  OR_GATE U12929 ( .I1(n12472), .I2(n12476), .O(n12475) );
  OR_GATE U12930 ( .I1(n12473), .I2(n12477), .O(n12474) );
  AND_GATE U12931 ( .I1(n12475), .I2(n12474), .O(n12482) );
  NAND_GATE U12932 ( .I1(n12476), .I2(n1015), .O(n12480) );
  NAND3_GATE U12933 ( .I1(n12480), .I2(n12479), .I3(n12478), .O(n12481) );
  NAND_GATE U12934 ( .I1(n12482), .I2(n12481), .O(n12875) );
  INV_GATE U12935 ( .I1(n12875), .O(n12878) );
  OR_GATE U12936 ( .I1(n12483), .I2(n12485), .O(n12496) );
  NAND_GATE U12937 ( .I1(n12485), .I2(n12484), .O(n12490) );
  NAND_GATE U12938 ( .I1(n12486), .I2(n12490), .O(n12494) );
  NAND_GATE U12939 ( .I1(n12488), .I2(n12487), .O(n12489) );
  NAND_GATE U12940 ( .I1(n12490), .I2(n12489), .O(n12491) );
  NAND_GATE U12941 ( .I1(n12492), .I2(n12491), .O(n12493) );
  NAND_GATE U12942 ( .I1(n12494), .I2(n12493), .O(n12495) );
  NAND_GATE U12943 ( .I1(n12496), .I2(n12495), .O(n12891) );
  OR_GATE U12944 ( .I1(n12497), .I2(n12501), .O(n12500) );
  OR_GATE U12945 ( .I1(n12498), .I2(n12502), .O(n12499) );
  AND_GATE U12946 ( .I1(n12500), .I2(n12499), .O(n12507) );
  NAND_GATE U12947 ( .I1(n12501), .I2(n1021), .O(n12505) );
  NAND3_GATE U12948 ( .I1(n12505), .I2(n12504), .I3(n12503), .O(n12506) );
  NAND_GATE U12949 ( .I1(n12507), .I2(n12506), .O(n12900) );
  INV_GATE U12950 ( .I1(n12900), .O(n12903) );
  OR_GATE U12951 ( .I1(n12508), .I2(n12510), .O(n12521) );
  NAND_GATE U12952 ( .I1(n12510), .I2(n12509), .O(n12515) );
  NAND_GATE U12953 ( .I1(n12511), .I2(n12515), .O(n12519) );
  NAND_GATE U12954 ( .I1(n12513), .I2(n12512), .O(n12514) );
  NAND_GATE U12955 ( .I1(n12515), .I2(n12514), .O(n12516) );
  NAND_GATE U12956 ( .I1(n12517), .I2(n12516), .O(n12518) );
  NAND_GATE U12957 ( .I1(n12519), .I2(n12518), .O(n12520) );
  NAND_GATE U12958 ( .I1(n12521), .I2(n12520), .O(n12916) );
  OR_GATE U12959 ( .I1(n12522), .I2(n12526), .O(n12525) );
  OR_GATE U12960 ( .I1(n12523), .I2(n12527), .O(n12524) );
  AND_GATE U12961 ( .I1(n12525), .I2(n12524), .O(n12532) );
  NAND_GATE U12962 ( .I1(n12526), .I2(n1115), .O(n12530) );
  NAND3_GATE U12963 ( .I1(n12530), .I2(n12529), .I3(n12528), .O(n12531) );
  NAND_GATE U12964 ( .I1(n12532), .I2(n12531), .O(n12925) );
  INV_GATE U12965 ( .I1(n12925), .O(n12928) );
  OR_GATE U12966 ( .I1(n12533), .I2(n12535), .O(n12546) );
  NAND_GATE U12967 ( .I1(n12535), .I2(n12534), .O(n12540) );
  NAND_GATE U12968 ( .I1(n12536), .I2(n12540), .O(n12544) );
  NAND_GATE U12969 ( .I1(n12538), .I2(n12537), .O(n12539) );
  NAND_GATE U12970 ( .I1(n12540), .I2(n12539), .O(n12541) );
  NAND_GATE U12971 ( .I1(n12542), .I2(n12541), .O(n12543) );
  NAND_GATE U12972 ( .I1(n12544), .I2(n12543), .O(n12545) );
  NAND_GATE U12973 ( .I1(n12546), .I2(n12545), .O(n12941) );
  OR_GATE U12974 ( .I1(n12547), .I2(n12551), .O(n12550) );
  OR_GATE U12975 ( .I1(n12548), .I2(n12552), .O(n12549) );
  AND_GATE U12976 ( .I1(n12550), .I2(n12549), .O(n12557) );
  NAND_GATE U12977 ( .I1(n12551), .I2(n1186), .O(n12555) );
  NAND3_GATE U12978 ( .I1(n12555), .I2(n12554), .I3(n12553), .O(n12556) );
  NAND_GATE U12979 ( .I1(n12557), .I2(n12556), .O(n12950) );
  INV_GATE U12980 ( .I1(n12950), .O(n12953) );
  INV_GATE U12981 ( .I1(n12558), .O(n12559) );
  NAND_GATE U12982 ( .I1(n12563), .I2(n12559), .O(n12571) );
  NAND_GATE U12983 ( .I1(n12561), .I2(n12565), .O(n12569) );
  NAND_GATE U12984 ( .I1(n12563), .I2(n12562), .O(n12564) );
  NAND_GATE U12985 ( .I1(n12565), .I2(n12564), .O(n12566) );
  NAND_GATE U12986 ( .I1(n12567), .I2(n12566), .O(n12568) );
  NAND_GATE U12987 ( .I1(n12569), .I2(n12568), .O(n12570) );
  NAND_GATE U12988 ( .I1(n12571), .I2(n12570), .O(n12966) );
  NAND_GATE U12989 ( .I1(n1370), .I2(A[0]), .O(n12572) );
  NAND_GATE U12990 ( .I1(n14781), .I2(n12572), .O(n12573) );
  NAND_GATE U12991 ( .I1(B[7]), .I2(n12573), .O(n12577) );
  NAND_GATE U12992 ( .I1(n1371), .I2(A[1]), .O(n12574) );
  NAND_GATE U12993 ( .I1(n14784), .I2(n12574), .O(n12575) );
  NAND_GATE U12994 ( .I1(B[6]), .I2(n12575), .O(n12576) );
  NAND_GATE U12995 ( .I1(n12577), .I2(n12576), .O(n12978) );
  NAND_GATE U12996 ( .I1(B[5]), .I2(A[2]), .O(n12982) );
  NAND3_GATE U12997 ( .I1(B[5]), .I2(B[6]), .I3(n1196), .O(n12975) );
  NAND_GATE U12998 ( .I1(n12982), .I2(n12975), .O(n12578) );
  NAND_GATE U12999 ( .I1(n12978), .I2(n12578), .O(n12579) );
  INV_GATE U13000 ( .I1(n12982), .O(n12976) );
  INV_GATE U13001 ( .I1(n12975), .O(n12977) );
  NAND_GATE U13002 ( .I1(n12976), .I2(n12977), .O(n12973) );
  NAND_GATE U13003 ( .I1(n12579), .I2(n12973), .O(n12967) );
  NAND_GATE U13004 ( .I1(n12966), .I2(n12967), .O(n12581) );
  NAND_GATE U13005 ( .I1(B[5]), .I2(A[3]), .O(n12968) );
  INV_GATE U13006 ( .I1(n12968), .O(n12580) );
  NAND_GATE U13007 ( .I1(n12966), .I2(n12580), .O(n12963) );
  NAND_GATE U13008 ( .I1(n12967), .I2(n12580), .O(n12962) );
  NAND3_GATE U13009 ( .I1(n12581), .I2(n12963), .I3(n12962), .O(n12952) );
  INV_GATE U13010 ( .I1(n12952), .O(n12949) );
  NAND_GATE U13011 ( .I1(B[5]), .I2(A[4]), .O(n12957) );
  NAND_GATE U13012 ( .I1(n12949), .I2(n12957), .O(n12582) );
  NAND_GATE U13013 ( .I1(n12953), .I2(n12582), .O(n12583) );
  INV_GATE U13014 ( .I1(n12957), .O(n12951) );
  NAND_GATE U13015 ( .I1(n12952), .I2(n12951), .O(n12948) );
  NAND_GATE U13016 ( .I1(n12583), .I2(n12948), .O(n12942) );
  NAND_GATE U13017 ( .I1(n12941), .I2(n12942), .O(n12585) );
  NAND_GATE U13018 ( .I1(B[5]), .I2(A[5]), .O(n12943) );
  INV_GATE U13019 ( .I1(n12943), .O(n12584) );
  NAND_GATE U13020 ( .I1(n12941), .I2(n12584), .O(n12938) );
  NAND_GATE U13021 ( .I1(n12942), .I2(n12584), .O(n12937) );
  NAND3_GATE U13022 ( .I1(n12585), .I2(n12938), .I3(n12937), .O(n12927) );
  INV_GATE U13023 ( .I1(n12927), .O(n12924) );
  NAND_GATE U13024 ( .I1(B[5]), .I2(A[6]), .O(n12932) );
  NAND_GATE U13025 ( .I1(n12924), .I2(n12932), .O(n12586) );
  NAND_GATE U13026 ( .I1(n12928), .I2(n12586), .O(n12587) );
  INV_GATE U13027 ( .I1(n12932), .O(n12926) );
  NAND_GATE U13028 ( .I1(n12927), .I2(n12926), .O(n12923) );
  NAND_GATE U13029 ( .I1(n12587), .I2(n12923), .O(n12917) );
  NAND_GATE U13030 ( .I1(n12916), .I2(n12917), .O(n12589) );
  NAND_GATE U13031 ( .I1(B[5]), .I2(A[7]), .O(n12918) );
  INV_GATE U13032 ( .I1(n12918), .O(n12588) );
  NAND_GATE U13033 ( .I1(n12916), .I2(n12588), .O(n12913) );
  NAND_GATE U13034 ( .I1(n12917), .I2(n12588), .O(n12912) );
  NAND3_GATE U13035 ( .I1(n12589), .I2(n12913), .I3(n12912), .O(n12902) );
  INV_GATE U13036 ( .I1(n12902), .O(n12899) );
  NAND_GATE U13037 ( .I1(B[5]), .I2(A[8]), .O(n12907) );
  NAND_GATE U13038 ( .I1(n12899), .I2(n12907), .O(n12590) );
  NAND_GATE U13039 ( .I1(n12903), .I2(n12590), .O(n12591) );
  INV_GATE U13040 ( .I1(n12907), .O(n12901) );
  NAND_GATE U13041 ( .I1(n12902), .I2(n12901), .O(n12898) );
  NAND_GATE U13042 ( .I1(n12591), .I2(n12898), .O(n12892) );
  NAND_GATE U13043 ( .I1(n12891), .I2(n12892), .O(n12593) );
  NAND_GATE U13044 ( .I1(B[5]), .I2(A[9]), .O(n12893) );
  INV_GATE U13045 ( .I1(n12893), .O(n12592) );
  NAND_GATE U13046 ( .I1(n12891), .I2(n12592), .O(n12888) );
  NAND_GATE U13047 ( .I1(n12892), .I2(n12592), .O(n12887) );
  NAND3_GATE U13048 ( .I1(n12593), .I2(n12888), .I3(n12887), .O(n12877) );
  INV_GATE U13049 ( .I1(n12877), .O(n12874) );
  NAND_GATE U13050 ( .I1(B[5]), .I2(A[10]), .O(n12882) );
  NAND_GATE U13051 ( .I1(n12874), .I2(n12882), .O(n12594) );
  NAND_GATE U13052 ( .I1(n12878), .I2(n12594), .O(n12595) );
  INV_GATE U13053 ( .I1(n12882), .O(n12876) );
  NAND_GATE U13054 ( .I1(n12877), .I2(n12876), .O(n12873) );
  NAND_GATE U13055 ( .I1(n12595), .I2(n12873), .O(n13018) );
  NAND_GATE U13056 ( .I1(n13017), .I2(n13018), .O(n12597) );
  NAND_GATE U13057 ( .I1(B[5]), .I2(A[11]), .O(n13019) );
  INV_GATE U13058 ( .I1(n13019), .O(n12596) );
  NAND_GATE U13059 ( .I1(n13018), .I2(n12596), .O(n13014) );
  NAND_GATE U13060 ( .I1(n13017), .I2(n12596), .O(n13013) );
  NAND3_GATE U13061 ( .I1(n12597), .I2(n13014), .I3(n13013), .O(n12864) );
  NAND_GATE U13062 ( .I1(B[5]), .I2(A[12]), .O(n12868) );
  OR_GATE U13063 ( .I1(n12598), .I2(n12603), .O(n12601) );
  OR_GATE U13064 ( .I1(n12599), .I2(n12602), .O(n12600) );
  AND_GATE U13065 ( .I1(n12601), .I2(n12600), .O(n12608) );
  NAND_GATE U13066 ( .I1(n12602), .I2(n1003), .O(n12606) );
  NAND3_GATE U13067 ( .I1(n12606), .I2(n12605), .I3(n12604), .O(n12607) );
  NAND_GATE U13068 ( .I1(n12608), .I2(n12607), .O(n12860) );
  NAND_GATE U13069 ( .I1(n12868), .I2(n12860), .O(n12609) );
  NAND_GATE U13070 ( .I1(n12864), .I2(n12609), .O(n12610) );
  INV_GATE U13071 ( .I1(n12868), .O(n12862) );
  INV_GATE U13072 ( .I1(n12860), .O(n12863) );
  NAND_GATE U13073 ( .I1(n12862), .I2(n12863), .O(n12858) );
  NAND_GATE U13074 ( .I1(n12610), .I2(n12858), .O(n13033) );
  NAND_GATE U13075 ( .I1(n13032), .I2(n13033), .O(n12612) );
  NAND_GATE U13076 ( .I1(B[5]), .I2(A[13]), .O(n13034) );
  INV_GATE U13077 ( .I1(n13034), .O(n12611) );
  NAND_GATE U13078 ( .I1(n13033), .I2(n12611), .O(n13029) );
  NAND_GATE U13079 ( .I1(n13032), .I2(n12611), .O(n13028) );
  NAND3_GATE U13080 ( .I1(n12612), .I2(n13029), .I3(n13028), .O(n12849) );
  NAND_GATE U13081 ( .I1(B[5]), .I2(A[14]), .O(n12853) );
  OR_GATE U13082 ( .I1(n12614), .I2(n12617), .O(n12615) );
  AND_GATE U13083 ( .I1(n12616), .I2(n12615), .O(n12623) );
  NAND_GATE U13084 ( .I1(n12617), .I2(n964), .O(n12621) );
  NAND3_GATE U13085 ( .I1(n12621), .I2(n12620), .I3(n12619), .O(n12622) );
  NAND_GATE U13086 ( .I1(n12623), .I2(n12622), .O(n12845) );
  NAND_GATE U13087 ( .I1(n12853), .I2(n12845), .O(n12624) );
  NAND_GATE U13088 ( .I1(n12849), .I2(n12624), .O(n12625) );
  INV_GATE U13089 ( .I1(n12853), .O(n12847) );
  INV_GATE U13090 ( .I1(n12845), .O(n12848) );
  NAND_GATE U13091 ( .I1(n12847), .I2(n12848), .O(n12843) );
  NAND_GATE U13092 ( .I1(n12625), .I2(n12843), .O(n13048) );
  NAND_GATE U13093 ( .I1(n13047), .I2(n13048), .O(n12627) );
  NAND_GATE U13094 ( .I1(B[5]), .I2(A[15]), .O(n13049) );
  INV_GATE U13095 ( .I1(n13049), .O(n12626) );
  NAND_GATE U13096 ( .I1(n13048), .I2(n12626), .O(n13044) );
  NAND_GATE U13097 ( .I1(n13047), .I2(n12626), .O(n13043) );
  NAND3_GATE U13098 ( .I1(n12627), .I2(n13044), .I3(n13043), .O(n12834) );
  NAND_GATE U13099 ( .I1(B[5]), .I2(A[16]), .O(n12838) );
  OR_GATE U13100 ( .I1(n12629), .I2(n12633), .O(n12630) );
  AND_GATE U13101 ( .I1(n12631), .I2(n12630), .O(n12639) );
  INV_GATE U13102 ( .I1(n12634), .O(n12632) );
  NAND_GATE U13103 ( .I1(n12633), .I2(n12632), .O(n12637) );
  NAND_GATE U13104 ( .I1(n1285), .I2(n12634), .O(n12636) );
  NAND3_GATE U13105 ( .I1(n12637), .I2(n12636), .I3(n12635), .O(n12638) );
  NAND_GATE U13106 ( .I1(n12639), .I2(n12638), .O(n12831) );
  NAND_GATE U13107 ( .I1(n12838), .I2(n12831), .O(n12640) );
  NAND_GATE U13108 ( .I1(n12834), .I2(n12640), .O(n12641) );
  INV_GATE U13109 ( .I1(n12838), .O(n12832) );
  INV_GATE U13110 ( .I1(n12831), .O(n12833) );
  NAND_GATE U13111 ( .I1(n12832), .I2(n12833), .O(n12830) );
  NAND_GATE U13112 ( .I1(n12641), .I2(n12830), .O(n13062) );
  NAND_GATE U13113 ( .I1(n13061), .I2(n13062), .O(n12643) );
  NAND_GATE U13114 ( .I1(B[5]), .I2(A[17]), .O(n13063) );
  INV_GATE U13115 ( .I1(n13063), .O(n12642) );
  NAND_GATE U13116 ( .I1(n13062), .I2(n12642), .O(n13058) );
  NAND3_GATE U13117 ( .I1(n12643), .I2(n13058), .I3(n13057), .O(n12823) );
  NAND_GATE U13118 ( .I1(B[5]), .I2(A[18]), .O(n12827) );
  OR_GATE U13119 ( .I1(n12644), .I2(n12649), .O(n12647) );
  OR_GATE U13120 ( .I1(n12645), .I2(n12648), .O(n12646) );
  AND_GATE U13121 ( .I1(n12647), .I2(n12646), .O(n12654) );
  NAND_GATE U13122 ( .I1(n12648), .I2(n929), .O(n12652) );
  NAND3_GATE U13123 ( .I1(n12652), .I2(n12651), .I3(n12650), .O(n12653) );
  NAND_GATE U13124 ( .I1(n12654), .I2(n12653), .O(n12820) );
  NAND_GATE U13125 ( .I1(n12827), .I2(n12820), .O(n12655) );
  NAND_GATE U13126 ( .I1(n12823), .I2(n12655), .O(n12656) );
  INV_GATE U13127 ( .I1(n12827), .O(n12822) );
  NAND_GATE U13128 ( .I1(n12822), .I2(n550), .O(n12819) );
  NAND_GATE U13129 ( .I1(n12656), .I2(n12819), .O(n13077) );
  NAND_GATE U13130 ( .I1(n13076), .I2(n13077), .O(n12658) );
  NAND_GATE U13131 ( .I1(B[5]), .I2(A[19]), .O(n13078) );
  INV_GATE U13132 ( .I1(n13078), .O(n12657) );
  NAND_GATE U13133 ( .I1(n13077), .I2(n12657), .O(n13073) );
  NAND_GATE U13134 ( .I1(n13076), .I2(n12657), .O(n13072) );
  NAND3_GATE U13135 ( .I1(n12658), .I2(n13073), .I3(n13072), .O(n12811) );
  NAND_GATE U13136 ( .I1(n12810), .I2(n12814), .O(n12659) );
  NAND_GATE U13137 ( .I1(n12811), .I2(n12659), .O(n12660) );
  NAND_GATE U13138 ( .I1(n12807), .I2(n12660), .O(n12801) );
  NAND_GATE U13139 ( .I1(n12674), .I2(n12801), .O(n12797) );
  INV_GATE U13140 ( .I1(n12661), .O(n12662) );
  NAND_GATE U13141 ( .I1(n12662), .I2(n12665), .O(n12673) );
  NAND_GATE U13142 ( .I1(n12663), .I2(n12667), .O(n12671) );
  NAND_GATE U13143 ( .I1(n12664), .I2(n507), .O(n12667) );
  NAND_GATE U13144 ( .I1(n625), .I2(n12665), .O(n12666) );
  NAND_GATE U13145 ( .I1(n12667), .I2(n12666), .O(n12668) );
  NAND_GATE U13146 ( .I1(n12669), .I2(n12668), .O(n12670) );
  NAND_GATE U13147 ( .I1(n12671), .I2(n12670), .O(n12672) );
  NAND_GATE U13148 ( .I1(n12673), .I2(n12672), .O(n12800) );
  NAND_GATE U13149 ( .I1(n12801), .I2(n12800), .O(n12675) );
  NAND3_GATE U13150 ( .I1(n12797), .I2(n12675), .I3(n12796), .O(n13092) );
  NAND_GATE U13151 ( .I1(n13091), .I2(n13096), .O(n12676) );
  NAND_GATE U13152 ( .I1(n13092), .I2(n12676), .O(n12689) );
  INV_GATE U13153 ( .I1(n12685), .O(n12679) );
  NAND_GATE U13154 ( .I1(n12680), .I2(n12679), .O(n12677) );
  NAND_GATE U13155 ( .I1(n339), .I2(n12677), .O(n12683) );
  NAND_GATE U13156 ( .I1(n12683), .I2(n12682), .O(n12688) );
  INV_GATE U13157 ( .I1(n12684), .O(n12686) );
  NAND_GATE U13158 ( .I1(n12686), .I2(n12685), .O(n12687) );
  NAND_GATE U13159 ( .I1(n12688), .I2(n12687), .O(n13106) );
  NAND3_GATE U13160 ( .I1(n12689), .I2(n13088), .I3(n13109), .O(n12690) );
  NAND_GATE U13161 ( .I1(n13106), .I2(n12690), .O(n12691) );
  NAND_GATE U13162 ( .I1(n13102), .I2(n12691), .O(n13124) );
  NAND_GATE U13163 ( .I1(n13117), .I2(n13119), .O(n12692) );
  NAND_GATE U13164 ( .I1(n13124), .I2(n12692), .O(n12784) );
  NAND_GATE U13165 ( .I1(n13123), .I2(n12784), .O(n12777) );
  NAND_GATE U13166 ( .I1(n12792), .I2(n12777), .O(n12693) );
  NAND3_GATE U13167 ( .I1(n12694), .I2(n12693), .I3(n12779), .O(n12773) );
  NAND_GATE U13168 ( .I1(n12765), .I2(n12766), .O(n12695) );
  NAND_GATE U13169 ( .I1(n12773), .I2(n12695), .O(n12696) );
  NAND_GATE U13170 ( .I1(n12772), .I2(n12696), .O(n12758) );
  NAND_GATE U13171 ( .I1(n12758), .I2(n13133), .O(n12697) );
  NAND_GATE U13172 ( .I1(n12760), .I2(n12758), .O(n12759) );
  NAND3_GATE U13173 ( .I1(n12698), .I2(n12697), .I3(n12759), .O(n13179) );
  NAND4_GATE U13174 ( .I1(n12701), .I2(n13187), .I3(n12700), .I4(n12699), .O(
        n12702) );
  NAND4_GATE U13175 ( .I1(n12704), .I2(n12703), .I3(n13179), .I4(n12702), .O(
        n12705) );
  NAND_GATE U13176 ( .I1(n12706), .I2(n12705), .O(n13160) );
  NAND_GATE U13177 ( .I1(n462), .I2(n13160), .O(n12708) );
  NAND3_GATE U13178 ( .I1(n13160), .I2(n12745), .I3(n12746), .O(n12707) );
  NAND3_GATE U13179 ( .I1(n12709), .I2(n12708), .I3(n12707), .O(n12742) );
  NAND3_GATE U13180 ( .I1(n12711), .I2(n12710), .I3(n12742), .O(n12712) );
  NAND_GATE U13181 ( .I1(n12719), .I2(n12717), .O(n12713) );
  NAND_GATE U13182 ( .I1(n12726), .I2(n12713), .O(n12714) );
  NAND_GATE U13183 ( .I1(n12725), .I2(n12714), .O(n15356) );
  NAND_GATE U13184 ( .I1(n488), .I2(n15356), .O(n12716) );
  AND_GATE U13185 ( .I1(n12716), .I2(n12715), .O(\A1[35] ) );
  NAND3_GATE U13186 ( .I1(n12717), .I2(n157), .I3(n12719), .O(n12724) );
  NAND_GATE U13187 ( .I1(n12718), .I2(n12726), .O(n12723) );
  NAND_GATE U13188 ( .I1(n12719), .I2(n157), .O(n12720) );
  NAND_GATE U13189 ( .I1(n12721), .I2(n12720), .O(n12722) );
  NAND3_GATE U13190 ( .I1(n12724), .I2(n12723), .I3(n12722), .O(n12729) );
  INV_GATE U13191 ( .I1(n12725), .O(n12727) );
  NAND_GATE U13192 ( .I1(n12727), .I2(n12726), .O(n12728) );
  NAND_GATE U13193 ( .I1(n12729), .I2(n12728), .O(n15358) );
  OR_GATE U13194 ( .I1(n12742), .I2(n12734), .O(n12732) );
  INV_GATE U13195 ( .I1(n12742), .O(n12737) );
  NAND_GATE U13196 ( .I1(n12730), .I2(n12737), .O(n12731) );
  NAND3_GATE U13197 ( .I1(n12733), .I2(n12732), .I3(n12731), .O(n12740) );
  NAND_GATE U13198 ( .I1(n12742), .I2(n1213), .O(n12739) );
  NAND3_GATE U13199 ( .I1(n12740), .I2(n12739), .I3(n12738), .O(n12744) );
  NAND_GATE U13200 ( .I1(n12744), .I2(n12743), .O(n13580) );
  NAND_GATE U13201 ( .I1(B[4]), .I2(A[31]), .O(n13581) );
  INV_GATE U13202 ( .I1(n13581), .O(n13577) );
  NAND_GATE U13203 ( .I1(n13580), .I2(n13577), .O(n13148) );
  NAND_GATE U13204 ( .I1(B[4]), .I2(A[30]), .O(n13171) );
  INV_GATE U13205 ( .I1(n13171), .O(n13152) );
  NAND_GATE U13206 ( .I1(n12746), .I2(n12745), .O(n13161) );
  NAND3_GATE U13207 ( .I1(n462), .I2(n13160), .I3(n13159), .O(n13158) );
  NAND3_GATE U13208 ( .I1(n13161), .I2(n624), .I3(n13163), .O(n12748) );
  NAND_GATE U13209 ( .I1(n13160), .I2(n13159), .O(n12747) );
  NAND_GATE U13210 ( .I1(n462), .I2(n13162), .O(n13157) );
  NAND3_GATE U13211 ( .I1(n12748), .I2(n12747), .I3(n13157), .O(n12749) );
  NAND_GATE U13212 ( .I1(n13158), .I2(n12749), .O(n13154) );
  NAND_GATE U13213 ( .I1(n13152), .I2(n13154), .O(n13145) );
  NAND_GATE U13214 ( .I1(n745), .I2(n400), .O(n12750) );
  NAND_GATE U13215 ( .I1(n13181), .I2(n12750), .O(n13186) );
  NAND3_GATE U13216 ( .I1(n13179), .I2(n1354), .I3(n13178), .O(n13185) );
  NAND_GATE U13217 ( .I1(n13178), .I2(n13179), .O(n12754) );
  NAND3_GATE U13218 ( .I1(n12752), .I2(n12751), .I3(n13178), .O(n12753) );
  NAND_GATE U13219 ( .I1(n12754), .I2(n12753), .O(n12755) );
  NAND_GATE U13220 ( .I1(n13185), .I2(n12755), .O(n13140) );
  NAND_GATE U13221 ( .I1(B[4]), .I2(A[29]), .O(n13569) );
  INV_GATE U13222 ( .I1(n13569), .O(n13175) );
  NAND_GATE U13223 ( .I1(n13188), .I2(n978), .O(n13143) );
  NAND3_GATE U13224 ( .I1(n12757), .I2(n12756), .I3(n12758), .O(n13136) );
  NAND_GATE U13225 ( .I1(n611), .I2(n13133), .O(n13134) );
  NAND_GATE U13226 ( .I1(B[4]), .I2(A[28]), .O(n13607) );
  NAND4_GATE U13227 ( .I1(n13136), .I2(n13134), .I3(n13135), .I4(n13607), .O(
        n12763) );
  NAND_GATE U13228 ( .I1(n13133), .I2(n920), .O(n12761) );
  AND_GATE U13229 ( .I1(n12763), .I2(n12762), .O(n13174) );
  NAND_GATE U13230 ( .I1(B[4]), .I2(A[27]), .O(n13561) );
  INV_GATE U13231 ( .I1(n13561), .O(n13196) );
  NAND_GATE U13232 ( .I1(n12764), .I2(n12773), .O(n12771) );
  NAND3_GATE U13233 ( .I1(n12765), .I2(n12766), .I3(n528), .O(n12770) );
  NAND_GATE U13234 ( .I1(n12766), .I2(n528), .O(n12767) );
  NAND_GATE U13235 ( .I1(n12768), .I2(n12767), .O(n12769) );
  NAND3_GATE U13236 ( .I1(n12771), .I2(n12770), .I3(n12769), .O(n12776) );
  INV_GATE U13237 ( .I1(n12772), .O(n12774) );
  NAND_GATE U13238 ( .I1(n12774), .I2(n12773), .O(n12775) );
  NAND_GATE U13239 ( .I1(n12776), .I2(n12775), .O(n13197) );
  NAND_GATE U13240 ( .I1(n13196), .I2(n13197), .O(n13132) );
  NAND_GATE U13241 ( .I1(B[4]), .I2(A[26]), .O(n13203) );
  INV_GATE U13242 ( .I1(n13203), .O(n13202) );
  NAND3_GATE U13243 ( .I1(n12778), .I2(n12791), .I3(n12792), .O(n12781) );
  OR_GATE U13244 ( .I1(n12779), .I2(n12792), .O(n12780) );
  INV_GATE U13245 ( .I1(n12782), .O(n12783) );
  NAND_GATE U13246 ( .I1(n12786), .I2(n12783), .O(n12790) );
  NAND3_GATE U13247 ( .I1(n13123), .I2(n12786), .I3(n12784), .O(n12789) );
  NAND3_GATE U13248 ( .I1(n12787), .I2(n12786), .I3(n12785), .O(n12788) );
  NAND3_GATE U13249 ( .I1(n12790), .I2(n12789), .I3(n12788), .O(n12794) );
  NAND_GATE U13250 ( .I1(n12792), .I2(n12791), .O(n12793) );
  NAND_GATE U13251 ( .I1(n12794), .I2(n12793), .O(n12795) );
  NAND_GATE U13252 ( .I1(n13202), .I2(n240), .O(n13209) );
  NAND_GATE U13253 ( .I1(B[4]), .I2(A[23]), .O(n13240) );
  INV_GATE U13254 ( .I1(n13240), .O(n13100) );
  OR_GATE U13255 ( .I1(n12796), .I2(n12801), .O(n12799) );
  OR_GATE U13256 ( .I1(n12800), .I2(n12797), .O(n12798) );
  AND_GATE U13257 ( .I1(n12799), .I2(n12798), .O(n12806) );
  NAND_GATE U13258 ( .I1(n116), .I2(n12800), .O(n12804) );
  NAND3_GATE U13259 ( .I1(n12804), .I2(n12803), .I3(n12802), .O(n12805) );
  NAND_GATE U13260 ( .I1(n12806), .I2(n12805), .O(n13248) );
  NAND_GATE U13261 ( .I1(B[4]), .I2(A[22]), .O(n13250) );
  INV_GATE U13262 ( .I1(n13250), .O(n13247) );
  INV_GATE U13263 ( .I1(n12807), .O(n12808) );
  NAND_GATE U13264 ( .I1(n12808), .I2(n12811), .O(n12818) );
  NAND_GATE U13265 ( .I1(n12809), .I2(n12813), .O(n12816) );
  NAND_GATE U13266 ( .I1(n12810), .I2(n124), .O(n12813) );
  NAND_GATE U13267 ( .I1(n12816), .I2(n12815), .O(n12817) );
  NAND_GATE U13268 ( .I1(n12818), .I2(n12817), .O(n13539) );
  INV_GATE U13269 ( .I1(n12823), .O(n12821) );
  NAND_GATE U13270 ( .I1(n12821), .I2(n12820), .O(n12825) );
  NAND_GATE U13271 ( .I1(n12822), .I2(n12825), .O(n12828) );
  NAND_GATE U13272 ( .I1(n12823), .I2(n550), .O(n12824) );
  NAND_GATE U13273 ( .I1(n12825), .I2(n12824), .O(n12826) );
  NAND_GATE U13274 ( .I1(n12832), .I2(n12836), .O(n12840) );
  NAND_GATE U13275 ( .I1(n12834), .I2(n12833), .O(n12835) );
  NAND_GATE U13276 ( .I1(n12836), .I2(n12835), .O(n12837) );
  NAND_GATE U13277 ( .I1(n12838), .I2(n12837), .O(n12839) );
  NAND_GATE U13278 ( .I1(n12840), .I2(n12839), .O(n12841) );
  INV_GATE U13279 ( .I1(n12843), .O(n12844) );
  NAND_GATE U13280 ( .I1(n12849), .I2(n12844), .O(n12857) );
  INV_GATE U13281 ( .I1(n12849), .O(n12846) );
  NAND_GATE U13282 ( .I1(n12846), .I2(n12845), .O(n12851) );
  NAND_GATE U13283 ( .I1(n12847), .I2(n12851), .O(n12855) );
  NAND_GATE U13284 ( .I1(n12849), .I2(n12848), .O(n12850) );
  NAND_GATE U13285 ( .I1(n12851), .I2(n12850), .O(n12852) );
  NAND_GATE U13286 ( .I1(n12853), .I2(n12852), .O(n12854) );
  NAND_GATE U13287 ( .I1(n12855), .I2(n12854), .O(n12856) );
  NAND_GATE U13288 ( .I1(n12857), .I2(n12856), .O(n13494) );
  INV_GATE U13289 ( .I1(n12858), .O(n12859) );
  NAND_GATE U13290 ( .I1(n12864), .I2(n12859), .O(n12872) );
  INV_GATE U13291 ( .I1(n12864), .O(n12861) );
  NAND_GATE U13292 ( .I1(n12861), .I2(n12860), .O(n12866) );
  NAND_GATE U13293 ( .I1(n12862), .I2(n12866), .O(n12870) );
  NAND_GATE U13294 ( .I1(n12864), .I2(n12863), .O(n12865) );
  NAND_GATE U13295 ( .I1(n12866), .I2(n12865), .O(n12867) );
  NAND_GATE U13296 ( .I1(n12868), .I2(n12867), .O(n12869) );
  NAND_GATE U13297 ( .I1(n12870), .I2(n12869), .O(n12871) );
  NAND_GATE U13298 ( .I1(n12872), .I2(n12871), .O(n13480) );
  OR_GATE U13299 ( .I1(n12873), .I2(n12875), .O(n12886) );
  NAND_GATE U13300 ( .I1(n12875), .I2(n12874), .O(n12880) );
  NAND_GATE U13301 ( .I1(n12876), .I2(n12880), .O(n12884) );
  NAND_GATE U13302 ( .I1(n12878), .I2(n12877), .O(n12879) );
  NAND_GATE U13303 ( .I1(n12880), .I2(n12879), .O(n12881) );
  NAND_GATE U13304 ( .I1(n12882), .I2(n12881), .O(n12883) );
  NAND_GATE U13305 ( .I1(n12884), .I2(n12883), .O(n12885) );
  NAND_GATE U13306 ( .I1(n12886), .I2(n12885), .O(n13465) );
  OR_GATE U13307 ( .I1(n12887), .I2(n12891), .O(n12890) );
  OR_GATE U13308 ( .I1(n12888), .I2(n12892), .O(n12889) );
  AND_GATE U13309 ( .I1(n12890), .I2(n12889), .O(n12897) );
  NAND_GATE U13310 ( .I1(n12891), .I2(n1019), .O(n12895) );
  NAND3_GATE U13311 ( .I1(n12895), .I2(n12894), .I3(n12893), .O(n12896) );
  NAND_GATE U13312 ( .I1(n12897), .I2(n12896), .O(n13323) );
  INV_GATE U13313 ( .I1(n13323), .O(n13326) );
  OR_GATE U13314 ( .I1(n12898), .I2(n12900), .O(n12911) );
  NAND_GATE U13315 ( .I1(n12900), .I2(n12899), .O(n12905) );
  NAND_GATE U13316 ( .I1(n12901), .I2(n12905), .O(n12909) );
  NAND_GATE U13317 ( .I1(n12903), .I2(n12902), .O(n12904) );
  NAND_GATE U13318 ( .I1(n12905), .I2(n12904), .O(n12906) );
  NAND_GATE U13319 ( .I1(n12907), .I2(n12906), .O(n12908) );
  NAND_GATE U13320 ( .I1(n12909), .I2(n12908), .O(n12910) );
  NAND_GATE U13321 ( .I1(n12911), .I2(n12910), .O(n13339) );
  OR_GATE U13322 ( .I1(n12912), .I2(n12916), .O(n12915) );
  OR_GATE U13323 ( .I1(n12913), .I2(n12917), .O(n12914) );
  AND_GATE U13324 ( .I1(n12915), .I2(n12914), .O(n12922) );
  NAND_GATE U13325 ( .I1(n12916), .I2(n1023), .O(n12920) );
  NAND3_GATE U13326 ( .I1(n12920), .I2(n12919), .I3(n12918), .O(n12921) );
  NAND_GATE U13327 ( .I1(n12922), .I2(n12921), .O(n13348) );
  INV_GATE U13328 ( .I1(n13348), .O(n13351) );
  OR_GATE U13329 ( .I1(n12923), .I2(n12925), .O(n12936) );
  NAND_GATE U13330 ( .I1(n12925), .I2(n12924), .O(n12930) );
  NAND_GATE U13331 ( .I1(n12926), .I2(n12930), .O(n12934) );
  NAND_GATE U13332 ( .I1(n12928), .I2(n12927), .O(n12929) );
  NAND_GATE U13333 ( .I1(n12930), .I2(n12929), .O(n12931) );
  NAND_GATE U13334 ( .I1(n12932), .I2(n12931), .O(n12933) );
  NAND_GATE U13335 ( .I1(n12934), .I2(n12933), .O(n12935) );
  NAND_GATE U13336 ( .I1(n12936), .I2(n12935), .O(n13364) );
  OR_GATE U13337 ( .I1(n12937), .I2(n12941), .O(n12940) );
  OR_GATE U13338 ( .I1(n12938), .I2(n12942), .O(n12939) );
  AND_GATE U13339 ( .I1(n12940), .I2(n12939), .O(n12947) );
  NAND_GATE U13340 ( .I1(n12941), .I2(n1116), .O(n12945) );
  NAND3_GATE U13341 ( .I1(n12945), .I2(n12944), .I3(n12943), .O(n12946) );
  NAND_GATE U13342 ( .I1(n12947), .I2(n12946), .O(n13373) );
  INV_GATE U13343 ( .I1(n13373), .O(n13376) );
  OR_GATE U13344 ( .I1(n12948), .I2(n12950), .O(n12961) );
  NAND_GATE U13345 ( .I1(n12950), .I2(n12949), .O(n12955) );
  NAND_GATE U13346 ( .I1(n12951), .I2(n12955), .O(n12959) );
  NAND_GATE U13347 ( .I1(n12953), .I2(n12952), .O(n12954) );
  NAND_GATE U13348 ( .I1(n12955), .I2(n12954), .O(n12956) );
  NAND_GATE U13349 ( .I1(n12957), .I2(n12956), .O(n12958) );
  NAND_GATE U13350 ( .I1(n12959), .I2(n12958), .O(n12960) );
  NAND_GATE U13351 ( .I1(n12961), .I2(n12960), .O(n13389) );
  OR_GATE U13352 ( .I1(n12962), .I2(n12966), .O(n12965) );
  OR_GATE U13353 ( .I1(n12963), .I2(n12967), .O(n12964) );
  AND_GATE U13354 ( .I1(n12965), .I2(n12964), .O(n12972) );
  NAND_GATE U13355 ( .I1(n12966), .I2(n1187), .O(n12970) );
  NAND3_GATE U13356 ( .I1(n12970), .I2(n12969), .I3(n12968), .O(n12971) );
  NAND_GATE U13357 ( .I1(n12972), .I2(n12971), .O(n13398) );
  INV_GATE U13358 ( .I1(n13398), .O(n13401) );
  INV_GATE U13359 ( .I1(n12973), .O(n12974) );
  NAND_GATE U13360 ( .I1(n12978), .I2(n12974), .O(n12986) );
  NAND_GATE U13361 ( .I1(n12976), .I2(n12980), .O(n12984) );
  NAND_GATE U13362 ( .I1(n12978), .I2(n12977), .O(n12979) );
  NAND_GATE U13363 ( .I1(n12980), .I2(n12979), .O(n12981) );
  NAND_GATE U13364 ( .I1(n12982), .I2(n12981), .O(n12983) );
  NAND_GATE U13365 ( .I1(n12984), .I2(n12983), .O(n12985) );
  NAND_GATE U13366 ( .I1(n12986), .I2(n12985), .O(n13414) );
  NAND_GATE U13367 ( .I1(n1369), .I2(A[0]), .O(n12987) );
  NAND_GATE U13368 ( .I1(n14781), .I2(n12987), .O(n12988) );
  NAND_GATE U13369 ( .I1(B[6]), .I2(n12988), .O(n12992) );
  NAND_GATE U13370 ( .I1(n1370), .I2(A[1]), .O(n12989) );
  NAND_GATE U13371 ( .I1(n14784), .I2(n12989), .O(n12990) );
  NAND_GATE U13372 ( .I1(B[5]), .I2(n12990), .O(n12991) );
  NAND_GATE U13373 ( .I1(n12992), .I2(n12991), .O(n13426) );
  NAND_GATE U13374 ( .I1(B[4]), .I2(A[2]), .O(n13430) );
  NAND3_GATE U13375 ( .I1(B[4]), .I2(B[5]), .I3(n1196), .O(n13423) );
  NAND_GATE U13376 ( .I1(n13430), .I2(n13423), .O(n12993) );
  NAND_GATE U13377 ( .I1(n13426), .I2(n12993), .O(n12994) );
  INV_GATE U13378 ( .I1(n13430), .O(n13424) );
  INV_GATE U13379 ( .I1(n13423), .O(n13425) );
  NAND_GATE U13380 ( .I1(n13424), .I2(n13425), .O(n13421) );
  NAND_GATE U13381 ( .I1(n12994), .I2(n13421), .O(n13415) );
  NAND_GATE U13382 ( .I1(n13414), .I2(n13415), .O(n12996) );
  NAND_GATE U13383 ( .I1(B[4]), .I2(A[3]), .O(n13416) );
  INV_GATE U13384 ( .I1(n13416), .O(n12995) );
  NAND_GATE U13385 ( .I1(n13414), .I2(n12995), .O(n13411) );
  NAND_GATE U13386 ( .I1(n13415), .I2(n12995), .O(n13410) );
  NAND3_GATE U13387 ( .I1(n12996), .I2(n13411), .I3(n13410), .O(n13400) );
  INV_GATE U13388 ( .I1(n13400), .O(n13397) );
  NAND_GATE U13389 ( .I1(B[4]), .I2(A[4]), .O(n13405) );
  NAND_GATE U13390 ( .I1(n13397), .I2(n13405), .O(n12997) );
  NAND_GATE U13391 ( .I1(n13401), .I2(n12997), .O(n12998) );
  INV_GATE U13392 ( .I1(n13405), .O(n13399) );
  NAND_GATE U13393 ( .I1(n13400), .I2(n13399), .O(n13396) );
  NAND_GATE U13394 ( .I1(n12998), .I2(n13396), .O(n13390) );
  NAND_GATE U13395 ( .I1(n13389), .I2(n13390), .O(n13000) );
  NAND_GATE U13396 ( .I1(B[4]), .I2(A[5]), .O(n13391) );
  INV_GATE U13397 ( .I1(n13391), .O(n12999) );
  NAND_GATE U13398 ( .I1(n13389), .I2(n12999), .O(n13386) );
  NAND_GATE U13399 ( .I1(n13390), .I2(n12999), .O(n13385) );
  NAND3_GATE U13400 ( .I1(n13000), .I2(n13386), .I3(n13385), .O(n13375) );
  INV_GATE U13401 ( .I1(n13375), .O(n13372) );
  NAND_GATE U13402 ( .I1(B[4]), .I2(A[6]), .O(n13380) );
  NAND_GATE U13403 ( .I1(n13372), .I2(n13380), .O(n13001) );
  NAND_GATE U13404 ( .I1(n13376), .I2(n13001), .O(n13002) );
  INV_GATE U13405 ( .I1(n13380), .O(n13374) );
  NAND_GATE U13406 ( .I1(n13375), .I2(n13374), .O(n13371) );
  NAND_GATE U13407 ( .I1(n13002), .I2(n13371), .O(n13365) );
  NAND_GATE U13408 ( .I1(n13364), .I2(n13365), .O(n13004) );
  NAND_GATE U13409 ( .I1(B[4]), .I2(A[7]), .O(n13366) );
  INV_GATE U13410 ( .I1(n13366), .O(n13003) );
  NAND_GATE U13411 ( .I1(n13364), .I2(n13003), .O(n13361) );
  NAND_GATE U13412 ( .I1(n13365), .I2(n13003), .O(n13360) );
  NAND3_GATE U13413 ( .I1(n13004), .I2(n13361), .I3(n13360), .O(n13350) );
  INV_GATE U13414 ( .I1(n13350), .O(n13347) );
  NAND_GATE U13415 ( .I1(B[4]), .I2(A[8]), .O(n13355) );
  NAND_GATE U13416 ( .I1(n13347), .I2(n13355), .O(n13005) );
  NAND_GATE U13417 ( .I1(n13351), .I2(n13005), .O(n13006) );
  INV_GATE U13418 ( .I1(n13355), .O(n13349) );
  NAND_GATE U13419 ( .I1(n13350), .I2(n13349), .O(n13346) );
  NAND_GATE U13420 ( .I1(n13006), .I2(n13346), .O(n13340) );
  NAND_GATE U13421 ( .I1(n13339), .I2(n13340), .O(n13008) );
  NAND_GATE U13422 ( .I1(B[4]), .I2(A[9]), .O(n13341) );
  INV_GATE U13423 ( .I1(n13341), .O(n13007) );
  NAND_GATE U13424 ( .I1(n13339), .I2(n13007), .O(n13336) );
  NAND_GATE U13425 ( .I1(n13340), .I2(n13007), .O(n13335) );
  NAND3_GATE U13426 ( .I1(n13008), .I2(n13336), .I3(n13335), .O(n13325) );
  INV_GATE U13427 ( .I1(n13325), .O(n13322) );
  NAND_GATE U13428 ( .I1(B[4]), .I2(A[10]), .O(n13330) );
  NAND_GATE U13429 ( .I1(n13322), .I2(n13330), .O(n13009) );
  NAND_GATE U13430 ( .I1(n13326), .I2(n13009), .O(n13010) );
  INV_GATE U13431 ( .I1(n13330), .O(n13324) );
  NAND_GATE U13432 ( .I1(n13325), .I2(n13324), .O(n13321) );
  NAND_GATE U13433 ( .I1(n13010), .I2(n13321), .O(n13466) );
  NAND_GATE U13434 ( .I1(n13465), .I2(n13466), .O(n13012) );
  NAND_GATE U13435 ( .I1(B[4]), .I2(A[11]), .O(n13467) );
  INV_GATE U13436 ( .I1(n13467), .O(n13011) );
  NAND_GATE U13437 ( .I1(n13466), .I2(n13011), .O(n13462) );
  NAND_GATE U13438 ( .I1(n13465), .I2(n13011), .O(n13461) );
  NAND3_GATE U13439 ( .I1(n13012), .I2(n13462), .I3(n13461), .O(n13312) );
  NAND_GATE U13440 ( .I1(B[4]), .I2(A[12]), .O(n13316) );
  OR_GATE U13441 ( .I1(n13013), .I2(n13018), .O(n13016) );
  OR_GATE U13442 ( .I1(n13014), .I2(n13017), .O(n13015) );
  AND_GATE U13443 ( .I1(n13016), .I2(n13015), .O(n13023) );
  NAND_GATE U13444 ( .I1(n13017), .I2(n1007), .O(n13021) );
  NAND3_GATE U13445 ( .I1(n13021), .I2(n13020), .I3(n13019), .O(n13022) );
  NAND_GATE U13446 ( .I1(n13023), .I2(n13022), .O(n13308) );
  NAND_GATE U13447 ( .I1(n13316), .I2(n13308), .O(n13024) );
  NAND_GATE U13448 ( .I1(n13312), .I2(n13024), .O(n13025) );
  INV_GATE U13449 ( .I1(n13316), .O(n13310) );
  INV_GATE U13450 ( .I1(n13308), .O(n13311) );
  NAND_GATE U13451 ( .I1(n13310), .I2(n13311), .O(n13306) );
  NAND_GATE U13452 ( .I1(n13025), .I2(n13306), .O(n13481) );
  NAND_GATE U13453 ( .I1(n13480), .I2(n13481), .O(n13027) );
  NAND_GATE U13454 ( .I1(B[4]), .I2(A[13]), .O(n13482) );
  INV_GATE U13455 ( .I1(n13482), .O(n13026) );
  NAND_GATE U13456 ( .I1(n13481), .I2(n13026), .O(n13477) );
  NAND_GATE U13457 ( .I1(n13480), .I2(n13026), .O(n13476) );
  NAND3_GATE U13458 ( .I1(n13027), .I2(n13477), .I3(n13476), .O(n13297) );
  NAND_GATE U13459 ( .I1(B[4]), .I2(A[14]), .O(n13301) );
  OR_GATE U13460 ( .I1(n13028), .I2(n13033), .O(n13031) );
  OR_GATE U13461 ( .I1(n13029), .I2(n13032), .O(n13030) );
  AND_GATE U13462 ( .I1(n13031), .I2(n13030), .O(n13038) );
  NAND_GATE U13463 ( .I1(n13032), .I2(n994), .O(n13036) );
  NAND3_GATE U13464 ( .I1(n13036), .I2(n13035), .I3(n13034), .O(n13037) );
  NAND_GATE U13465 ( .I1(n13038), .I2(n13037), .O(n13293) );
  NAND_GATE U13466 ( .I1(n13301), .I2(n13293), .O(n13039) );
  NAND_GATE U13467 ( .I1(n13297), .I2(n13039), .O(n13040) );
  INV_GATE U13468 ( .I1(n13301), .O(n13295) );
  INV_GATE U13469 ( .I1(n13293), .O(n13296) );
  NAND_GATE U13470 ( .I1(n13295), .I2(n13296), .O(n13291) );
  NAND_GATE U13471 ( .I1(n13040), .I2(n13291), .O(n13495) );
  NAND_GATE U13472 ( .I1(n13494), .I2(n13495), .O(n13042) );
  NAND_GATE U13473 ( .I1(B[4]), .I2(A[15]), .O(n13496) );
  INV_GATE U13474 ( .I1(n13496), .O(n13041) );
  NAND_GATE U13475 ( .I1(n13495), .I2(n13041), .O(n13491) );
  NAND_GATE U13476 ( .I1(n13494), .I2(n13041), .O(n13490) );
  NAND3_GATE U13477 ( .I1(n13042), .I2(n13491), .I3(n13490), .O(n13284) );
  NAND_GATE U13478 ( .I1(B[4]), .I2(A[16]), .O(n13286) );
  OR_GATE U13479 ( .I1(n13043), .I2(n13048), .O(n13046) );
  OR_GATE U13480 ( .I1(n13044), .I2(n13047), .O(n13045) );
  NAND_GATE U13481 ( .I1(n13047), .I2(n932), .O(n13051) );
  NAND3_GATE U13482 ( .I1(n13051), .I2(n13050), .I3(n13049), .O(n13052) );
  NAND_GATE U13483 ( .I1(n13286), .I2(n13280), .O(n13053) );
  NAND_GATE U13484 ( .I1(n13284), .I2(n13053), .O(n13054) );
  INV_GATE U13485 ( .I1(n13286), .O(n13282) );
  INV_GATE U13486 ( .I1(n13280), .O(n13283) );
  NAND_GATE U13487 ( .I1(n13282), .I2(n13283), .O(n13278) );
  NAND_GATE U13488 ( .I1(n13054), .I2(n13278), .O(n13511) );
  NAND_GATE U13489 ( .I1(n13510), .I2(n13511), .O(n13056) );
  NAND_GATE U13490 ( .I1(B[4]), .I2(A[17]), .O(n13512) );
  INV_GATE U13491 ( .I1(n13512), .O(n13055) );
  NAND_GATE U13492 ( .I1(n13511), .I2(n13055), .O(n13506) );
  NAND_GATE U13493 ( .I1(n13510), .I2(n13055), .O(n13505) );
  NAND3_GATE U13494 ( .I1(n13056), .I2(n13506), .I3(n13505), .O(n13271) );
  NAND_GATE U13495 ( .I1(B[4]), .I2(A[18]), .O(n13273) );
  OR_GATE U13496 ( .I1(n13057), .I2(n13062), .O(n13060) );
  OR_GATE U13497 ( .I1(n13058), .I2(n13061), .O(n13059) );
  AND_GATE U13498 ( .I1(n13060), .I2(n13059), .O(n13067) );
  NAND_GATE U13499 ( .I1(n13061), .I2(n960), .O(n13065) );
  NAND3_GATE U13500 ( .I1(n13065), .I2(n13064), .I3(n13063), .O(n13066) );
  NAND_GATE U13501 ( .I1(n13067), .I2(n13066), .O(n13268) );
  NAND_GATE U13502 ( .I1(n13273), .I2(n13268), .O(n13068) );
  NAND_GATE U13503 ( .I1(n13271), .I2(n13068), .O(n13069) );
  INV_GATE U13504 ( .I1(n13273), .O(n13269) );
  INV_GATE U13505 ( .I1(n13268), .O(n13270) );
  NAND_GATE U13506 ( .I1(n13269), .I2(n13270), .O(n13267) );
  NAND_GATE U13507 ( .I1(n13069), .I2(n13267), .O(n13526) );
  NAND_GATE U13508 ( .I1(n13525), .I2(n13526), .O(n13071) );
  NAND_GATE U13509 ( .I1(B[4]), .I2(A[19]), .O(n13527) );
  INV_GATE U13510 ( .I1(n13527), .O(n13070) );
  NAND_GATE U13511 ( .I1(n13526), .I2(n13070), .O(n13522) );
  NAND_GATE U13512 ( .I1(n13525), .I2(n13070), .O(n13521) );
  NAND3_GATE U13513 ( .I1(n13071), .I2(n13522), .I3(n13521), .O(n13261) );
  NAND_GATE U13514 ( .I1(B[4]), .I2(A[20]), .O(n13262) );
  OR_GATE U13515 ( .I1(n13072), .I2(n13077), .O(n13075) );
  OR_GATE U13516 ( .I1(n13073), .I2(n13076), .O(n13074) );
  NAND_GATE U13517 ( .I1(n13076), .I2(n360), .O(n13080) );
  NAND3_GATE U13518 ( .I1(n13080), .I2(n13079), .I3(n13078), .O(n13081) );
  NAND_GATE U13519 ( .I1(n13262), .I2(n13258), .O(n13082) );
  NAND_GATE U13520 ( .I1(n13261), .I2(n13082), .O(n13083) );
  INV_GATE U13521 ( .I1(n13262), .O(n13257) );
  NAND_GATE U13522 ( .I1(n13257), .I2(n13260), .O(n13254) );
  NAND_GATE U13523 ( .I1(n13083), .I2(n13254), .O(n13540) );
  NAND_GATE U13524 ( .I1(n13539), .I2(n13540), .O(n13085) );
  NAND_GATE U13525 ( .I1(B[4]), .I2(A[21]), .O(n13541) );
  INV_GATE U13526 ( .I1(n13541), .O(n13084) );
  NAND_GATE U13527 ( .I1(n13540), .I2(n13084), .O(n13536) );
  NAND_GATE U13528 ( .I1(n13539), .I2(n13084), .O(n13535) );
  NAND3_GATE U13529 ( .I1(n13085), .I2(n13536), .I3(n13535), .O(n13249) );
  NAND_GATE U13530 ( .I1(n13248), .I2(n13250), .O(n13086) );
  NAND_GATE U13531 ( .I1(n13249), .I2(n13086), .O(n13087) );
  NAND_GATE U13532 ( .I1(n13245), .I2(n13087), .O(n13239) );
  NAND_GATE U13533 ( .I1(n13089), .I2(n13094), .O(n13098) );
  NAND_GATE U13534 ( .I1(n13091), .I2(n13090), .O(n13094) );
  NAND_GATE U13535 ( .I1(n1325), .I2(n13092), .O(n13093) );
  NAND_GATE U13536 ( .I1(n13094), .I2(n13093), .O(n13095) );
  NAND_GATE U13537 ( .I1(n13239), .I2(n13238), .O(n13101) );
  NAND3_GATE U13538 ( .I1(n13235), .I2(n13101), .I3(n13234), .O(n13228) );
  NAND_GATE U13539 ( .I1(B[4]), .I2(A[24]), .O(n13231) );
  OR_GATE U13540 ( .I1(n13106), .I2(n13102), .O(n13105) );
  NAND3_GATE U13541 ( .I1(n336), .I2(n13106), .I3(n13103), .O(n13104) );
  AND_GATE U13542 ( .I1(n13105), .I2(n13104), .O(n13111) );
  NAND_GATE U13543 ( .I1(n336), .I2(n13106), .O(n13107) );
  NAND3_GATE U13544 ( .I1(n13109), .I2(n13108), .I3(n13107), .O(n13110) );
  NAND_GATE U13545 ( .I1(n13111), .I2(n13110), .O(n13224) );
  NAND_GATE U13546 ( .I1(n13231), .I2(n13224), .O(n13112) );
  NAND_GATE U13547 ( .I1(n13228), .I2(n13112), .O(n13114) );
  INV_GATE U13548 ( .I1(n13231), .O(n13226) );
  INV_GATE U13549 ( .I1(n13224), .O(n13227) );
  NAND_GATE U13550 ( .I1(n13226), .I2(n13227), .O(n13113) );
  NAND_GATE U13551 ( .I1(n13114), .I2(n13113), .O(n13214) );
  NAND_GATE U13552 ( .I1(n231), .I2(n13124), .O(n13122) );
  NAND_GATE U13553 ( .I1(n13119), .I2(n13118), .O(n13115) );
  NAND_GATE U13554 ( .I1(n13116), .I2(n13115), .O(n13121) );
  NAND3_GATE U13555 ( .I1(n13119), .I2(n13118), .I3(n13117), .O(n13120) );
  NAND3_GATE U13556 ( .I1(n13122), .I2(n13121), .I3(n13120), .O(n13126) );
  NAND_GATE U13557 ( .I1(n13126), .I2(n13125), .O(n13215) );
  NAND_GATE U13558 ( .I1(n13214), .I2(n13215), .O(n13128) );
  NAND_GATE U13559 ( .I1(B[4]), .I2(A[25]), .O(n13220) );
  INV_GATE U13560 ( .I1(n13220), .O(n13127) );
  NAND_GATE U13561 ( .I1(n13127), .I2(n13215), .O(n13213) );
  NAND_GATE U13562 ( .I1(n13127), .I2(n13214), .O(n13216) );
  NAND3_GATE U13563 ( .I1(n13128), .I2(n13213), .I3(n13216), .O(n13210) );
  NAND_GATE U13564 ( .I1(n13203), .I2(n13205), .O(n13129) );
  NAND_GATE U13565 ( .I1(n13210), .I2(n13129), .O(n13130) );
  NAND_GATE U13566 ( .I1(n13209), .I2(n13130), .O(n13194) );
  NAND_GATE U13567 ( .I1(n13194), .I2(n13197), .O(n13131) );
  NAND_GATE U13568 ( .I1(n13196), .I2(n13194), .O(n13195) );
  NAND3_GATE U13569 ( .I1(n13136), .I2(n13135), .I3(n13134), .O(n13137) );
  NAND_GATE U13570 ( .I1(n477), .I2(n523), .O(n13173) );
  NAND_GATE U13571 ( .I1(n13139), .I2(n13173), .O(n13191) );
  NAND_GATE U13572 ( .I1(n13191), .I2(n13175), .O(n13142) );
  NAND3_GATE U13573 ( .I1(n13191), .I2(n13140), .I3(n13188), .O(n13141) );
  NAND3_GATE U13574 ( .I1(n13143), .I2(n13142), .I3(n13141), .O(n13168) );
  NAND_GATE U13575 ( .I1(n13168), .I2(n13154), .O(n13144) );
  NAND_GATE U13576 ( .I1(n13152), .I2(n13168), .O(n13153) );
  NAND3_GATE U13577 ( .I1(n13145), .I2(n13144), .I3(n13153), .O(n13578) );
  NAND_GATE U13578 ( .I1(n13578), .I2(n13577), .O(n13147) );
  NAND_GATE U13579 ( .I1(n13580), .I2(n13578), .O(n13146) );
  NAND3_GATE U13580 ( .I1(n13148), .I2(n13147), .I3(n13146), .O(n15357) );
  INV_GATE U13581 ( .I1(n15357), .O(n13149) );
  NAND_GATE U13582 ( .I1(n15358), .I2(n13149), .O(n13150) );
  NAND_GATE U13583 ( .I1(n13151), .I2(n13150), .O(\A1[34] ) );
  NAND3_GATE U13584 ( .I1(n13152), .I2(n13164), .I3(n13154), .O(n13156) );
  OR_GATE U13585 ( .I1(n13154), .I2(n13153), .O(n13155) );
  NAND_GATE U13586 ( .I1(n624), .I2(n13161), .O(n13162) );
  NAND3_GATE U13587 ( .I1(n13166), .I2(n13164), .I3(n13165), .O(n13170) );
  NAND_GATE U13588 ( .I1(n13166), .I2(n13165), .O(n13167) );
  NAND_GATE U13589 ( .I1(n13168), .I2(n13167), .O(n13169) );
  NAND3_GATE U13590 ( .I1(n13171), .I2(n13170), .I3(n13169), .O(n13172) );
  NAND_GATE U13591 ( .I1(B[3]), .I2(A[31]), .O(n14010) );
  NAND_GATE U13592 ( .I1(B[3]), .I2(A[30]), .O(n13591) );
  INV_GATE U13593 ( .I1(n13591), .O(n13593) );
  OR_GATE U13594 ( .I1(n13569), .I2(n13173), .O(n13177) );
  NAND3_GATE U13595 ( .I1(n467), .I2(n13175), .I3(n13174), .O(n13176) );
  NAND_GATE U13596 ( .I1(n13177), .I2(n13176), .O(n13183) );
  NAND_GATE U13597 ( .I1(n13178), .I2(n12750), .O(n13184) );
  NAND_GATE U13598 ( .I1(n1354), .I2(n13179), .O(n13181) );
  NAND3_GATE U13599 ( .I1(n400), .I2(n13187), .I3(n745), .O(n13180) );
  NAND3_GATE U13600 ( .I1(n13184), .I2(n13181), .I3(n13180), .O(n13182) );
  NAND3_GATE U13601 ( .I1(n13185), .I2(n13183), .I3(n13182), .O(n13571) );
  NAND3_GATE U13602 ( .I1(n13188), .I2(n978), .I3(n512), .O(n13570) );
  NAND_GATE U13603 ( .I1(n13187), .I2(n13186), .O(n13188) );
  NAND3_GATE U13604 ( .I1(n512), .I2(n13189), .I3(n13188), .O(n13567) );
  NAND_GATE U13605 ( .I1(n13189), .I2(n13188), .O(n13190) );
  NAND_GATE U13606 ( .I1(n13191), .I2(n13190), .O(n13568) );
  NAND3_GATE U13607 ( .I1(n13567), .I2(n13568), .I3(n13569), .O(n13589) );
  NAND3_GATE U13608 ( .I1(n13593), .I2(n1201), .I3(n13589), .O(n13587) );
  NAND_GATE U13609 ( .I1(B[3]), .I2(A[29]), .O(n13603) );
  INV_GATE U13610 ( .I1(n13603), .O(n13613) );
  NAND_GATE U13611 ( .I1(n477), .I2(n13192), .O(n13608) );
  NAND3_GATE U13612 ( .I1(n467), .I2(n523), .I3(n477), .O(n13609) );
  NAND_GATE U13613 ( .I1(n467), .I2(n523), .O(n13193) );
  NAND_GATE U13614 ( .I1(n13193), .I2(n13192), .O(n13606) );
  NAND_GATE U13615 ( .I1(n13607), .I2(n13606), .O(n13601) );
  NAND3_GATE U13616 ( .I1(n13613), .I2(n13602), .I3(n13601), .O(n13566) );
  NAND_GATE U13617 ( .I1(B[3]), .I2(A[28]), .O(n13991) );
  NAND_GATE U13618 ( .I1(n452), .I2(n13197), .O(n13560) );
  AND3_GATE U13619 ( .I1(n13560), .I2(n13561), .I3(n13559), .O(n13200) );
  OR_GATE U13620 ( .I1(n13197), .I2(n13195), .O(n13199) );
  NAND3_GATE U13621 ( .I1(n452), .I2(n13197), .I3(n13196), .O(n13198) );
  NAND_GATE U13622 ( .I1(n13199), .I2(n13198), .O(n13558) );
  OR_GATE U13623 ( .I1(n13200), .I2(n13558), .O(n13992) );
  NAND_GATE U13624 ( .I1(n13205), .I2(n13204), .O(n13201) );
  NAND_GATE U13625 ( .I1(n13202), .I2(n13201), .O(n13208) );
  NAND_GATE U13626 ( .I1(n240), .I2(n13210), .O(n13207) );
  NAND3_GATE U13627 ( .I1(n13205), .I2(n13204), .I3(n13203), .O(n13206) );
  NAND3_GATE U13628 ( .I1(n13208), .I2(n13207), .I3(n13206), .O(n13212) );
  NAND_GATE U13629 ( .I1(n13212), .I2(n13211), .O(n13619) );
  NAND3_GATE U13630 ( .I1(n13220), .I2(n13219), .I3(n13218), .O(n13217) );
  NAND3_GATE U13631 ( .I1(n13222), .I2(n13217), .I3(n13221), .O(n13979) );
  NAND_GATE U13632 ( .I1(B[3]), .I2(A[26]), .O(n13975) );
  INV_GATE U13633 ( .I1(n13975), .O(n13981) );
  NAND_GATE U13634 ( .I1(n13977), .I2(n13981), .O(n13974) );
  NAND4_GATE U13635 ( .I1(n13220), .I2(n13219), .I3(n13218), .I4(n13975), .O(
        n13554) );
  NAND_GATE U13636 ( .I1(n13222), .I2(n13221), .O(n13223) );
  NAND_GATE U13637 ( .I1(n13975), .I2(n13223), .O(n13553) );
  NAND_GATE U13638 ( .I1(n13228), .I2(n13227), .O(n13225) );
  NAND3_GATE U13639 ( .I1(n13226), .I2(n13225), .I3(n13229), .O(n13233) );
  NAND_GATE U13640 ( .I1(n13229), .I2(n13225), .O(n13230) );
  NAND_GATE U13641 ( .I1(n13231), .I2(n13230), .O(n13232) );
  OR_GATE U13642 ( .I1(n13234), .I2(n13239), .O(n13237) );
  OR_GATE U13643 ( .I1(n13238), .I2(n13235), .O(n13236) );
  AND_GATE U13644 ( .I1(n13237), .I2(n13236), .O(n13244) );
  NAND_GATE U13645 ( .I1(n372), .I2(n13238), .O(n13242) );
  NAND3_GATE U13646 ( .I1(n13242), .I2(n13241), .I3(n13240), .O(n13243) );
  NAND_GATE U13647 ( .I1(n13244), .I2(n13243), .O(n13633) );
  NAND_GATE U13648 ( .I1(B[3]), .I2(A[24]), .O(n13638) );
  INV_GATE U13649 ( .I1(n13638), .O(n13632) );
  NAND_GATE U13650 ( .I1(n1324), .I2(n13632), .O(n13631) );
  NAND_GATE U13651 ( .I1(n367), .I2(n13249), .O(n13253) );
  NAND_GATE U13652 ( .I1(n13247), .I2(n13246), .O(n13251) );
  NAND_GATE U13653 ( .I1(n13253), .I2(n13252), .O(n13955) );
  INV_GATE U13654 ( .I1(n13254), .O(n13255) );
  NAND_GATE U13655 ( .I1(n13261), .I2(n13255), .O(n13266) );
  NAND_GATE U13656 ( .I1(n13259), .I2(n13258), .O(n13256) );
  NAND_GATE U13657 ( .I1(n13257), .I2(n13256), .O(n13264) );
  NAND_GATE U13658 ( .I1(n13264), .I2(n13263), .O(n13265) );
  NAND_GATE U13659 ( .I1(n13266), .I2(n13265), .O(n13941) );
  NAND_GATE U13660 ( .I1(n13269), .I2(n13272), .O(n13275) );
  NAND_GATE U13661 ( .I1(n13275), .I2(n13274), .O(n13276) );
  NAND_GATE U13662 ( .I1(n13277), .I2(n13276), .O(n13927) );
  INV_GATE U13663 ( .I1(n13278), .O(n13279) );
  NAND_GATE U13664 ( .I1(n13284), .I2(n13279), .O(n13290) );
  INV_GATE U13665 ( .I1(n13284), .O(n13281) );
  NAND_GATE U13666 ( .I1(n13281), .I2(n13280), .O(n13285) );
  NAND_GATE U13667 ( .I1(n13282), .I2(n13285), .O(n13288) );
  NAND_GATE U13668 ( .I1(n13288), .I2(n13287), .O(n13289) );
  NAND_GATE U13669 ( .I1(n13290), .I2(n13289), .O(n13912) );
  INV_GATE U13670 ( .I1(n13291), .O(n13292) );
  NAND_GATE U13671 ( .I1(n13297), .I2(n13292), .O(n13305) );
  INV_GATE U13672 ( .I1(n13297), .O(n13294) );
  NAND_GATE U13673 ( .I1(n13294), .I2(n13293), .O(n13299) );
  NAND_GATE U13674 ( .I1(n13295), .I2(n13299), .O(n13303) );
  NAND_GATE U13675 ( .I1(n13297), .I2(n13296), .O(n13298) );
  NAND_GATE U13676 ( .I1(n13299), .I2(n13298), .O(n13300) );
  NAND_GATE U13677 ( .I1(n13301), .I2(n13300), .O(n13302) );
  NAND_GATE U13678 ( .I1(n13303), .I2(n13302), .O(n13304) );
  NAND_GATE U13679 ( .I1(n13305), .I2(n13304), .O(n13898) );
  INV_GATE U13680 ( .I1(n13306), .O(n13307) );
  NAND_GATE U13681 ( .I1(n13312), .I2(n13307), .O(n13320) );
  INV_GATE U13682 ( .I1(n13312), .O(n13309) );
  NAND_GATE U13683 ( .I1(n13309), .I2(n13308), .O(n13314) );
  NAND_GATE U13684 ( .I1(n13310), .I2(n13314), .O(n13318) );
  NAND_GATE U13685 ( .I1(n13312), .I2(n13311), .O(n13313) );
  NAND_GATE U13686 ( .I1(n13314), .I2(n13313), .O(n13315) );
  NAND_GATE U13687 ( .I1(n13316), .I2(n13315), .O(n13317) );
  NAND_GATE U13688 ( .I1(n13318), .I2(n13317), .O(n13319) );
  NAND_GATE U13689 ( .I1(n13320), .I2(n13319), .O(n13884) );
  OR_GATE U13690 ( .I1(n13321), .I2(n13323), .O(n13334) );
  NAND_GATE U13691 ( .I1(n13323), .I2(n13322), .O(n13328) );
  NAND_GATE U13692 ( .I1(n13324), .I2(n13328), .O(n13332) );
  NAND_GATE U13693 ( .I1(n13326), .I2(n13325), .O(n13327) );
  NAND_GATE U13694 ( .I1(n13328), .I2(n13327), .O(n13329) );
  NAND_GATE U13695 ( .I1(n13330), .I2(n13329), .O(n13331) );
  NAND_GATE U13696 ( .I1(n13332), .I2(n13331), .O(n13333) );
  NAND_GATE U13697 ( .I1(n13334), .I2(n13333), .O(n13869) );
  OR_GATE U13698 ( .I1(n13335), .I2(n13339), .O(n13338) );
  OR_GATE U13699 ( .I1(n13336), .I2(n13340), .O(n13337) );
  AND_GATE U13700 ( .I1(n13338), .I2(n13337), .O(n13345) );
  NAND_GATE U13701 ( .I1(n13339), .I2(n1022), .O(n13343) );
  NAND3_GATE U13702 ( .I1(n13343), .I2(n13342), .I3(n13341), .O(n13344) );
  NAND_GATE U13703 ( .I1(n13345), .I2(n13344), .O(n13727) );
  INV_GATE U13704 ( .I1(n13727), .O(n13730) );
  OR_GATE U13705 ( .I1(n13346), .I2(n13348), .O(n13359) );
  NAND_GATE U13706 ( .I1(n13348), .I2(n13347), .O(n13353) );
  NAND_GATE U13707 ( .I1(n13349), .I2(n13353), .O(n13357) );
  NAND_GATE U13708 ( .I1(n13351), .I2(n13350), .O(n13352) );
  NAND_GATE U13709 ( .I1(n13353), .I2(n13352), .O(n13354) );
  NAND_GATE U13710 ( .I1(n13355), .I2(n13354), .O(n13356) );
  NAND_GATE U13711 ( .I1(n13357), .I2(n13356), .O(n13358) );
  NAND_GATE U13712 ( .I1(n13359), .I2(n13358), .O(n13743) );
  OR_GATE U13713 ( .I1(n13360), .I2(n13364), .O(n13363) );
  OR_GATE U13714 ( .I1(n13361), .I2(n13365), .O(n13362) );
  AND_GATE U13715 ( .I1(n13363), .I2(n13362), .O(n13370) );
  NAND_GATE U13716 ( .I1(n13364), .I2(n1026), .O(n13368) );
  NAND3_GATE U13717 ( .I1(n13368), .I2(n13367), .I3(n13366), .O(n13369) );
  NAND_GATE U13718 ( .I1(n13370), .I2(n13369), .O(n13752) );
  INV_GATE U13719 ( .I1(n13752), .O(n13755) );
  OR_GATE U13720 ( .I1(n13371), .I2(n13373), .O(n13384) );
  NAND_GATE U13721 ( .I1(n13373), .I2(n13372), .O(n13378) );
  NAND_GATE U13722 ( .I1(n13374), .I2(n13378), .O(n13382) );
  NAND_GATE U13723 ( .I1(n13376), .I2(n13375), .O(n13377) );
  NAND_GATE U13724 ( .I1(n13378), .I2(n13377), .O(n13379) );
  NAND_GATE U13725 ( .I1(n13380), .I2(n13379), .O(n13381) );
  NAND_GATE U13726 ( .I1(n13382), .I2(n13381), .O(n13383) );
  NAND_GATE U13727 ( .I1(n13384), .I2(n13383), .O(n13768) );
  OR_GATE U13728 ( .I1(n13385), .I2(n13389), .O(n13388) );
  OR_GATE U13729 ( .I1(n13386), .I2(n13390), .O(n13387) );
  AND_GATE U13730 ( .I1(n13388), .I2(n13387), .O(n13395) );
  NAND_GATE U13731 ( .I1(n13389), .I2(n1118), .O(n13393) );
  NAND3_GATE U13732 ( .I1(n13393), .I2(n13392), .I3(n13391), .O(n13394) );
  NAND_GATE U13733 ( .I1(n13395), .I2(n13394), .O(n13777) );
  INV_GATE U13734 ( .I1(n13777), .O(n13780) );
  OR_GATE U13735 ( .I1(n13396), .I2(n13398), .O(n13409) );
  NAND_GATE U13736 ( .I1(n13398), .I2(n13397), .O(n13403) );
  NAND_GATE U13737 ( .I1(n13399), .I2(n13403), .O(n13407) );
  NAND_GATE U13738 ( .I1(n13401), .I2(n13400), .O(n13402) );
  NAND_GATE U13739 ( .I1(n13403), .I2(n13402), .O(n13404) );
  NAND_GATE U13740 ( .I1(n13405), .I2(n13404), .O(n13406) );
  NAND_GATE U13741 ( .I1(n13407), .I2(n13406), .O(n13408) );
  NAND_GATE U13742 ( .I1(n13409), .I2(n13408), .O(n13793) );
  OR_GATE U13743 ( .I1(n13410), .I2(n13414), .O(n13413) );
  OR_GATE U13744 ( .I1(n13411), .I2(n13415), .O(n13412) );
  AND_GATE U13745 ( .I1(n13413), .I2(n13412), .O(n13420) );
  NAND_GATE U13746 ( .I1(n13414), .I2(n1188), .O(n13418) );
  NAND3_GATE U13747 ( .I1(n13418), .I2(n13417), .I3(n13416), .O(n13419) );
  NAND_GATE U13748 ( .I1(n13420), .I2(n13419), .O(n13802) );
  INV_GATE U13749 ( .I1(n13802), .O(n13805) );
  INV_GATE U13750 ( .I1(n13421), .O(n13422) );
  NAND_GATE U13751 ( .I1(n13426), .I2(n13422), .O(n13434) );
  NAND_GATE U13752 ( .I1(n13424), .I2(n13428), .O(n13432) );
  NAND_GATE U13753 ( .I1(n13426), .I2(n13425), .O(n13427) );
  NAND_GATE U13754 ( .I1(n13428), .I2(n13427), .O(n13429) );
  NAND_GATE U13755 ( .I1(n13430), .I2(n13429), .O(n13431) );
  NAND_GATE U13756 ( .I1(n13432), .I2(n13431), .O(n13433) );
  NAND_GATE U13757 ( .I1(n13434), .I2(n13433), .O(n13818) );
  NAND_GATE U13758 ( .I1(n1368), .I2(A[0]), .O(n13435) );
  NAND_GATE U13759 ( .I1(n14781), .I2(n13435), .O(n13436) );
  NAND_GATE U13760 ( .I1(B[5]), .I2(n13436), .O(n13440) );
  NAND_GATE U13761 ( .I1(n1369), .I2(A[1]), .O(n13437) );
  NAND_GATE U13762 ( .I1(n14784), .I2(n13437), .O(n13438) );
  NAND_GATE U13763 ( .I1(B[4]), .I2(n13438), .O(n13439) );
  NAND_GATE U13764 ( .I1(n13440), .I2(n13439), .O(n13830) );
  NAND_GATE U13765 ( .I1(B[3]), .I2(A[2]), .O(n13834) );
  NAND3_GATE U13766 ( .I1(B[3]), .I2(B[4]), .I3(n1196), .O(n13827) );
  NAND_GATE U13767 ( .I1(n13834), .I2(n13827), .O(n13441) );
  NAND_GATE U13768 ( .I1(n13830), .I2(n13441), .O(n13442) );
  INV_GATE U13769 ( .I1(n13834), .O(n13828) );
  INV_GATE U13770 ( .I1(n13827), .O(n13829) );
  NAND_GATE U13771 ( .I1(n13828), .I2(n13829), .O(n13825) );
  NAND_GATE U13772 ( .I1(n13442), .I2(n13825), .O(n13819) );
  NAND_GATE U13773 ( .I1(n13818), .I2(n13819), .O(n13444) );
  NAND_GATE U13774 ( .I1(B[3]), .I2(A[3]), .O(n13820) );
  INV_GATE U13775 ( .I1(n13820), .O(n13443) );
  NAND_GATE U13776 ( .I1(n13818), .I2(n13443), .O(n13815) );
  NAND_GATE U13777 ( .I1(n13819), .I2(n13443), .O(n13814) );
  NAND3_GATE U13778 ( .I1(n13444), .I2(n13815), .I3(n13814), .O(n13804) );
  INV_GATE U13779 ( .I1(n13804), .O(n13801) );
  NAND_GATE U13780 ( .I1(B[3]), .I2(A[4]), .O(n13809) );
  NAND_GATE U13781 ( .I1(n13801), .I2(n13809), .O(n13445) );
  NAND_GATE U13782 ( .I1(n13805), .I2(n13445), .O(n13446) );
  INV_GATE U13783 ( .I1(n13809), .O(n13803) );
  NAND_GATE U13784 ( .I1(n13804), .I2(n13803), .O(n13800) );
  NAND_GATE U13785 ( .I1(n13446), .I2(n13800), .O(n13794) );
  NAND_GATE U13786 ( .I1(n13793), .I2(n13794), .O(n13448) );
  NAND_GATE U13787 ( .I1(B[3]), .I2(A[5]), .O(n13795) );
  INV_GATE U13788 ( .I1(n13795), .O(n13447) );
  NAND_GATE U13789 ( .I1(n13793), .I2(n13447), .O(n13790) );
  NAND_GATE U13790 ( .I1(n13794), .I2(n13447), .O(n13789) );
  NAND3_GATE U13791 ( .I1(n13448), .I2(n13790), .I3(n13789), .O(n13779) );
  INV_GATE U13792 ( .I1(n13779), .O(n13776) );
  NAND_GATE U13793 ( .I1(B[3]), .I2(A[6]), .O(n13784) );
  NAND_GATE U13794 ( .I1(n13776), .I2(n13784), .O(n13449) );
  NAND_GATE U13795 ( .I1(n13780), .I2(n13449), .O(n13450) );
  INV_GATE U13796 ( .I1(n13784), .O(n13778) );
  NAND_GATE U13797 ( .I1(n13779), .I2(n13778), .O(n13775) );
  NAND_GATE U13798 ( .I1(n13450), .I2(n13775), .O(n13769) );
  NAND_GATE U13799 ( .I1(n13768), .I2(n13769), .O(n13452) );
  NAND_GATE U13800 ( .I1(B[3]), .I2(A[7]), .O(n13770) );
  INV_GATE U13801 ( .I1(n13770), .O(n13451) );
  NAND_GATE U13802 ( .I1(n13768), .I2(n13451), .O(n13765) );
  NAND_GATE U13803 ( .I1(n13769), .I2(n13451), .O(n13764) );
  NAND3_GATE U13804 ( .I1(n13452), .I2(n13765), .I3(n13764), .O(n13754) );
  INV_GATE U13805 ( .I1(n13754), .O(n13751) );
  NAND_GATE U13806 ( .I1(B[3]), .I2(A[8]), .O(n13759) );
  NAND_GATE U13807 ( .I1(n13751), .I2(n13759), .O(n13453) );
  NAND_GATE U13808 ( .I1(n13755), .I2(n13453), .O(n13454) );
  INV_GATE U13809 ( .I1(n13759), .O(n13753) );
  NAND_GATE U13810 ( .I1(n13754), .I2(n13753), .O(n13750) );
  NAND_GATE U13811 ( .I1(n13454), .I2(n13750), .O(n13744) );
  NAND_GATE U13812 ( .I1(n13743), .I2(n13744), .O(n13456) );
  NAND_GATE U13813 ( .I1(B[3]), .I2(A[9]), .O(n13745) );
  INV_GATE U13814 ( .I1(n13745), .O(n13455) );
  NAND_GATE U13815 ( .I1(n13743), .I2(n13455), .O(n13740) );
  NAND_GATE U13816 ( .I1(n13744), .I2(n13455), .O(n13739) );
  NAND3_GATE U13817 ( .I1(n13456), .I2(n13740), .I3(n13739), .O(n13729) );
  INV_GATE U13818 ( .I1(n13729), .O(n13726) );
  NAND_GATE U13819 ( .I1(B[3]), .I2(A[10]), .O(n13734) );
  NAND_GATE U13820 ( .I1(n13726), .I2(n13734), .O(n13457) );
  NAND_GATE U13821 ( .I1(n13730), .I2(n13457), .O(n13458) );
  INV_GATE U13822 ( .I1(n13734), .O(n13728) );
  NAND_GATE U13823 ( .I1(n13729), .I2(n13728), .O(n13725) );
  NAND_GATE U13824 ( .I1(n13458), .I2(n13725), .O(n13870) );
  NAND_GATE U13825 ( .I1(n13869), .I2(n13870), .O(n13460) );
  NAND_GATE U13826 ( .I1(B[3]), .I2(A[11]), .O(n13871) );
  INV_GATE U13827 ( .I1(n13871), .O(n13459) );
  NAND_GATE U13828 ( .I1(n13870), .I2(n13459), .O(n13866) );
  NAND_GATE U13829 ( .I1(n13869), .I2(n13459), .O(n13865) );
  NAND3_GATE U13830 ( .I1(n13460), .I2(n13866), .I3(n13865), .O(n13716) );
  NAND_GATE U13831 ( .I1(B[3]), .I2(A[12]), .O(n13720) );
  OR_GATE U13832 ( .I1(n13461), .I2(n13466), .O(n13464) );
  OR_GATE U13833 ( .I1(n13462), .I2(n13465), .O(n13463) );
  AND_GATE U13834 ( .I1(n13464), .I2(n13463), .O(n13471) );
  NAND_GATE U13835 ( .I1(n13465), .I2(n1012), .O(n13469) );
  NAND3_GATE U13836 ( .I1(n13469), .I2(n13468), .I3(n13467), .O(n13470) );
  NAND_GATE U13837 ( .I1(n13471), .I2(n13470), .O(n13712) );
  NAND_GATE U13838 ( .I1(n13720), .I2(n13712), .O(n13472) );
  NAND_GATE U13839 ( .I1(n13716), .I2(n13472), .O(n13473) );
  INV_GATE U13840 ( .I1(n13720), .O(n13714) );
  INV_GATE U13841 ( .I1(n13712), .O(n13715) );
  NAND_GATE U13842 ( .I1(n13714), .I2(n13715), .O(n13710) );
  NAND_GATE U13843 ( .I1(n13473), .I2(n13710), .O(n13885) );
  NAND_GATE U13844 ( .I1(n13884), .I2(n13885), .O(n13475) );
  NAND_GATE U13845 ( .I1(B[3]), .I2(A[13]), .O(n13886) );
  INV_GATE U13846 ( .I1(n13886), .O(n13474) );
  NAND_GATE U13847 ( .I1(n13885), .I2(n13474), .O(n13881) );
  NAND_GATE U13848 ( .I1(n13884), .I2(n13474), .O(n13880) );
  NAND3_GATE U13849 ( .I1(n13475), .I2(n13881), .I3(n13880), .O(n13701) );
  NAND_GATE U13850 ( .I1(B[3]), .I2(A[14]), .O(n13705) );
  OR_GATE U13851 ( .I1(n13476), .I2(n13481), .O(n13479) );
  OR_GATE U13852 ( .I1(n13477), .I2(n13480), .O(n13478) );
  NAND_GATE U13853 ( .I1(n13480), .I2(n1002), .O(n13484) );
  NAND3_GATE U13854 ( .I1(n13484), .I2(n13483), .I3(n13482), .O(n13485) );
  NAND_GATE U13855 ( .I1(n13705), .I2(n13697), .O(n13486) );
  NAND_GATE U13856 ( .I1(n13701), .I2(n13486), .O(n13487) );
  INV_GATE U13857 ( .I1(n13705), .O(n13699) );
  INV_GATE U13858 ( .I1(n13697), .O(n13700) );
  NAND_GATE U13859 ( .I1(n13699), .I2(n13700), .O(n13695) );
  NAND_GATE U13860 ( .I1(n13487), .I2(n13695), .O(n13899) );
  NAND_GATE U13861 ( .I1(n13898), .I2(n13899), .O(n13489) );
  NAND_GATE U13862 ( .I1(B[3]), .I2(A[15]), .O(n13900) );
  INV_GATE U13863 ( .I1(n13900), .O(n13488) );
  NAND_GATE U13864 ( .I1(n13899), .I2(n13488), .O(n13895) );
  NAND_GATE U13865 ( .I1(n13898), .I2(n13488), .O(n13894) );
  NAND3_GATE U13866 ( .I1(n13489), .I2(n13895), .I3(n13894), .O(n13686) );
  NAND_GATE U13867 ( .I1(B[3]), .I2(A[16]), .O(n13690) );
  OR_GATE U13868 ( .I1(n13490), .I2(n13495), .O(n13493) );
  OR_GATE U13869 ( .I1(n13491), .I2(n13494), .O(n13492) );
  AND_GATE U13870 ( .I1(n13493), .I2(n13492), .O(n13500) );
  NAND_GATE U13871 ( .I1(n13494), .I2(n963), .O(n13498) );
  NAND3_GATE U13872 ( .I1(n13498), .I2(n13497), .I3(n13496), .O(n13499) );
  NAND_GATE U13873 ( .I1(n13500), .I2(n13499), .O(n13682) );
  NAND_GATE U13874 ( .I1(n13690), .I2(n13682), .O(n13501) );
  NAND_GATE U13875 ( .I1(n13686), .I2(n13501), .O(n13502) );
  INV_GATE U13876 ( .I1(n13690), .O(n13684) );
  INV_GATE U13877 ( .I1(n13682), .O(n13685) );
  NAND_GATE U13878 ( .I1(n13684), .I2(n13685), .O(n13680) );
  NAND_GATE U13879 ( .I1(n13502), .I2(n13680), .O(n13913) );
  NAND_GATE U13880 ( .I1(n13912), .I2(n13913), .O(n13504) );
  NAND_GATE U13881 ( .I1(B[3]), .I2(A[17]), .O(n13914) );
  INV_GATE U13882 ( .I1(n13914), .O(n13503) );
  NAND_GATE U13883 ( .I1(n13913), .I2(n13503), .O(n13909) );
  NAND_GATE U13884 ( .I1(n13912), .I2(n13503), .O(n13908) );
  NAND3_GATE U13885 ( .I1(n13504), .I2(n13909), .I3(n13908), .O(n13672) );
  NAND_GATE U13886 ( .I1(B[3]), .I2(A[18]), .O(n13675) );
  OR_GATE U13887 ( .I1(n13506), .I2(n13510), .O(n13507) );
  AND_GATE U13888 ( .I1(n13508), .I2(n13507), .O(n13516) );
  INV_GATE U13889 ( .I1(n13511), .O(n13509) );
  NAND_GATE U13890 ( .I1(n13510), .I2(n13509), .O(n13514) );
  NAND_GATE U13891 ( .I1(n1284), .I2(n13511), .O(n13513) );
  NAND3_GATE U13892 ( .I1(n13514), .I2(n13513), .I3(n13512), .O(n13515) );
  NAND_GATE U13893 ( .I1(n13516), .I2(n13515), .O(n13670) );
  NAND_GATE U13894 ( .I1(n13675), .I2(n13670), .O(n13517) );
  NAND_GATE U13895 ( .I1(n13672), .I2(n13517), .O(n13518) );
  INV_GATE U13896 ( .I1(n13675), .O(n13671) );
  NAND_GATE U13897 ( .I1(n13671), .I2(n50), .O(n13669) );
  NAND_GATE U13898 ( .I1(n13518), .I2(n13669), .O(n13928) );
  NAND_GATE U13899 ( .I1(n13927), .I2(n13928), .O(n13520) );
  NAND_GATE U13900 ( .I1(B[3]), .I2(A[19]), .O(n13929) );
  INV_GATE U13901 ( .I1(n13929), .O(n13519) );
  NAND3_GATE U13902 ( .I1(n13520), .I2(n13924), .I3(n13923), .O(n13660) );
  NAND_GATE U13903 ( .I1(B[3]), .I2(A[20]), .O(n13664) );
  OR_GATE U13904 ( .I1(n13521), .I2(n13526), .O(n13524) );
  OR_GATE U13905 ( .I1(n13522), .I2(n13525), .O(n13523) );
  NAND_GATE U13906 ( .I1(n13525), .I2(n927), .O(n13529) );
  NAND3_GATE U13907 ( .I1(n13529), .I2(n13528), .I3(n13527), .O(n13530) );
  NAND_GATE U13908 ( .I1(n13664), .I2(n13656), .O(n13531) );
  NAND_GATE U13909 ( .I1(n13660), .I2(n13531), .O(n13532) );
  INV_GATE U13910 ( .I1(n13664), .O(n13658) );
  INV_GATE U13911 ( .I1(n13656), .O(n13659) );
  NAND_GATE U13912 ( .I1(n13658), .I2(n13659), .O(n13654) );
  NAND_GATE U13913 ( .I1(n13532), .I2(n13654), .O(n13942) );
  NAND_GATE U13914 ( .I1(n13941), .I2(n13942), .O(n13534) );
  NAND_GATE U13915 ( .I1(B[3]), .I2(A[21]), .O(n13943) );
  INV_GATE U13916 ( .I1(n13943), .O(n13533) );
  NAND_GATE U13917 ( .I1(n13942), .I2(n13533), .O(n13938) );
  NAND_GATE U13918 ( .I1(n13941), .I2(n13533), .O(n13937) );
  NAND3_GATE U13919 ( .I1(n13534), .I2(n13938), .I3(n13937), .O(n13648) );
  NAND_GATE U13920 ( .I1(B[3]), .I2(A[22]), .O(n13649) );
  OR_GATE U13921 ( .I1(n13535), .I2(n13540), .O(n13538) );
  OR_GATE U13922 ( .I1(n13536), .I2(n13539), .O(n13537) );
  NAND_GATE U13923 ( .I1(n13539), .I2(n923), .O(n13543) );
  NAND3_GATE U13924 ( .I1(n13543), .I2(n13542), .I3(n13541), .O(n13544) );
  NAND_GATE U13925 ( .I1(n13649), .I2(n13645), .O(n13545) );
  NAND_GATE U13926 ( .I1(n13648), .I2(n13545), .O(n13546) );
  INV_GATE U13927 ( .I1(n13649), .O(n13644) );
  NAND_GATE U13928 ( .I1(n13644), .I2(n13647), .O(n13641) );
  NAND_GATE U13929 ( .I1(n13546), .I2(n13641), .O(n13956) );
  NAND_GATE U13930 ( .I1(n13955), .I2(n13956), .O(n13548) );
  NAND_GATE U13931 ( .I1(B[3]), .I2(A[23]), .O(n13957) );
  INV_GATE U13932 ( .I1(n13957), .O(n13547) );
  NAND_GATE U13933 ( .I1(n13956), .I2(n13547), .O(n13952) );
  NAND_GATE U13934 ( .I1(n13955), .I2(n13547), .O(n13951) );
  NAND_GATE U13935 ( .I1(n13633), .I2(n13638), .O(n13549) );
  NAND_GATE U13936 ( .I1(n13634), .I2(n13549), .O(n13550) );
  NAND_GATE U13937 ( .I1(n13631), .I2(n13550), .O(n13626) );
  NAND_GATE U13938 ( .I1(B[3]), .I2(A[25]), .O(n13969) );
  INV_GATE U13939 ( .I1(n13969), .O(n13551) );
  NAND_GATE U13940 ( .I1(n13551), .I2(n13626), .O(n13629) );
  NAND3_GATE U13941 ( .I1(n13552), .I2(n13629), .I3(n13627), .O(n13976) );
  NAND3_GATE U13942 ( .I1(n13554), .I2(n13553), .I3(n13976), .O(n13555) );
  NAND_GATE U13943 ( .I1(n13974), .I2(n13555), .O(n13622) );
  NAND_GATE U13944 ( .I1(n13619), .I2(n13622), .O(n13557) );
  NAND_GATE U13945 ( .I1(B[3]), .I2(A[27]), .O(n13616) );
  INV_GATE U13946 ( .I1(n13616), .O(n13556) );
  NAND_GATE U13947 ( .I1(n13556), .I2(n13622), .O(n13620) );
  NAND_GATE U13948 ( .I1(n13556), .I2(n13619), .O(n13621) );
  NAND3_GATE U13949 ( .I1(n13557), .I2(n13620), .I3(n13621), .O(n13997) );
  NAND4_GATE U13950 ( .I1(n13561), .I2(n13991), .I3(n13560), .I4(n13559), .O(
        n13562) );
  NAND3_GATE U13951 ( .I1(n13997), .I2(n13563), .I3(n13562), .O(n13564) );
  NAND_GATE U13952 ( .I1(n13996), .I2(n13564), .O(n13600) );
  NAND3_GATE U13953 ( .I1(n13602), .I2(n13601), .I3(n13600), .O(n13565) );
  NAND_GATE U13954 ( .I1(n13613), .I2(n13600), .O(n13610) );
  NAND3_GATE U13955 ( .I1(n13566), .I2(n13565), .I3(n13610), .O(n13590) );
  NAND4_GATE U13956 ( .I1(n13569), .I2(n13591), .I3(n13568), .I4(n13567), .O(
        n13574) );
  NAND_GATE U13957 ( .I1(n13571), .I2(n13570), .O(n13572) );
  NAND_GATE U13958 ( .I1(n13591), .I2(n13572), .O(n13573) );
  NAND3_GATE U13959 ( .I1(n13590), .I2(n13574), .I3(n13573), .O(n13575) );
  NAND_GATE U13960 ( .I1(n13587), .I2(n13575), .O(n14016) );
  NAND_GATE U13961 ( .I1(n14012), .I2(n14010), .O(n13576) );
  INV_GATE U13962 ( .I1(n13578), .O(n13579) );
  NAND3_GATE U13963 ( .I1(n13577), .I2(n13579), .I3(n13580), .O(n15362) );
  NAND3_GATE U13964 ( .I1(n13578), .I2(n13577), .I3(n606), .O(n15361) );
  NAND_GATE U13965 ( .I1(n457), .I2(n12744), .O(n13583) );
  NAND_GATE U13966 ( .I1(n13580), .I2(n13579), .O(n13582) );
  NAND3_GATE U13967 ( .I1(n13583), .I2(n13582), .I3(n13581), .O(n15360) );
  NAND3_GATE U13968 ( .I1(n15362), .I2(n15361), .I3(n15360), .O(n13584) );
  NAND_GATE U13969 ( .I1(n1265), .I2(n13584), .O(n13586) );
  AND_GATE U13970 ( .I1(n13586), .I2(n13585), .O(\A1[33] ) );
  NAND_GATE U13971 ( .I1(n1365), .I2(A[31]), .O(n14450) );
  INV_GATE U13972 ( .I1(n14450), .O(n14445) );
  INV_GATE U13973 ( .I1(n13587), .O(n13588) );
  NAND_GATE U13974 ( .I1(n13588), .I2(n13590), .O(n13598) );
  NAND_GATE U13975 ( .I1(n1201), .I2(n13589), .O(n13592) );
  NAND3_GATE U13976 ( .I1(n13591), .I2(n514), .I3(n13592), .O(n13595) );
  NAND3_GATE U13977 ( .I1(n13596), .I2(n13595), .I3(n13594), .O(n13597) );
  NAND_GATE U13978 ( .I1(n13598), .I2(n13597), .O(n14449) );
  NAND_GATE U13979 ( .I1(n14445), .I2(n14449), .O(n14009) );
  NAND_GATE U13980 ( .I1(n13601), .I2(n13602), .O(n13599) );
  NAND_GATE U13981 ( .I1(n13600), .I2(n13599), .O(n13605) );
  NAND3_GATE U13982 ( .I1(n13612), .I2(n13602), .I3(n13601), .O(n13604) );
  NAND3_GATE U13983 ( .I1(n13605), .I2(n13604), .I3(n13603), .O(n14003) );
  OR_GATE U13984 ( .I1(n13611), .I2(n13610), .O(n13615) );
  NAND3_GATE U13985 ( .I1(n13613), .I2(n13612), .I3(n13611), .O(n13614) );
  AND_GATE U13986 ( .I1(n13615), .I2(n13614), .O(n14004) );
  NAND_GATE U13987 ( .I1(n1365), .I2(A[30]), .O(n14021) );
  INV_GATE U13988 ( .I1(n14021), .O(n14023) );
  NAND3_GATE U13989 ( .I1(n14003), .I2(n14004), .I3(n14023), .O(n14027) );
  NAND_GATE U13990 ( .I1(n13619), .I2(n401), .O(n13618) );
  NAND3_GATE U13991 ( .I1(n13618), .I2(n13617), .I3(n13616), .O(n13625) );
  OR_GATE U13992 ( .I1(n13620), .I2(n13619), .O(n13624) );
  OR_GATE U13993 ( .I1(n13622), .I2(n13621), .O(n13623) );
  NAND3_GATE U13994 ( .I1(n13625), .I2(n13624), .I3(n13623), .O(n14430) );
  INV_GATE U13995 ( .I1(n14430), .O(n14426) );
  NAND_GATE U13996 ( .I1(n1365), .I2(A[28]), .O(n14428) );
  INV_GATE U13997 ( .I1(n14428), .O(n14432) );
  INV_GATE U13998 ( .I1(n13626), .O(n13628) );
  NAND_GATE U13999 ( .I1(n1264), .I2(n13628), .O(n13967) );
  NAND_GATE U14000 ( .I1(n1365), .I2(A[26]), .O(n14412) );
  NAND4_GATE U14001 ( .I1(n13969), .I2(n13968), .I3(n13967), .I4(n14412), .O(
        n13966) );
  NAND_GATE U14002 ( .I1(n13632), .I2(n13636), .O(n13639) );
  NAND_GATE U14003 ( .I1(n13633), .I2(n734), .O(n13636) );
  NAND_GATE U14004 ( .I1(n1324), .I2(n13634), .O(n13635) );
  NAND_GATE U14005 ( .I1(n13636), .I2(n13635), .O(n13637) );
  INV_GATE U14006 ( .I1(n13641), .O(n13642) );
  NAND_GATE U14007 ( .I1(n13648), .I2(n13642), .O(n13653) );
  NAND_GATE U14008 ( .I1(n13646), .I2(n13645), .O(n13643) );
  NAND_GATE U14009 ( .I1(n13644), .I2(n13643), .O(n13651) );
  NAND_GATE U14010 ( .I1(n13651), .I2(n13650), .O(n13652) );
  NAND_GATE U14011 ( .I1(n13653), .I2(n13652), .O(n14394) );
  INV_GATE U14012 ( .I1(n13654), .O(n13655) );
  NAND_GATE U14013 ( .I1(n13660), .I2(n13655), .O(n13668) );
  INV_GATE U14014 ( .I1(n13660), .O(n13657) );
  NAND_GATE U14015 ( .I1(n13657), .I2(n13656), .O(n13662) );
  NAND_GATE U14016 ( .I1(n13658), .I2(n13662), .O(n13666) );
  NAND_GATE U14017 ( .I1(n13660), .I2(n13659), .O(n13661) );
  NAND_GATE U14018 ( .I1(n13662), .I2(n13661), .O(n13663) );
  NAND_GATE U14019 ( .I1(n13664), .I2(n13663), .O(n13665) );
  NAND_GATE U14020 ( .I1(n13666), .I2(n13665), .O(n13667) );
  NAND_GATE U14021 ( .I1(n13668), .I2(n13667), .O(n14379) );
  NAND_GATE U14022 ( .I1(n13671), .I2(n13674), .O(n13677) );
  NAND_GATE U14023 ( .I1(n13672), .I2(n50), .O(n13673) );
  NAND_GATE U14024 ( .I1(n13677), .I2(n13676), .O(n13678) );
  NAND_GATE U14025 ( .I1(n13679), .I2(n13678), .O(n14365) );
  INV_GATE U14026 ( .I1(n13680), .O(n13681) );
  NAND_GATE U14027 ( .I1(n13686), .I2(n13681), .O(n13694) );
  INV_GATE U14028 ( .I1(n13686), .O(n13683) );
  NAND_GATE U14029 ( .I1(n13683), .I2(n13682), .O(n13688) );
  NAND_GATE U14030 ( .I1(n13684), .I2(n13688), .O(n13692) );
  NAND_GATE U14031 ( .I1(n13686), .I2(n13685), .O(n13687) );
  NAND_GATE U14032 ( .I1(n13688), .I2(n13687), .O(n13689) );
  NAND_GATE U14033 ( .I1(n13690), .I2(n13689), .O(n13691) );
  NAND_GATE U14034 ( .I1(n13692), .I2(n13691), .O(n13693) );
  NAND_GATE U14035 ( .I1(n13694), .I2(n13693), .O(n14349) );
  INV_GATE U14036 ( .I1(n13695), .O(n13696) );
  NAND_GATE U14037 ( .I1(n13701), .I2(n13696), .O(n13709) );
  INV_GATE U14038 ( .I1(n13701), .O(n13698) );
  NAND_GATE U14039 ( .I1(n13698), .I2(n13697), .O(n13703) );
  NAND_GATE U14040 ( .I1(n13699), .I2(n13703), .O(n13707) );
  NAND_GATE U14041 ( .I1(n13701), .I2(n13700), .O(n13702) );
  NAND_GATE U14042 ( .I1(n13703), .I2(n13702), .O(n13704) );
  NAND_GATE U14043 ( .I1(n13705), .I2(n13704), .O(n13706) );
  NAND_GATE U14044 ( .I1(n13707), .I2(n13706), .O(n13708) );
  NAND_GATE U14045 ( .I1(n13709), .I2(n13708), .O(n14335) );
  INV_GATE U14046 ( .I1(n13710), .O(n13711) );
  NAND_GATE U14047 ( .I1(n13716), .I2(n13711), .O(n13724) );
  INV_GATE U14048 ( .I1(n13716), .O(n13713) );
  NAND_GATE U14049 ( .I1(n13713), .I2(n13712), .O(n13718) );
  NAND_GATE U14050 ( .I1(n13714), .I2(n13718), .O(n13722) );
  NAND_GATE U14051 ( .I1(n13716), .I2(n13715), .O(n13717) );
  NAND_GATE U14052 ( .I1(n13718), .I2(n13717), .O(n13719) );
  NAND_GATE U14053 ( .I1(n13720), .I2(n13719), .O(n13721) );
  NAND_GATE U14054 ( .I1(n13722), .I2(n13721), .O(n13723) );
  NAND_GATE U14055 ( .I1(n13724), .I2(n13723), .O(n14320) );
  OR_GATE U14056 ( .I1(n13725), .I2(n13727), .O(n13738) );
  NAND_GATE U14057 ( .I1(n13727), .I2(n13726), .O(n13732) );
  NAND_GATE U14058 ( .I1(n13728), .I2(n13732), .O(n13736) );
  NAND_GATE U14059 ( .I1(n13730), .I2(n13729), .O(n13731) );
  NAND_GATE U14060 ( .I1(n13732), .I2(n13731), .O(n13733) );
  NAND_GATE U14061 ( .I1(n13734), .I2(n13733), .O(n13735) );
  NAND_GATE U14062 ( .I1(n13736), .I2(n13735), .O(n13737) );
  NAND_GATE U14063 ( .I1(n13738), .I2(n13737), .O(n14305) );
  OR_GATE U14064 ( .I1(n13739), .I2(n13743), .O(n13742) );
  OR_GATE U14065 ( .I1(n13740), .I2(n13744), .O(n13741) );
  AND_GATE U14066 ( .I1(n13742), .I2(n13741), .O(n13749) );
  NAND_GATE U14067 ( .I1(n13743), .I2(n1024), .O(n13747) );
  NAND3_GATE U14068 ( .I1(n13747), .I2(n13746), .I3(n13745), .O(n13748) );
  NAND_GATE U14069 ( .I1(n13749), .I2(n13748), .O(n14163) );
  INV_GATE U14070 ( .I1(n14163), .O(n14166) );
  OR_GATE U14071 ( .I1(n13750), .I2(n13752), .O(n13763) );
  NAND_GATE U14072 ( .I1(n13752), .I2(n13751), .O(n13757) );
  NAND_GATE U14073 ( .I1(n13753), .I2(n13757), .O(n13761) );
  NAND_GATE U14074 ( .I1(n13755), .I2(n13754), .O(n13756) );
  NAND_GATE U14075 ( .I1(n13757), .I2(n13756), .O(n13758) );
  NAND_GATE U14076 ( .I1(n13759), .I2(n13758), .O(n13760) );
  NAND_GATE U14077 ( .I1(n13761), .I2(n13760), .O(n13762) );
  NAND_GATE U14078 ( .I1(n13763), .I2(n13762), .O(n14179) );
  OR_GATE U14079 ( .I1(n13764), .I2(n13768), .O(n13767) );
  OR_GATE U14080 ( .I1(n13765), .I2(n13769), .O(n13766) );
  AND_GATE U14081 ( .I1(n13767), .I2(n13766), .O(n13774) );
  NAND_GATE U14082 ( .I1(n13768), .I2(n1028), .O(n13772) );
  NAND3_GATE U14083 ( .I1(n13772), .I2(n13771), .I3(n13770), .O(n13773) );
  NAND_GATE U14084 ( .I1(n13774), .I2(n13773), .O(n14188) );
  INV_GATE U14085 ( .I1(n14188), .O(n14191) );
  OR_GATE U14086 ( .I1(n13775), .I2(n13777), .O(n13788) );
  NAND_GATE U14087 ( .I1(n13777), .I2(n13776), .O(n13782) );
  NAND_GATE U14088 ( .I1(n13778), .I2(n13782), .O(n13786) );
  NAND_GATE U14089 ( .I1(n13780), .I2(n13779), .O(n13781) );
  NAND_GATE U14090 ( .I1(n13782), .I2(n13781), .O(n13783) );
  NAND_GATE U14091 ( .I1(n13784), .I2(n13783), .O(n13785) );
  NAND_GATE U14092 ( .I1(n13786), .I2(n13785), .O(n13787) );
  NAND_GATE U14093 ( .I1(n13788), .I2(n13787), .O(n14204) );
  OR_GATE U14094 ( .I1(n13789), .I2(n13793), .O(n13792) );
  OR_GATE U14095 ( .I1(n13790), .I2(n13794), .O(n13791) );
  AND_GATE U14096 ( .I1(n13792), .I2(n13791), .O(n13799) );
  NAND_GATE U14097 ( .I1(n13793), .I2(n1120), .O(n13797) );
  NAND3_GATE U14098 ( .I1(n13797), .I2(n13796), .I3(n13795), .O(n13798) );
  NAND_GATE U14099 ( .I1(n13799), .I2(n13798), .O(n14213) );
  INV_GATE U14100 ( .I1(n14213), .O(n14216) );
  OR_GATE U14101 ( .I1(n13800), .I2(n13802), .O(n13813) );
  NAND_GATE U14102 ( .I1(n13802), .I2(n13801), .O(n13807) );
  NAND_GATE U14103 ( .I1(n13803), .I2(n13807), .O(n13811) );
  NAND_GATE U14104 ( .I1(n13805), .I2(n13804), .O(n13806) );
  NAND_GATE U14105 ( .I1(n13807), .I2(n13806), .O(n13808) );
  NAND_GATE U14106 ( .I1(n13809), .I2(n13808), .O(n13810) );
  NAND_GATE U14107 ( .I1(n13811), .I2(n13810), .O(n13812) );
  NAND_GATE U14108 ( .I1(n13813), .I2(n13812), .O(n14229) );
  OR_GATE U14109 ( .I1(n13814), .I2(n13818), .O(n13817) );
  OR_GATE U14110 ( .I1(n13815), .I2(n13819), .O(n13816) );
  AND_GATE U14111 ( .I1(n13817), .I2(n13816), .O(n13824) );
  NAND_GATE U14112 ( .I1(n13818), .I2(n1189), .O(n13822) );
  NAND3_GATE U14113 ( .I1(n13822), .I2(n13821), .I3(n13820), .O(n13823) );
  NAND_GATE U14114 ( .I1(n13824), .I2(n13823), .O(n14238) );
  INV_GATE U14115 ( .I1(n14238), .O(n14241) );
  INV_GATE U14116 ( .I1(n13825), .O(n13826) );
  NAND_GATE U14117 ( .I1(n13830), .I2(n13826), .O(n13838) );
  NAND_GATE U14118 ( .I1(n13828), .I2(n13832), .O(n13836) );
  NAND_GATE U14119 ( .I1(n13830), .I2(n13829), .O(n13831) );
  NAND_GATE U14120 ( .I1(n13832), .I2(n13831), .O(n13833) );
  NAND_GATE U14121 ( .I1(n13834), .I2(n13833), .O(n13835) );
  NAND_GATE U14122 ( .I1(n13836), .I2(n13835), .O(n13837) );
  NAND_GATE U14123 ( .I1(n13838), .I2(n13837), .O(n14254) );
  NAND_GATE U14124 ( .I1(n1367), .I2(A[0]), .O(n13839) );
  NAND_GATE U14125 ( .I1(n14781), .I2(n13839), .O(n13840) );
  NAND_GATE U14126 ( .I1(B[4]), .I2(n13840), .O(n13844) );
  NAND_GATE U14127 ( .I1(n1368), .I2(A[1]), .O(n13841) );
  NAND_GATE U14128 ( .I1(n14784), .I2(n13841), .O(n13842) );
  NAND_GATE U14129 ( .I1(B[3]), .I2(n13842), .O(n13843) );
  NAND_GATE U14130 ( .I1(n13844), .I2(n13843), .O(n14266) );
  NAND_GATE U14131 ( .I1(n1365), .I2(A[2]), .O(n14270) );
  NAND3_GATE U14132 ( .I1(n1365), .I2(B[3]), .I3(n1196), .O(n14263) );
  NAND_GATE U14133 ( .I1(n14270), .I2(n14263), .O(n13845) );
  NAND_GATE U14134 ( .I1(n14266), .I2(n13845), .O(n13846) );
  INV_GATE U14135 ( .I1(n14270), .O(n14264) );
  INV_GATE U14136 ( .I1(n14263), .O(n14265) );
  NAND_GATE U14137 ( .I1(n14264), .I2(n14265), .O(n14261) );
  NAND_GATE U14138 ( .I1(n13846), .I2(n14261), .O(n14255) );
  NAND_GATE U14139 ( .I1(n14254), .I2(n14255), .O(n13848) );
  NAND_GATE U14140 ( .I1(n1365), .I2(A[3]), .O(n14256) );
  INV_GATE U14141 ( .I1(n14256), .O(n13847) );
  NAND_GATE U14142 ( .I1(n14254), .I2(n13847), .O(n14251) );
  NAND_GATE U14143 ( .I1(n14255), .I2(n13847), .O(n14250) );
  NAND3_GATE U14144 ( .I1(n13848), .I2(n14251), .I3(n14250), .O(n14240) );
  INV_GATE U14145 ( .I1(n14240), .O(n14237) );
  NAND_GATE U14146 ( .I1(n1365), .I2(A[4]), .O(n14245) );
  NAND_GATE U14147 ( .I1(n14237), .I2(n14245), .O(n13849) );
  NAND_GATE U14148 ( .I1(n14241), .I2(n13849), .O(n13850) );
  INV_GATE U14149 ( .I1(n14245), .O(n14239) );
  NAND_GATE U14150 ( .I1(n14240), .I2(n14239), .O(n14236) );
  NAND_GATE U14151 ( .I1(n13850), .I2(n14236), .O(n14230) );
  NAND_GATE U14152 ( .I1(n14229), .I2(n14230), .O(n13852) );
  NAND_GATE U14153 ( .I1(n1365), .I2(A[5]), .O(n14231) );
  INV_GATE U14154 ( .I1(n14231), .O(n13851) );
  NAND_GATE U14155 ( .I1(n14229), .I2(n13851), .O(n14226) );
  NAND_GATE U14156 ( .I1(n14230), .I2(n13851), .O(n14225) );
  NAND3_GATE U14157 ( .I1(n13852), .I2(n14226), .I3(n14225), .O(n14215) );
  INV_GATE U14158 ( .I1(n14215), .O(n14212) );
  NAND_GATE U14159 ( .I1(n1365), .I2(A[6]), .O(n14220) );
  NAND_GATE U14160 ( .I1(n14212), .I2(n14220), .O(n13853) );
  NAND_GATE U14161 ( .I1(n14216), .I2(n13853), .O(n13854) );
  INV_GATE U14162 ( .I1(n14220), .O(n14214) );
  NAND_GATE U14163 ( .I1(n14215), .I2(n14214), .O(n14211) );
  NAND_GATE U14164 ( .I1(n13854), .I2(n14211), .O(n14205) );
  NAND_GATE U14165 ( .I1(n14204), .I2(n14205), .O(n13856) );
  NAND_GATE U14166 ( .I1(n1365), .I2(A[7]), .O(n14206) );
  INV_GATE U14167 ( .I1(n14206), .O(n13855) );
  NAND_GATE U14168 ( .I1(n14204), .I2(n13855), .O(n14201) );
  NAND_GATE U14169 ( .I1(n14205), .I2(n13855), .O(n14200) );
  NAND3_GATE U14170 ( .I1(n13856), .I2(n14201), .I3(n14200), .O(n14190) );
  INV_GATE U14171 ( .I1(n14190), .O(n14187) );
  NAND_GATE U14172 ( .I1(n1365), .I2(A[8]), .O(n14195) );
  NAND_GATE U14173 ( .I1(n14187), .I2(n14195), .O(n13857) );
  NAND_GATE U14174 ( .I1(n14191), .I2(n13857), .O(n13858) );
  INV_GATE U14175 ( .I1(n14195), .O(n14189) );
  NAND_GATE U14176 ( .I1(n14190), .I2(n14189), .O(n14186) );
  NAND_GATE U14177 ( .I1(n13858), .I2(n14186), .O(n14180) );
  NAND_GATE U14178 ( .I1(n14179), .I2(n14180), .O(n13860) );
  NAND_GATE U14179 ( .I1(n1365), .I2(A[9]), .O(n14181) );
  INV_GATE U14180 ( .I1(n14181), .O(n13859) );
  NAND_GATE U14181 ( .I1(n14179), .I2(n13859), .O(n14176) );
  NAND_GATE U14182 ( .I1(n14180), .I2(n13859), .O(n14175) );
  NAND3_GATE U14183 ( .I1(n13860), .I2(n14176), .I3(n14175), .O(n14165) );
  INV_GATE U14184 ( .I1(n14165), .O(n14162) );
  NAND_GATE U14185 ( .I1(n1365), .I2(A[10]), .O(n14170) );
  NAND_GATE U14186 ( .I1(n14162), .I2(n14170), .O(n13861) );
  NAND_GATE U14187 ( .I1(n14166), .I2(n13861), .O(n13862) );
  INV_GATE U14188 ( .I1(n14170), .O(n14164) );
  NAND_GATE U14189 ( .I1(n14165), .I2(n14164), .O(n14161) );
  NAND_GATE U14190 ( .I1(n13862), .I2(n14161), .O(n14306) );
  NAND_GATE U14191 ( .I1(n14305), .I2(n14306), .O(n13864) );
  NAND_GATE U14192 ( .I1(n1365), .I2(A[11]), .O(n14307) );
  INV_GATE U14193 ( .I1(n14307), .O(n13863) );
  NAND_GATE U14194 ( .I1(n14306), .I2(n13863), .O(n14302) );
  NAND_GATE U14195 ( .I1(n14305), .I2(n13863), .O(n14301) );
  NAND3_GATE U14196 ( .I1(n13864), .I2(n14302), .I3(n14301), .O(n14152) );
  NAND_GATE U14197 ( .I1(n1365), .I2(A[12]), .O(n14156) );
  OR_GATE U14198 ( .I1(n13865), .I2(n13870), .O(n13868) );
  OR_GATE U14199 ( .I1(n13866), .I2(n13869), .O(n13867) );
  AND_GATE U14200 ( .I1(n13868), .I2(n13867), .O(n13875) );
  NAND_GATE U14201 ( .I1(n13869), .I2(n1016), .O(n13873) );
  NAND3_GATE U14202 ( .I1(n13873), .I2(n13872), .I3(n13871), .O(n13874) );
  NAND_GATE U14203 ( .I1(n13875), .I2(n13874), .O(n14148) );
  NAND_GATE U14204 ( .I1(n14156), .I2(n14148), .O(n13876) );
  NAND_GATE U14205 ( .I1(n14152), .I2(n13876), .O(n13877) );
  INV_GATE U14206 ( .I1(n14156), .O(n14150) );
  INV_GATE U14207 ( .I1(n14148), .O(n14151) );
  NAND_GATE U14208 ( .I1(n14150), .I2(n14151), .O(n14146) );
  NAND_GATE U14209 ( .I1(n13877), .I2(n14146), .O(n14321) );
  NAND_GATE U14210 ( .I1(n14320), .I2(n14321), .O(n13879) );
  NAND_GATE U14211 ( .I1(n1365), .I2(A[13]), .O(n14322) );
  INV_GATE U14212 ( .I1(n14322), .O(n13878) );
  NAND_GATE U14213 ( .I1(n14321), .I2(n13878), .O(n14317) );
  NAND_GATE U14214 ( .I1(n14320), .I2(n13878), .O(n14316) );
  NAND3_GATE U14215 ( .I1(n13879), .I2(n14317), .I3(n14316), .O(n14137) );
  NAND_GATE U14216 ( .I1(n1365), .I2(A[14]), .O(n14141) );
  OR_GATE U14217 ( .I1(n13880), .I2(n13885), .O(n13883) );
  OR_GATE U14218 ( .I1(n13881), .I2(n13884), .O(n13882) );
  NAND_GATE U14219 ( .I1(n13884), .I2(n1006), .O(n13888) );
  NAND3_GATE U14220 ( .I1(n13888), .I2(n13887), .I3(n13886), .O(n13889) );
  NAND_GATE U14221 ( .I1(n14141), .I2(n14133), .O(n13890) );
  NAND_GATE U14222 ( .I1(n14137), .I2(n13890), .O(n13891) );
  INV_GATE U14223 ( .I1(n14141), .O(n14135) );
  INV_GATE U14224 ( .I1(n14133), .O(n14136) );
  NAND_GATE U14225 ( .I1(n14135), .I2(n14136), .O(n14131) );
  NAND_GATE U14226 ( .I1(n13891), .I2(n14131), .O(n14336) );
  NAND_GATE U14227 ( .I1(n14335), .I2(n14336), .O(n13893) );
  NAND_GATE U14228 ( .I1(n1365), .I2(A[15]), .O(n14337) );
  INV_GATE U14229 ( .I1(n14337), .O(n13892) );
  NAND_GATE U14230 ( .I1(n14336), .I2(n13892), .O(n14332) );
  NAND_GATE U14231 ( .I1(n14335), .I2(n13892), .O(n14331) );
  NAND3_GATE U14232 ( .I1(n13893), .I2(n14332), .I3(n14331), .O(n14122) );
  NAND_GATE U14233 ( .I1(n1365), .I2(A[16]), .O(n14126) );
  OR_GATE U14234 ( .I1(n13894), .I2(n13899), .O(n13897) );
  OR_GATE U14235 ( .I1(n13895), .I2(n13898), .O(n13896) );
  NAND_GATE U14236 ( .I1(n13898), .I2(n993), .O(n13902) );
  NAND3_GATE U14237 ( .I1(n13902), .I2(n13901), .I3(n13900), .O(n13903) );
  NAND_GATE U14238 ( .I1(n14126), .I2(n14118), .O(n13904) );
  NAND_GATE U14239 ( .I1(n14122), .I2(n13904), .O(n13905) );
  INV_GATE U14240 ( .I1(n14126), .O(n14120) );
  INV_GATE U14241 ( .I1(n14118), .O(n14121) );
  NAND_GATE U14242 ( .I1(n14120), .I2(n14121), .O(n14116) );
  NAND_GATE U14243 ( .I1(n13905), .I2(n14116), .O(n14350) );
  NAND_GATE U14244 ( .I1(n14349), .I2(n14350), .O(n13907) );
  NAND_GATE U14245 ( .I1(n1365), .I2(A[17]), .O(n14351) );
  INV_GATE U14246 ( .I1(n14351), .O(n13906) );
  NAND_GATE U14247 ( .I1(n14350), .I2(n13906), .O(n14346) );
  NAND_GATE U14248 ( .I1(n14349), .I2(n13906), .O(n14345) );
  NAND3_GATE U14249 ( .I1(n13907), .I2(n14346), .I3(n14345), .O(n14107) );
  NAND_GATE U14250 ( .I1(n1365), .I2(A[18]), .O(n14111) );
  OR_GATE U14251 ( .I1(n13909), .I2(n13912), .O(n13910) );
  AND_GATE U14252 ( .I1(n13911), .I2(n13910), .O(n13918) );
  NAND_GATE U14253 ( .I1(n13912), .I2(n930), .O(n13916) );
  NAND3_GATE U14254 ( .I1(n13916), .I2(n13915), .I3(n13914), .O(n13917) );
  NAND_GATE U14255 ( .I1(n13918), .I2(n13917), .O(n14104) );
  NAND_GATE U14256 ( .I1(n14111), .I2(n14104), .O(n13919) );
  NAND_GATE U14257 ( .I1(n14107), .I2(n13919), .O(n13920) );
  INV_GATE U14258 ( .I1(n14111), .O(n14105) );
  INV_GATE U14259 ( .I1(n14104), .O(n14106) );
  NAND_GATE U14260 ( .I1(n14105), .I2(n14106), .O(n14102) );
  NAND_GATE U14261 ( .I1(n13920), .I2(n14102), .O(n14366) );
  NAND_GATE U14262 ( .I1(n14365), .I2(n14366), .O(n13922) );
  NAND_GATE U14263 ( .I1(n1365), .I2(A[19]), .O(n14367) );
  INV_GATE U14264 ( .I1(n14367), .O(n13921) );
  NAND_GATE U14265 ( .I1(n14366), .I2(n13921), .O(n14361) );
  NAND_GATE U14266 ( .I1(n14365), .I2(n13921), .O(n14360) );
  NAND3_GATE U14267 ( .I1(n13922), .I2(n14361), .I3(n14360), .O(n14093) );
  NAND_GATE U14268 ( .I1(n1365), .I2(A[20]), .O(n14097) );
  OR_GATE U14269 ( .I1(n13923), .I2(n13928), .O(n13926) );
  OR_GATE U14270 ( .I1(n13924), .I2(n13927), .O(n13925) );
  AND_GATE U14271 ( .I1(n13926), .I2(n13925), .O(n13933) );
  NAND_GATE U14272 ( .I1(n13927), .I2(n49), .O(n13931) );
  NAND3_GATE U14273 ( .I1(n13931), .I2(n13930), .I3(n13929), .O(n13932) );
  NAND_GATE U14274 ( .I1(n13933), .I2(n13932), .O(n14090) );
  NAND_GATE U14275 ( .I1(n14097), .I2(n14090), .O(n13934) );
  NAND_GATE U14276 ( .I1(n14093), .I2(n13934), .O(n13935) );
  INV_GATE U14277 ( .I1(n14097), .O(n14091) );
  INV_GATE U14278 ( .I1(n14090), .O(n14092) );
  NAND_GATE U14279 ( .I1(n14091), .I2(n14092), .O(n14088) );
  NAND_GATE U14280 ( .I1(n13935), .I2(n14088), .O(n14380) );
  NAND_GATE U14281 ( .I1(n1365), .I2(A[21]), .O(n14381) );
  INV_GATE U14282 ( .I1(n14381), .O(n13936) );
  NAND_GATE U14283 ( .I1(n14380), .I2(n13936), .O(n14376) );
  NAND_GATE U14284 ( .I1(n1365), .I2(A[22]), .O(n14083) );
  OR_GATE U14285 ( .I1(n13937), .I2(n13942), .O(n13940) );
  OR_GATE U14286 ( .I1(n13938), .I2(n13941), .O(n13939) );
  NAND_GATE U14287 ( .I1(n13941), .I2(n361), .O(n13945) );
  NAND3_GATE U14288 ( .I1(n13945), .I2(n13944), .I3(n13943), .O(n13946) );
  NAND_GATE U14289 ( .I1(n14083), .I2(n14080), .O(n13947) );
  NAND_GATE U14290 ( .I1(n14081), .I2(n13947), .O(n13948) );
  NAND_GATE U14291 ( .I1(n13948), .I2(n14078), .O(n14395) );
  NAND_GATE U14292 ( .I1(n14394), .I2(n14395), .O(n13950) );
  NAND_GATE U14293 ( .I1(n1365), .I2(A[23]), .O(n14396) );
  INV_GATE U14294 ( .I1(n14396), .O(n13949) );
  NAND_GATE U14295 ( .I1(n14394), .I2(n13949), .O(n14390) );
  NAND3_GATE U14296 ( .I1(n13950), .I2(n14391), .I3(n14390), .O(n14069) );
  NAND_GATE U14297 ( .I1(n1365), .I2(A[24]), .O(n14073) );
  OR_GATE U14298 ( .I1(n13951), .I2(n13956), .O(n13954) );
  OR_GATE U14299 ( .I1(n13952), .I2(n13955), .O(n13953) );
  NAND_GATE U14300 ( .I1(n13955), .I2(n365), .O(n13959) );
  NAND3_GATE U14301 ( .I1(n13959), .I2(n13958), .I3(n13957), .O(n13960) );
  NAND_GATE U14302 ( .I1(n14073), .I2(n14066), .O(n13961) );
  NAND_GATE U14303 ( .I1(n14069), .I2(n13961), .O(n13962) );
  INV_GATE U14304 ( .I1(n14073), .O(n14065) );
  INV_GATE U14305 ( .I1(n14066), .O(n14068) );
  NAND_GATE U14306 ( .I1(n14065), .I2(n14068), .O(n14063) );
  NAND_GATE U14307 ( .I1(n13962), .I2(n14063), .O(n14053) );
  NAND_GATE U14308 ( .I1(n14057), .I2(n14053), .O(n13964) );
  NAND_GATE U14309 ( .I1(n1365), .I2(A[25]), .O(n14054) );
  INV_GATE U14310 ( .I1(n14054), .O(n13963) );
  NAND_GATE U14311 ( .I1(n14053), .I2(n13963), .O(n14058) );
  NAND_GATE U14312 ( .I1(n14057), .I2(n13963), .O(n14061) );
  NAND3_GATE U14313 ( .I1(n13966), .I2(n13965), .I3(n652), .O(n13973) );
  NAND3_GATE U14314 ( .I1(n13969), .I2(n13968), .I3(n13967), .O(n13971) );
  NAND3_GATE U14315 ( .I1(n13972), .I2(n13971), .I3(n13970), .O(n14413) );
  INV_GATE U14316 ( .I1(n14413), .O(n14411) );
  NAND_GATE U14317 ( .I1(n13973), .I2(n14409), .O(n14046) );
  NAND_GATE U14318 ( .I1(n1365), .I2(A[27]), .O(n14043) );
  INV_GATE U14319 ( .I1(n14043), .O(n13987) );
  NAND_GATE U14320 ( .I1(n14046), .I2(n13987), .O(n14049) );
  NAND3_GATE U14321 ( .I1(n13979), .I2(n13978), .I3(n13975), .O(n13984) );
  NAND_GATE U14322 ( .I1(n13977), .I2(n13976), .O(n13983) );
  NAND_GATE U14323 ( .I1(n13979), .I2(n13978), .O(n13980) );
  NAND_GATE U14324 ( .I1(n13981), .I2(n13980), .O(n13982) );
  NAND3_GATE U14325 ( .I1(n13984), .I2(n13983), .I3(n13982), .O(n13985) );
  NAND_GATE U14326 ( .I1(n13986), .I2(n13985), .O(n14048) );
  NAND_GATE U14327 ( .I1(n14048), .I2(n13987), .O(n14047) );
  NAND_GATE U14328 ( .I1(n14046), .I2(n14048), .O(n13988) );
  NAND3_GATE U14329 ( .I1(n14049), .I2(n14047), .I3(n13988), .O(n14427) );
  NAND_GATE U14330 ( .I1(n14430), .I2(n14428), .O(n13989) );
  NAND_GATE U14331 ( .I1(n14427), .I2(n13989), .O(n13990) );
  NAND_GATE U14332 ( .I1(n14424), .I2(n13990), .O(n14033) );
  NAND3_GATE U14333 ( .I1(n13992), .I2(n506), .I3(n13991), .O(n13993) );
  NAND3_GATE U14334 ( .I1(n13995), .I2(n13994), .I3(n13993), .O(n14000) );
  INV_GATE U14335 ( .I1(n13996), .O(n13998) );
  NAND_GATE U14336 ( .I1(n13998), .I2(n13997), .O(n13999) );
  NAND_GATE U14337 ( .I1(n14000), .I2(n13999), .O(n14034) );
  NAND_GATE U14338 ( .I1(n14033), .I2(n14034), .O(n14002) );
  NAND_GATE U14339 ( .I1(n1365), .I2(A[29]), .O(n14042) );
  INV_GATE U14340 ( .I1(n14042), .O(n14001) );
  NAND_GATE U14341 ( .I1(n14001), .I2(n14034), .O(n14032) );
  NAND3_GATE U14342 ( .I1(n14002), .I2(n14032), .I3(n14035), .O(n14028) );
  NAND_GATE U14343 ( .I1(n14004), .I2(n14003), .O(n14022) );
  NAND_GATE U14344 ( .I1(n14021), .I2(n14022), .O(n14005) );
  NAND_GATE U14345 ( .I1(n14028), .I2(n14005), .O(n14006) );
  NAND_GATE U14346 ( .I1(n14027), .I2(n14006), .O(n14448) );
  NAND_GATE U14347 ( .I1(n14448), .I2(n14449), .O(n14008) );
  NAND_GATE U14348 ( .I1(n14445), .I2(n14448), .O(n14007) );
  NAND3_GATE U14349 ( .I1(n14009), .I2(n14008), .I3(n14007), .O(n15364) );
  NAND3_GATE U14350 ( .I1(n14010), .I2(n14011), .I3(n14012), .O(n14015) );
  NAND3_GATE U14351 ( .I1(n14015), .I2(n14014), .I3(n14013), .O(n14018) );
  NAND_GATE U14352 ( .I1(n1267), .I2(n14016), .O(n14017) );
  NAND_GATE U14353 ( .I1(n14018), .I2(n14017), .O(n15363) );
  NAND_GATE U14354 ( .I1(n15364), .I2(n665), .O(n14019) );
  NAND_GATE U14355 ( .I1(n14020), .I2(n14019), .O(\A1[32] ) );
  NAND3_GATE U14356 ( .I1(n14022), .I2(n568), .I3(n14021), .O(n14025) );
  NAND_GATE U14357 ( .I1(n14023), .I2(n14028), .O(n14024) );
  NAND4_GATE U14358 ( .I1(n14026), .I2(n14025), .I3(n14027), .I4(n14024), .O(
        n14031) );
  INV_GATE U14359 ( .I1(n14027), .O(n14029) );
  NAND_GATE U14360 ( .I1(n14029), .I2(n14028), .O(n14030) );
  NAND_GATE U14361 ( .I1(n14031), .I2(n14030), .O(n14457) );
  NAND_GATE U14362 ( .I1(n14033), .I2(n604), .O(n14041) );
  NAND3_GATE U14363 ( .I1(n14042), .I2(n14041), .I3(n14040), .O(n14036) );
  NAND_GATE U14364 ( .I1(B[1]), .I2(A[30]), .O(n14473) );
  INV_GATE U14365 ( .I1(n14473), .O(n14468) );
  NAND_GATE U14366 ( .I1(n1249), .I2(n14468), .O(n14466) );
  NAND_GATE U14367 ( .I1(n14038), .I2(n14037), .O(n14039) );
  NAND_GATE U14368 ( .I1(n14473), .I2(n14039), .O(n14441) );
  NAND4_GATE U14369 ( .I1(n14042), .I2(n14041), .I3(n14040), .I4(n14473), .O(
        n14440) );
  NAND_GATE U14370 ( .I1(n14046), .I2(n599), .O(n14044) );
  NAND3_GATE U14371 ( .I1(n14045), .I2(n14044), .I3(n14043), .O(n14052) );
  OR_GATE U14372 ( .I1(n14047), .I2(n14046), .O(n14051) );
  OR_GATE U14373 ( .I1(n14049), .I2(n14048), .O(n14050) );
  NAND3_GATE U14374 ( .I1(n14052), .I2(n14051), .I3(n14050), .O(n14482) );
  INV_GATE U14375 ( .I1(n14482), .O(n14484) );
  NAND_GATE U14376 ( .I1(B[1]), .I2(A[28]), .O(n14487) );
  INV_GATE U14377 ( .I1(n14487), .O(n14481) );
  NAND_GATE U14378 ( .I1(n14484), .I2(n14481), .O(n14478) );
  NAND_GATE U14379 ( .I1(B[1]), .I2(A[26]), .O(n14858) );
  NAND_GATE U14380 ( .I1(n14057), .I2(n14062), .O(n14056) );
  NAND_GATE U14381 ( .I1(n1333), .I2(n14053), .O(n14055) );
  NAND3_GATE U14382 ( .I1(n14056), .I2(n14055), .I3(n14054), .O(n14060) );
  OR_GATE U14383 ( .I1(n14058), .I2(n14057), .O(n14059) );
  NAND_GATE U14384 ( .I1(n14060), .I2(n14059), .O(n14407) );
  NAND_GATE U14385 ( .I1(n14858), .I2(n14407), .O(n14406) );
  NAND_GATE U14386 ( .I1(n281), .I2(n14858), .O(n14405) );
  INV_GATE U14387 ( .I1(n14063), .O(n14064) );
  NAND_GATE U14388 ( .I1(n14069), .I2(n14064), .O(n14077) );
  NAND_GATE U14389 ( .I1(n14065), .I2(n14071), .O(n14075) );
  NAND_GATE U14390 ( .I1(n14067), .I2(n14066), .O(n14071) );
  NAND_GATE U14391 ( .I1(n14069), .I2(n14068), .O(n14070) );
  NAND_GATE U14392 ( .I1(n14071), .I2(n14070), .O(n14072) );
  NAND_GATE U14393 ( .I1(n14073), .I2(n14072), .O(n14074) );
  NAND_GATE U14394 ( .I1(n14075), .I2(n14074), .O(n14076) );
  NAND_GATE U14395 ( .I1(n14077), .I2(n14076), .O(n14497) );
  INV_GATE U14396 ( .I1(n14078), .O(n14079) );
  NAND_GATE U14397 ( .I1(n14081), .I2(n14079), .O(n14087) );
  NAND_GATE U14398 ( .I1(n684), .I2(n14082), .O(n14085) );
  NAND_GATE U14399 ( .I1(n14085), .I2(n14084), .O(n14086) );
  NAND_GATE U14400 ( .I1(n14087), .I2(n14086), .O(n14506) );
  INV_GATE U14401 ( .I1(n14088), .O(n14089) );
  NAND_GATE U14402 ( .I1(n14093), .I2(n14089), .O(n14101) );
  NAND_GATE U14403 ( .I1(n63), .I2(n14090), .O(n14095) );
  NAND_GATE U14404 ( .I1(n14091), .I2(n14095), .O(n14099) );
  NAND_GATE U14405 ( .I1(n14093), .I2(n14092), .O(n14094) );
  NAND_GATE U14406 ( .I1(n14095), .I2(n14094), .O(n14096) );
  NAND_GATE U14407 ( .I1(n14097), .I2(n14096), .O(n14098) );
  NAND_GATE U14408 ( .I1(n14099), .I2(n14098), .O(n14100) );
  NAND_GATE U14409 ( .I1(n14101), .I2(n14100), .O(n14532) );
  INV_GATE U14410 ( .I1(n14102), .O(n14103) );
  NAND_GATE U14411 ( .I1(n14107), .I2(n14103), .O(n14115) );
  NAND_GATE U14412 ( .I1(n14105), .I2(n14109), .O(n14113) );
  NAND_GATE U14413 ( .I1(n14107), .I2(n14106), .O(n14108) );
  NAND_GATE U14414 ( .I1(n14109), .I2(n14108), .O(n14110) );
  NAND_GATE U14415 ( .I1(n14111), .I2(n14110), .O(n14112) );
  NAND_GATE U14416 ( .I1(n14113), .I2(n14112), .O(n14114) );
  NAND_GATE U14417 ( .I1(n14115), .I2(n14114), .O(n14556) );
  INV_GATE U14418 ( .I1(n14116), .O(n14117) );
  NAND_GATE U14419 ( .I1(n14122), .I2(n14117), .O(n14130) );
  INV_GATE U14420 ( .I1(n14122), .O(n14119) );
  NAND_GATE U14421 ( .I1(n14119), .I2(n14118), .O(n14124) );
  NAND_GATE U14422 ( .I1(n14120), .I2(n14124), .O(n14128) );
  NAND_GATE U14423 ( .I1(n14122), .I2(n14121), .O(n14123) );
  NAND_GATE U14424 ( .I1(n14124), .I2(n14123), .O(n14125) );
  NAND_GATE U14425 ( .I1(n14126), .I2(n14125), .O(n14127) );
  NAND_GATE U14426 ( .I1(n14128), .I2(n14127), .O(n14129) );
  NAND_GATE U14427 ( .I1(n14130), .I2(n14129), .O(n14581) );
  INV_GATE U14428 ( .I1(n14131), .O(n14132) );
  NAND_GATE U14429 ( .I1(n14137), .I2(n14132), .O(n14145) );
  INV_GATE U14430 ( .I1(n14137), .O(n14134) );
  NAND_GATE U14431 ( .I1(n14134), .I2(n14133), .O(n14139) );
  NAND_GATE U14432 ( .I1(n14135), .I2(n14139), .O(n14143) );
  NAND_GATE U14433 ( .I1(n14137), .I2(n14136), .O(n14138) );
  NAND_GATE U14434 ( .I1(n14139), .I2(n14138), .O(n14140) );
  NAND_GATE U14435 ( .I1(n14141), .I2(n14140), .O(n14142) );
  NAND_GATE U14436 ( .I1(n14143), .I2(n14142), .O(n14144) );
  NAND_GATE U14437 ( .I1(n14145), .I2(n14144), .O(n14607) );
  INV_GATE U14438 ( .I1(n14146), .O(n14147) );
  NAND_GATE U14439 ( .I1(n14152), .I2(n14147), .O(n14160) );
  INV_GATE U14440 ( .I1(n14152), .O(n14149) );
  NAND_GATE U14441 ( .I1(n14149), .I2(n14148), .O(n14154) );
  NAND_GATE U14442 ( .I1(n14150), .I2(n14154), .O(n14158) );
  NAND_GATE U14443 ( .I1(n14152), .I2(n14151), .O(n14153) );
  NAND_GATE U14444 ( .I1(n14154), .I2(n14153), .O(n14155) );
  NAND_GATE U14445 ( .I1(n14156), .I2(n14155), .O(n14157) );
  NAND_GATE U14446 ( .I1(n14158), .I2(n14157), .O(n14159) );
  NAND_GATE U14447 ( .I1(n14160), .I2(n14159), .O(n14633) );
  OR_GATE U14448 ( .I1(n14161), .I2(n14163), .O(n14174) );
  NAND_GATE U14449 ( .I1(n14163), .I2(n14162), .O(n14168) );
  NAND_GATE U14450 ( .I1(n14164), .I2(n14168), .O(n14172) );
  NAND_GATE U14451 ( .I1(n14166), .I2(n14165), .O(n14167) );
  NAND_GATE U14452 ( .I1(n14168), .I2(n14167), .O(n14169) );
  NAND_GATE U14453 ( .I1(n14170), .I2(n14169), .O(n14171) );
  NAND_GATE U14454 ( .I1(n14172), .I2(n14171), .O(n14173) );
  NAND_GATE U14455 ( .I1(n14174), .I2(n14173), .O(n14659) );
  OR_GATE U14456 ( .I1(n14175), .I2(n14179), .O(n14178) );
  OR_GATE U14457 ( .I1(n14176), .I2(n14180), .O(n14177) );
  AND_GATE U14458 ( .I1(n14178), .I2(n14177), .O(n14185) );
  NAND_GATE U14459 ( .I1(n14179), .I2(n1027), .O(n14183) );
  NAND3_GATE U14460 ( .I1(n14183), .I2(n14182), .I3(n14181), .O(n14184) );
  NAND_GATE U14461 ( .I1(n14185), .I2(n14184), .O(n14668) );
  INV_GATE U14462 ( .I1(n14668), .O(n14671) );
  OR_GATE U14463 ( .I1(n14186), .I2(n14188), .O(n14199) );
  NAND_GATE U14464 ( .I1(n14188), .I2(n14187), .O(n14193) );
  NAND_GATE U14465 ( .I1(n14189), .I2(n14193), .O(n14197) );
  NAND_GATE U14466 ( .I1(n14191), .I2(n14190), .O(n14192) );
  NAND_GATE U14467 ( .I1(n14193), .I2(n14192), .O(n14194) );
  NAND_GATE U14468 ( .I1(n14195), .I2(n14194), .O(n14196) );
  NAND_GATE U14469 ( .I1(n14197), .I2(n14196), .O(n14198) );
  NAND_GATE U14470 ( .I1(n14199), .I2(n14198), .O(n14684) );
  OR_GATE U14471 ( .I1(n14200), .I2(n14204), .O(n14203) );
  OR_GATE U14472 ( .I1(n14201), .I2(n14205), .O(n14202) );
  AND_GATE U14473 ( .I1(n14203), .I2(n14202), .O(n14210) );
  NAND_GATE U14474 ( .I1(n14204), .I2(n1030), .O(n14208) );
  NAND3_GATE U14475 ( .I1(n14208), .I2(n14207), .I3(n14206), .O(n14209) );
  NAND_GATE U14476 ( .I1(n14210), .I2(n14209), .O(n14693) );
  INV_GATE U14477 ( .I1(n14693), .O(n14696) );
  OR_GATE U14478 ( .I1(n14211), .I2(n14213), .O(n14224) );
  NAND_GATE U14479 ( .I1(n14213), .I2(n14212), .O(n14218) );
  NAND_GATE U14480 ( .I1(n14214), .I2(n14218), .O(n14222) );
  NAND_GATE U14481 ( .I1(n14216), .I2(n14215), .O(n14217) );
  NAND_GATE U14482 ( .I1(n14218), .I2(n14217), .O(n14219) );
  NAND_GATE U14483 ( .I1(n14220), .I2(n14219), .O(n14221) );
  NAND_GATE U14484 ( .I1(n14222), .I2(n14221), .O(n14223) );
  NAND_GATE U14485 ( .I1(n14224), .I2(n14223), .O(n14709) );
  OR_GATE U14486 ( .I1(n14225), .I2(n14229), .O(n14228) );
  OR_GATE U14487 ( .I1(n14226), .I2(n14230), .O(n14227) );
  AND_GATE U14488 ( .I1(n14228), .I2(n14227), .O(n14235) );
  NAND_GATE U14489 ( .I1(n14229), .I2(n1121), .O(n14233) );
  NAND3_GATE U14490 ( .I1(n14233), .I2(n14232), .I3(n14231), .O(n14234) );
  NAND_GATE U14491 ( .I1(n14235), .I2(n14234), .O(n14718) );
  INV_GATE U14492 ( .I1(n14718), .O(n14721) );
  OR_GATE U14493 ( .I1(n14236), .I2(n14238), .O(n14249) );
  NAND_GATE U14494 ( .I1(n14238), .I2(n14237), .O(n14243) );
  NAND_GATE U14495 ( .I1(n14239), .I2(n14243), .O(n14247) );
  NAND_GATE U14496 ( .I1(n14241), .I2(n14240), .O(n14242) );
  NAND_GATE U14497 ( .I1(n14243), .I2(n14242), .O(n14244) );
  NAND_GATE U14498 ( .I1(n14245), .I2(n14244), .O(n14246) );
  NAND_GATE U14499 ( .I1(n14247), .I2(n14246), .O(n14248) );
  NAND_GATE U14500 ( .I1(n14249), .I2(n14248), .O(n14734) );
  OR_GATE U14501 ( .I1(n14250), .I2(n14254), .O(n14253) );
  OR_GATE U14502 ( .I1(n14251), .I2(n14255), .O(n14252) );
  AND_GATE U14503 ( .I1(n14253), .I2(n14252), .O(n14260) );
  NAND_GATE U14504 ( .I1(n14254), .I2(n1190), .O(n14258) );
  NAND3_GATE U14505 ( .I1(n14258), .I2(n14257), .I3(n14256), .O(n14259) );
  NAND_GATE U14506 ( .I1(n14260), .I2(n14259), .O(n14743) );
  INV_GATE U14507 ( .I1(n14743), .O(n14746) );
  INV_GATE U14508 ( .I1(n14261), .O(n14262) );
  NAND_GATE U14509 ( .I1(n14266), .I2(n14262), .O(n14274) );
  NAND_GATE U14510 ( .I1(n14264), .I2(n14268), .O(n14272) );
  NAND_GATE U14511 ( .I1(n14266), .I2(n14265), .O(n14267) );
  NAND_GATE U14512 ( .I1(n14268), .I2(n14267), .O(n14269) );
  NAND_GATE U14513 ( .I1(n14270), .I2(n14269), .O(n14271) );
  NAND_GATE U14514 ( .I1(n14272), .I2(n14271), .O(n14273) );
  NAND_GATE U14515 ( .I1(n14274), .I2(n14273), .O(n14759) );
  NAND_GATE U14516 ( .I1(n1366), .I2(A[0]), .O(n14275) );
  NAND_GATE U14517 ( .I1(n14781), .I2(n14275), .O(n14276) );
  NAND_GATE U14518 ( .I1(B[3]), .I2(n14276), .O(n14280) );
  NAND_GATE U14519 ( .I1(n1367), .I2(A[1]), .O(n14277) );
  NAND_GATE U14520 ( .I1(n14784), .I2(n14277), .O(n14278) );
  NAND_GATE U14521 ( .I1(n1365), .I2(n14278), .O(n14279) );
  NAND_GATE U14522 ( .I1(n14280), .I2(n14279), .O(n14771) );
  NAND_GATE U14523 ( .I1(B[1]), .I2(A[2]), .O(n14775) );
  NAND3_GATE U14524 ( .I1(B[1]), .I2(n1365), .I3(n1196), .O(n14768) );
  NAND_GATE U14525 ( .I1(n14775), .I2(n14768), .O(n14281) );
  NAND_GATE U14526 ( .I1(n14771), .I2(n14281), .O(n14282) );
  INV_GATE U14527 ( .I1(n14775), .O(n14769) );
  INV_GATE U14528 ( .I1(n14768), .O(n14770) );
  NAND_GATE U14529 ( .I1(n14769), .I2(n14770), .O(n14766) );
  NAND_GATE U14530 ( .I1(n14282), .I2(n14766), .O(n14760) );
  NAND_GATE U14531 ( .I1(n14759), .I2(n14760), .O(n14284) );
  NAND_GATE U14532 ( .I1(B[1]), .I2(A[3]), .O(n14761) );
  INV_GATE U14533 ( .I1(n14761), .O(n14283) );
  NAND_GATE U14534 ( .I1(n14759), .I2(n14283), .O(n14756) );
  NAND_GATE U14535 ( .I1(n14760), .I2(n14283), .O(n14755) );
  NAND3_GATE U14536 ( .I1(n14284), .I2(n14756), .I3(n14755), .O(n14745) );
  INV_GATE U14537 ( .I1(n14745), .O(n14742) );
  NAND_GATE U14538 ( .I1(B[1]), .I2(A[4]), .O(n14750) );
  NAND_GATE U14539 ( .I1(n14742), .I2(n14750), .O(n14285) );
  NAND_GATE U14540 ( .I1(n14746), .I2(n14285), .O(n14286) );
  INV_GATE U14541 ( .I1(n14750), .O(n14744) );
  NAND_GATE U14542 ( .I1(n14745), .I2(n14744), .O(n14741) );
  NAND_GATE U14543 ( .I1(n14286), .I2(n14741), .O(n14735) );
  NAND_GATE U14544 ( .I1(n14734), .I2(n14735), .O(n14288) );
  NAND_GATE U14545 ( .I1(B[1]), .I2(A[5]), .O(n14736) );
  INV_GATE U14546 ( .I1(n14736), .O(n14287) );
  NAND_GATE U14547 ( .I1(n14734), .I2(n14287), .O(n14731) );
  NAND_GATE U14548 ( .I1(n14735), .I2(n14287), .O(n14730) );
  NAND3_GATE U14549 ( .I1(n14288), .I2(n14731), .I3(n14730), .O(n14720) );
  INV_GATE U14550 ( .I1(n14720), .O(n14717) );
  NAND_GATE U14551 ( .I1(B[1]), .I2(A[6]), .O(n14725) );
  NAND_GATE U14552 ( .I1(n14717), .I2(n14725), .O(n14289) );
  NAND_GATE U14553 ( .I1(n14721), .I2(n14289), .O(n14290) );
  INV_GATE U14554 ( .I1(n14725), .O(n14719) );
  NAND_GATE U14555 ( .I1(n14720), .I2(n14719), .O(n14716) );
  NAND_GATE U14556 ( .I1(n14290), .I2(n14716), .O(n14710) );
  NAND_GATE U14557 ( .I1(n14709), .I2(n14710), .O(n14292) );
  NAND_GATE U14558 ( .I1(B[1]), .I2(A[7]), .O(n14711) );
  INV_GATE U14559 ( .I1(n14711), .O(n14291) );
  NAND_GATE U14560 ( .I1(n14709), .I2(n14291), .O(n14706) );
  NAND_GATE U14561 ( .I1(n14710), .I2(n14291), .O(n14705) );
  NAND3_GATE U14562 ( .I1(n14292), .I2(n14706), .I3(n14705), .O(n14695) );
  INV_GATE U14563 ( .I1(n14695), .O(n14692) );
  NAND_GATE U14564 ( .I1(B[1]), .I2(A[8]), .O(n14700) );
  NAND_GATE U14565 ( .I1(n14692), .I2(n14700), .O(n14293) );
  NAND_GATE U14566 ( .I1(n14696), .I2(n14293), .O(n14294) );
  INV_GATE U14567 ( .I1(n14700), .O(n14694) );
  NAND_GATE U14568 ( .I1(n14695), .I2(n14694), .O(n14691) );
  NAND_GATE U14569 ( .I1(n14294), .I2(n14691), .O(n14685) );
  NAND_GATE U14570 ( .I1(n14684), .I2(n14685), .O(n14296) );
  NAND_GATE U14571 ( .I1(B[1]), .I2(A[9]), .O(n14686) );
  INV_GATE U14572 ( .I1(n14686), .O(n14295) );
  NAND_GATE U14573 ( .I1(n14684), .I2(n14295), .O(n14681) );
  NAND_GATE U14574 ( .I1(n14685), .I2(n14295), .O(n14680) );
  NAND3_GATE U14575 ( .I1(n14296), .I2(n14681), .I3(n14680), .O(n14670) );
  INV_GATE U14576 ( .I1(n14670), .O(n14667) );
  NAND_GATE U14577 ( .I1(B[1]), .I2(A[10]), .O(n14675) );
  NAND_GATE U14578 ( .I1(n14667), .I2(n14675), .O(n14297) );
  NAND_GATE U14579 ( .I1(n14671), .I2(n14297), .O(n14298) );
  INV_GATE U14580 ( .I1(n14675), .O(n14669) );
  NAND_GATE U14581 ( .I1(n14670), .I2(n14669), .O(n14666) );
  NAND_GATE U14582 ( .I1(n14298), .I2(n14666), .O(n14660) );
  NAND_GATE U14583 ( .I1(n14659), .I2(n14660), .O(n14300) );
  NAND_GATE U14584 ( .I1(B[1]), .I2(A[11]), .O(n14661) );
  INV_GATE U14585 ( .I1(n14661), .O(n14299) );
  NAND_GATE U14586 ( .I1(n14660), .I2(n14299), .O(n14656) );
  NAND_GATE U14587 ( .I1(n14659), .I2(n14299), .O(n14655) );
  NAND3_GATE U14588 ( .I1(n14300), .I2(n14656), .I3(n14655), .O(n14646) );
  NAND_GATE U14589 ( .I1(B[1]), .I2(A[12]), .O(n14650) );
  OR_GATE U14590 ( .I1(n14301), .I2(n14306), .O(n14304) );
  OR_GATE U14591 ( .I1(n14302), .I2(n14305), .O(n14303) );
  AND_GATE U14592 ( .I1(n14304), .I2(n14303), .O(n14311) );
  NAND_GATE U14593 ( .I1(n14305), .I2(n1020), .O(n14309) );
  NAND3_GATE U14594 ( .I1(n14309), .I2(n14308), .I3(n14307), .O(n14310) );
  NAND_GATE U14595 ( .I1(n14311), .I2(n14310), .O(n14642) );
  NAND_GATE U14596 ( .I1(n14650), .I2(n14642), .O(n14312) );
  NAND_GATE U14597 ( .I1(n14646), .I2(n14312), .O(n14313) );
  INV_GATE U14598 ( .I1(n14650), .O(n14644) );
  INV_GATE U14599 ( .I1(n14642), .O(n14645) );
  NAND_GATE U14600 ( .I1(n14644), .I2(n14645), .O(n14640) );
  NAND_GATE U14601 ( .I1(n14313), .I2(n14640), .O(n14634) );
  NAND_GATE U14602 ( .I1(n14633), .I2(n14634), .O(n14315) );
  NAND_GATE U14603 ( .I1(B[1]), .I2(A[13]), .O(n14635) );
  INV_GATE U14604 ( .I1(n14635), .O(n14314) );
  NAND_GATE U14605 ( .I1(n14634), .I2(n14314), .O(n14630) );
  NAND_GATE U14606 ( .I1(n14633), .I2(n14314), .O(n14629) );
  NAND3_GATE U14607 ( .I1(n14315), .I2(n14630), .I3(n14629), .O(n14620) );
  NAND_GATE U14608 ( .I1(B[1]), .I2(A[14]), .O(n14624) );
  OR_GATE U14609 ( .I1(n14316), .I2(n14321), .O(n14319) );
  OR_GATE U14610 ( .I1(n14317), .I2(n14320), .O(n14318) );
  AND_GATE U14611 ( .I1(n14319), .I2(n14318), .O(n14326) );
  NAND_GATE U14612 ( .I1(n14320), .I2(n1011), .O(n14324) );
  NAND3_GATE U14613 ( .I1(n14324), .I2(n14323), .I3(n14322), .O(n14325) );
  NAND_GATE U14614 ( .I1(n14326), .I2(n14325), .O(n14616) );
  NAND_GATE U14615 ( .I1(n14624), .I2(n14616), .O(n14327) );
  NAND_GATE U14616 ( .I1(n14620), .I2(n14327), .O(n14328) );
  INV_GATE U14617 ( .I1(n14624), .O(n14618) );
  INV_GATE U14618 ( .I1(n14616), .O(n14619) );
  NAND_GATE U14619 ( .I1(n14618), .I2(n14619), .O(n14614) );
  NAND_GATE U14620 ( .I1(n14328), .I2(n14614), .O(n14608) );
  NAND_GATE U14621 ( .I1(n14607), .I2(n14608), .O(n14330) );
  NAND_GATE U14622 ( .I1(B[1]), .I2(A[15]), .O(n14609) );
  INV_GATE U14623 ( .I1(n14609), .O(n14329) );
  NAND_GATE U14624 ( .I1(n14608), .I2(n14329), .O(n14604) );
  NAND_GATE U14625 ( .I1(n14607), .I2(n14329), .O(n14603) );
  NAND3_GATE U14626 ( .I1(n14330), .I2(n14604), .I3(n14603), .O(n14594) );
  NAND_GATE U14627 ( .I1(B[1]), .I2(A[16]), .O(n14598) );
  OR_GATE U14628 ( .I1(n14331), .I2(n14336), .O(n14334) );
  OR_GATE U14629 ( .I1(n14332), .I2(n14335), .O(n14333) );
  NAND_GATE U14630 ( .I1(n14335), .I2(n1001), .O(n14339) );
  NAND3_GATE U14631 ( .I1(n14339), .I2(n14338), .I3(n14337), .O(n14340) );
  NAND_GATE U14632 ( .I1(n14598), .I2(n14590), .O(n14341) );
  NAND_GATE U14633 ( .I1(n14594), .I2(n14341), .O(n14342) );
  INV_GATE U14634 ( .I1(n14598), .O(n14592) );
  INV_GATE U14635 ( .I1(n14590), .O(n14593) );
  NAND_GATE U14636 ( .I1(n14592), .I2(n14593), .O(n14588) );
  NAND_GATE U14637 ( .I1(n14342), .I2(n14588), .O(n14582) );
  NAND_GATE U14638 ( .I1(n14581), .I2(n14582), .O(n14344) );
  NAND_GATE U14639 ( .I1(B[1]), .I2(A[17]), .O(n14583) );
  INV_GATE U14640 ( .I1(n14583), .O(n14343) );
  NAND_GATE U14641 ( .I1(n14582), .I2(n14343), .O(n14578) );
  NAND_GATE U14642 ( .I1(n14581), .I2(n14343), .O(n14577) );
  NAND3_GATE U14643 ( .I1(n14344), .I2(n14578), .I3(n14577), .O(n14568) );
  NAND_GATE U14644 ( .I1(B[1]), .I2(A[18]), .O(n14572) );
  OR_GATE U14645 ( .I1(n14345), .I2(n14350), .O(n14348) );
  OR_GATE U14646 ( .I1(n14346), .I2(n14349), .O(n14347) );
  AND_GATE U14647 ( .I1(n14348), .I2(n14347), .O(n14355) );
  NAND_GATE U14648 ( .I1(n14349), .I2(n962), .O(n14353) );
  NAND3_GATE U14649 ( .I1(n14353), .I2(n14352), .I3(n14351), .O(n14354) );
  NAND_GATE U14650 ( .I1(n14355), .I2(n14354), .O(n14565) );
  NAND_GATE U14651 ( .I1(n14572), .I2(n14565), .O(n14356) );
  NAND_GATE U14652 ( .I1(n14568), .I2(n14356), .O(n14357) );
  INV_GATE U14653 ( .I1(n14572), .O(n14567) );
  NAND_GATE U14654 ( .I1(n14567), .I2(n644), .O(n14563) );
  NAND_GATE U14655 ( .I1(n14357), .I2(n14563), .O(n14557) );
  NAND_GATE U14656 ( .I1(n14556), .I2(n14557), .O(n14359) );
  NAND_GATE U14657 ( .I1(B[1]), .I2(A[19]), .O(n14558) );
  INV_GATE U14658 ( .I1(n14558), .O(n14358) );
  NAND_GATE U14659 ( .I1(n14557), .I2(n14358), .O(n14553) );
  NAND_GATE U14660 ( .I1(n14556), .I2(n14358), .O(n14552) );
  NAND3_GATE U14661 ( .I1(n14359), .I2(n14553), .I3(n14552), .O(n14543) );
  NAND_GATE U14662 ( .I1(B[1]), .I2(A[20]), .O(n14547) );
  OR_GATE U14663 ( .I1(n14361), .I2(n14365), .O(n14362) );
  AND_GATE U14664 ( .I1(n14363), .I2(n14362), .O(n14371) );
  INV_GATE U14665 ( .I1(n14366), .O(n14364) );
  NAND_GATE U14666 ( .I1(n14365), .I2(n14364), .O(n14369) );
  NAND_GATE U14667 ( .I1(n1283), .I2(n14366), .O(n14368) );
  NAND3_GATE U14668 ( .I1(n14369), .I2(n14368), .I3(n14367), .O(n14370) );
  NAND_GATE U14669 ( .I1(n14371), .I2(n14370), .O(n14540) );
  NAND_GATE U14670 ( .I1(n14547), .I2(n14540), .O(n14372) );
  NAND_GATE U14671 ( .I1(n14543), .I2(n14372), .O(n14373) );
  INV_GATE U14672 ( .I1(n14547), .O(n14541) );
  INV_GATE U14673 ( .I1(n14540), .O(n14542) );
  NAND_GATE U14674 ( .I1(n14541), .I2(n14542), .O(n14539) );
  NAND_GATE U14675 ( .I1(n14373), .I2(n14539), .O(n14533) );
  NAND_GATE U14676 ( .I1(n14532), .I2(n14533), .O(n14375) );
  NAND_GATE U14677 ( .I1(B[1]), .I2(A[21]), .O(n14534) );
  INV_GATE U14678 ( .I1(n14534), .O(n14374) );
  NAND_GATE U14679 ( .I1(n14533), .I2(n14374), .O(n14529) );
  NAND_GATE U14680 ( .I1(n14532), .I2(n14374), .O(n14528) );
  NAND3_GATE U14681 ( .I1(n14375), .I2(n14529), .I3(n14528), .O(n14519) );
  NAND_GATE U14682 ( .I1(B[1]), .I2(A[22]), .O(n14523) );
  OR_GATE U14683 ( .I1(n14376), .I2(n14379), .O(n14377) );
  AND_GATE U14684 ( .I1(n14378), .I2(n14377), .O(n14385) );
  NAND_GATE U14685 ( .I1(n14379), .I2(n556), .O(n14383) );
  NAND3_GATE U14686 ( .I1(n14383), .I2(n14382), .I3(n14381), .O(n14384) );
  NAND_GATE U14687 ( .I1(n14385), .I2(n14384), .O(n14515) );
  NAND_GATE U14688 ( .I1(n14523), .I2(n14515), .O(n14386) );
  NAND_GATE U14689 ( .I1(n14519), .I2(n14386), .O(n14387) );
  INV_GATE U14690 ( .I1(n14523), .O(n14517) );
  INV_GATE U14691 ( .I1(n14515), .O(n14518) );
  NAND_GATE U14692 ( .I1(n14517), .I2(n14518), .O(n14513) );
  NAND_GATE U14693 ( .I1(n14387), .I2(n14513), .O(n14507) );
  NAND_GATE U14694 ( .I1(n14506), .I2(n14507), .O(n14389) );
  NAND_GATE U14695 ( .I1(B[1]), .I2(A[23]), .O(n14508) );
  INV_GATE U14696 ( .I1(n14508), .O(n14388) );
  NAND_GATE U14697 ( .I1(n14507), .I2(n14388), .O(n14503) );
  NAND_GATE U14698 ( .I1(n14506), .I2(n14388), .O(n14502) );
  NAND3_GATE U14699 ( .I1(n14389), .I2(n14503), .I3(n14502), .O(n14840) );
  NAND_GATE U14700 ( .I1(B[1]), .I2(A[24]), .O(n14843) );
  OR_GATE U14701 ( .I1(n14391), .I2(n14394), .O(n14392) );
  AND_GATE U14702 ( .I1(n14393), .I2(n14392), .O(n14400) );
  NAND_GATE U14703 ( .I1(n14394), .I2(n418), .O(n14398) );
  NAND3_GATE U14704 ( .I1(n14398), .I2(n14397), .I3(n14396), .O(n14399) );
  NAND_GATE U14705 ( .I1(n14400), .I2(n14399), .O(n14838) );
  NAND_GATE U14706 ( .I1(n14843), .I2(n14838), .O(n14401) );
  NAND_GATE U14707 ( .I1(n14840), .I2(n14401), .O(n14402) );
  INV_GATE U14708 ( .I1(n14843), .O(n14837) );
  NAND_GATE U14709 ( .I1(n14837), .I2(n14839), .O(n14834) );
  NAND_GATE U14710 ( .I1(n14402), .I2(n14834), .O(n14495) );
  NAND_GATE U14711 ( .I1(B[1]), .I2(A[25]), .O(n14492) );
  INV_GATE U14712 ( .I1(n14492), .O(n14403) );
  NAND_GATE U14713 ( .I1(n14495), .I2(n14403), .O(n14498) );
  NAND3_GATE U14714 ( .I1(n14404), .I2(n14498), .I3(n14496), .O(n14856) );
  NAND3_GATE U14715 ( .I1(n14406), .I2(n14405), .I3(n14856), .O(n14408) );
  INV_GATE U14716 ( .I1(n14858), .O(n14854) );
  NAND_GATE U14717 ( .I1(n14854), .I2(n1357), .O(n14852) );
  NAND_GATE U14718 ( .I1(n14408), .I2(n14852), .O(n14867) );
  NAND_GATE U14719 ( .I1(B[1]), .I2(A[27]), .O(n14864) );
  INV_GATE U14720 ( .I1(n14864), .O(n14420) );
  NAND_GATE U14721 ( .I1(n14867), .I2(n14420), .O(n14870) );
  INV_GATE U14722 ( .I1(n14409), .O(n14410) );
  NAND_GATE U14723 ( .I1(n652), .I2(n14410), .O(n14419) );
  NAND_GATE U14724 ( .I1(n652), .I2(n14411), .O(n14417) );
  NAND3_GATE U14725 ( .I1(n14413), .I2(n862), .I3(n14412), .O(n14416) );
  NAND_GATE U14726 ( .I1(n862), .I2(n14413), .O(n14414) );
  NAND_GATE U14727 ( .I1(n466), .I2(n14414), .O(n14415) );
  NAND3_GATE U14728 ( .I1(n14417), .I2(n14416), .I3(n14415), .O(n14418) );
  NAND_GATE U14729 ( .I1(n14419), .I2(n14418), .O(n14869) );
  NAND_GATE U14730 ( .I1(n14869), .I2(n14420), .O(n14868) );
  NAND_GATE U14731 ( .I1(n14869), .I2(n14867), .O(n14421) );
  NAND3_GATE U14732 ( .I1(n14870), .I2(n14868), .I3(n14421), .O(n14483) );
  NAND_GATE U14733 ( .I1(n14482), .I2(n14487), .O(n14422) );
  NAND_GATE U14734 ( .I1(n14483), .I2(n14422), .O(n14423) );
  NAND_GATE U14735 ( .I1(n14478), .I2(n14423), .O(n14884) );
  NAND_GATE U14736 ( .I1(B[1]), .I2(A[29]), .O(n14886) );
  INV_GATE U14737 ( .I1(n14886), .O(n14438) );
  INV_GATE U14738 ( .I1(n14424), .O(n14425) );
  NAND_GATE U14739 ( .I1(n14425), .I2(n14427), .O(n14437) );
  NAND_GATE U14740 ( .I1(n14426), .I2(n14427), .O(n14435) );
  NAND3_GATE U14741 ( .I1(n14428), .I2(n14429), .I3(n14430), .O(n14434) );
  NAND_GATE U14742 ( .I1(n14430), .I2(n14429), .O(n14431) );
  NAND_GATE U14743 ( .I1(n14432), .I2(n14431), .O(n14433) );
  NAND3_GATE U14744 ( .I1(n14435), .I2(n14434), .I3(n14433), .O(n14436) );
  NAND_GATE U14745 ( .I1(n14437), .I2(n14436), .O(n14883) );
  NAND_GATE U14746 ( .I1(n14883), .I2(n14438), .O(n14878) );
  NAND_GATE U14747 ( .I1(n14883), .I2(n14884), .O(n14439) );
  NAND3_GATE U14748 ( .I1(n14879), .I2(n14878), .I3(n14439), .O(n14469) );
  NAND3_GATE U14749 ( .I1(n14441), .I2(n14440), .I3(n14469), .O(n14442) );
  NAND_GATE U14750 ( .I1(n14466), .I2(n14442), .O(n14462) );
  NAND_GATE U14751 ( .I1(n14457), .I2(n14462), .O(n14444) );
  NAND_GATE U14752 ( .I1(B[1]), .I2(A[31]), .O(n14458) );
  INV_GATE U14753 ( .I1(n14458), .O(n14443) );
  NAND_GATE U14754 ( .I1(n14443), .I2(n14462), .O(n14456) );
  NAND_GATE U14755 ( .I1(n14443), .I2(n14457), .O(n14461) );
  NAND3_GATE U14756 ( .I1(n14444), .I2(n14456), .I3(n14461), .O(n15365) );
  NAND3_GATE U14757 ( .I1(n14445), .I2(n592), .I3(n14449), .O(n14446) );
  NAND_GATE U14758 ( .I1(n592), .I2(n14449), .O(n14451) );
  NAND3_GATE U14759 ( .I1(n14452), .I2(n14451), .I3(n14450), .O(n14453) );
  NAND_GATE U14760 ( .I1(n15365), .I2(n1308), .O(n14454) );
  AND_GATE U14761 ( .I1(n14455), .I2(n14454), .O(\A1[31] ) );
  OR_GATE U14762 ( .I1(n14456), .I2(n14457), .O(n14465) );
  NAND_GATE U14763 ( .I1(n14457), .I2(n601), .O(n14460) );
  NAND3_GATE U14764 ( .I1(n14460), .I2(n14459), .I3(n14458), .O(n14464) );
  OR_GATE U14765 ( .I1(n14462), .I2(n14461), .O(n14463) );
  INV_GATE U14766 ( .I1(n14466), .O(n14467) );
  NAND_GATE U14767 ( .I1(n14467), .I2(n14469), .O(n14477) );
  NAND_GATE U14768 ( .I1(n14468), .I2(n14471), .O(n14475) );
  NAND_GATE U14769 ( .I1(n1249), .I2(n14469), .O(n14470) );
  NAND_GATE U14770 ( .I1(n14471), .I2(n14470), .O(n14472) );
  NAND_GATE U14771 ( .I1(n14473), .I2(n14472), .O(n14474) );
  NAND_GATE U14772 ( .I1(n14475), .I2(n14474), .O(n14476) );
  NAND_GATE U14773 ( .I1(n14477), .I2(n14476), .O(n14907) );
  NAND_GATE U14774 ( .I1(A[31]), .I2(B[0]), .O(n14902) );
  NAND_GATE U14775 ( .I1(A[30]), .I2(B[0]), .O(n14914) );
  INV_GATE U14776 ( .I1(n14478), .O(n14479) );
  NAND_GATE U14777 ( .I1(n14479), .I2(n14483), .O(n14491) );
  NAND_GATE U14778 ( .I1(n14482), .I2(n626), .O(n14480) );
  NAND_GATE U14779 ( .I1(n14481), .I2(n14480), .O(n14489) );
  NAND_GATE U14780 ( .I1(n14484), .I2(n14483), .O(n14485) );
  NAND_GATE U14781 ( .I1(n14480), .I2(n14485), .O(n14486) );
  NAND_GATE U14782 ( .I1(n14487), .I2(n14486), .O(n14488) );
  NAND_GATE U14783 ( .I1(n14489), .I2(n14488), .O(n14490) );
  NAND_GATE U14784 ( .I1(n14491), .I2(n14490), .O(n14929) );
  NAND_GATE U14785 ( .I1(A[29]), .I2(B[0]), .O(n14924) );
  NAND_GATE U14786 ( .I1(A[28]), .I2(B[0]), .O(n14937) );
  NAND_GATE U14787 ( .I1(A[27]), .I2(B[0]), .O(n14946) );
  INV_GATE U14788 ( .I1(n14946), .O(n14942) );
  NAND_GATE U14789 ( .I1(n14497), .I2(n435), .O(n14494) );
  NAND3_GATE U14790 ( .I1(n14494), .I2(n14493), .I3(n14492), .O(n14501) );
  OR_GATE U14791 ( .I1(n14496), .I2(n14495), .O(n14500) );
  OR_GATE U14792 ( .I1(n14498), .I2(n14497), .O(n14499) );
  NAND3_GATE U14793 ( .I1(n14501), .I2(n14500), .I3(n14499), .O(n14963) );
  NAND_GATE U14794 ( .I1(A[25]), .I2(B[0]), .O(n14972) );
  INV_GATE U14795 ( .I1(n14972), .O(n14968) );
  OR_GATE U14796 ( .I1(n14502), .I2(n14507), .O(n14505) );
  OR_GATE U14797 ( .I1(n14503), .I2(n14506), .O(n14504) );
  AND_GATE U14798 ( .I1(n14505), .I2(n14504), .O(n14512) );
  NAND_GATE U14799 ( .I1(n14506), .I2(n984), .O(n14510) );
  NAND3_GATE U14800 ( .I1(n14510), .I2(n14509), .I3(n14508), .O(n14511) );
  NAND_GATE U14801 ( .I1(n14512), .I2(n14511), .O(n14988) );
  INV_GATE U14802 ( .I1(n14988), .O(n14981) );
  INV_GATE U14803 ( .I1(n14513), .O(n14514) );
  NAND_GATE U14804 ( .I1(n14519), .I2(n14514), .O(n14527) );
  INV_GATE U14805 ( .I1(n14519), .O(n14516) );
  NAND_GATE U14806 ( .I1(n14516), .I2(n14515), .O(n14521) );
  NAND_GATE U14807 ( .I1(n14517), .I2(n14521), .O(n14525) );
  NAND_GATE U14808 ( .I1(n14519), .I2(n14518), .O(n14520) );
  NAND_GATE U14809 ( .I1(n14521), .I2(n14520), .O(n14522) );
  NAND_GATE U14810 ( .I1(n14523), .I2(n14522), .O(n14524) );
  NAND_GATE U14811 ( .I1(n14525), .I2(n14524), .O(n14526) );
  NAND_GATE U14812 ( .I1(n14527), .I2(n14526), .O(n15003) );
  OR_GATE U14813 ( .I1(n14528), .I2(n14533), .O(n14531) );
  OR_GATE U14814 ( .I1(n14529), .I2(n14532), .O(n14530) );
  AND_GATE U14815 ( .I1(n14531), .I2(n14530), .O(n14538) );
  NAND_GATE U14816 ( .I1(n14532), .I2(n966), .O(n14536) );
  NAND3_GATE U14817 ( .I1(n14536), .I2(n14535), .I3(n14534), .O(n14537) );
  NAND_GATE U14818 ( .I1(n14541), .I2(n14545), .O(n14549) );
  NAND_GATE U14819 ( .I1(n14543), .I2(n14542), .O(n14544) );
  NAND_GATE U14820 ( .I1(n14545), .I2(n14544), .O(n14546) );
  NAND_GATE U14821 ( .I1(n14547), .I2(n14546), .O(n14548) );
  NAND_GATE U14822 ( .I1(n14549), .I2(n14548), .O(n14550) );
  NAND_GATE U14823 ( .I1(n14551), .I2(n14550), .O(n15029) );
  OR_GATE U14824 ( .I1(n14552), .I2(n14557), .O(n14555) );
  OR_GATE U14825 ( .I1(n14553), .I2(n14556), .O(n14554) );
  AND_GATE U14826 ( .I1(n14555), .I2(n14554), .O(n14562) );
  NAND_GATE U14827 ( .I1(n14556), .I2(n934), .O(n14560) );
  NAND3_GATE U14828 ( .I1(n14560), .I2(n14559), .I3(n14558), .O(n14561) );
  NAND_GATE U14829 ( .I1(n14562), .I2(n14561), .O(n15041) );
  INV_GATE U14830 ( .I1(n15041), .O(n15034) );
  INV_GATE U14831 ( .I1(n14563), .O(n14564) );
  NAND_GATE U14832 ( .I1(n14568), .I2(n14564), .O(n14576) );
  INV_GATE U14833 ( .I1(n14568), .O(n14566) );
  NAND_GATE U14834 ( .I1(n14566), .I2(n14565), .O(n14570) );
  NAND_GATE U14835 ( .I1(n14567), .I2(n14570), .O(n14574) );
  NAND_GATE U14836 ( .I1(n14568), .I2(n644), .O(n14569) );
  NAND_GATE U14837 ( .I1(n14570), .I2(n14569), .O(n14571) );
  NAND_GATE U14838 ( .I1(n14572), .I2(n14571), .O(n14573) );
  NAND_GATE U14839 ( .I1(n14574), .I2(n14573), .O(n14575) );
  NAND_GATE U14840 ( .I1(n14576), .I2(n14575), .O(n15056) );
  OR_GATE U14841 ( .I1(n14577), .I2(n14582), .O(n14580) );
  OR_GATE U14842 ( .I1(n14578), .I2(n14581), .O(n14579) );
  AND_GATE U14843 ( .I1(n14580), .I2(n14579), .O(n14587) );
  NAND_GATE U14844 ( .I1(n14581), .I2(n995), .O(n14585) );
  NAND3_GATE U14845 ( .I1(n14585), .I2(n14584), .I3(n14583), .O(n14586) );
  NAND_GATE U14846 ( .I1(n14587), .I2(n14586), .O(n15069) );
  INV_GATE U14847 ( .I1(n15069), .O(n15062) );
  INV_GATE U14848 ( .I1(n14588), .O(n14589) );
  NAND_GATE U14849 ( .I1(n14594), .I2(n14589), .O(n14602) );
  INV_GATE U14850 ( .I1(n14594), .O(n14591) );
  NAND_GATE U14851 ( .I1(n14591), .I2(n14590), .O(n14596) );
  NAND_GATE U14852 ( .I1(n14592), .I2(n14596), .O(n14600) );
  NAND_GATE U14853 ( .I1(n14594), .I2(n14593), .O(n14595) );
  NAND_GATE U14854 ( .I1(n14596), .I2(n14595), .O(n14597) );
  NAND_GATE U14855 ( .I1(n14598), .I2(n14597), .O(n14599) );
  NAND_GATE U14856 ( .I1(n14600), .I2(n14599), .O(n14601) );
  NAND_GATE U14857 ( .I1(n14602), .I2(n14601), .O(n15085) );
  OR_GATE U14858 ( .I1(n14603), .I2(n14608), .O(n14606) );
  OR_GATE U14859 ( .I1(n14604), .I2(n14607), .O(n14605) );
  AND_GATE U14860 ( .I1(n14606), .I2(n14605), .O(n14613) );
  NAND_GATE U14861 ( .I1(n14607), .I2(n1008), .O(n14611) );
  NAND3_GATE U14862 ( .I1(n14611), .I2(n14610), .I3(n14609), .O(n14612) );
  NAND_GATE U14863 ( .I1(n14613), .I2(n14612), .O(n15098) );
  INV_GATE U14864 ( .I1(n15098), .O(n15091) );
  INV_GATE U14865 ( .I1(n14614), .O(n14615) );
  NAND_GATE U14866 ( .I1(n14620), .I2(n14615), .O(n14628) );
  INV_GATE U14867 ( .I1(n14620), .O(n14617) );
  NAND_GATE U14868 ( .I1(n14617), .I2(n14616), .O(n14622) );
  NAND_GATE U14869 ( .I1(n14618), .I2(n14622), .O(n14626) );
  NAND_GATE U14870 ( .I1(n14620), .I2(n14619), .O(n14621) );
  NAND_GATE U14871 ( .I1(n14622), .I2(n14621), .O(n14623) );
  NAND_GATE U14872 ( .I1(n14624), .I2(n14623), .O(n14625) );
  NAND_GATE U14873 ( .I1(n14626), .I2(n14625), .O(n14627) );
  NAND_GATE U14874 ( .I1(n14628), .I2(n14627), .O(n15114) );
  OR_GATE U14875 ( .I1(n14629), .I2(n14634), .O(n14632) );
  OR_GATE U14876 ( .I1(n14630), .I2(n14633), .O(n14631) );
  AND_GATE U14877 ( .I1(n14632), .I2(n14631), .O(n14639) );
  NAND_GATE U14878 ( .I1(n14633), .I2(n1017), .O(n14637) );
  NAND3_GATE U14879 ( .I1(n14637), .I2(n14636), .I3(n14635), .O(n14638) );
  NAND_GATE U14880 ( .I1(n14639), .I2(n14638), .O(n15127) );
  INV_GATE U14881 ( .I1(n15127), .O(n15120) );
  INV_GATE U14882 ( .I1(n14640), .O(n14641) );
  NAND_GATE U14883 ( .I1(n14646), .I2(n14641), .O(n14654) );
  INV_GATE U14884 ( .I1(n14646), .O(n14643) );
  NAND_GATE U14885 ( .I1(n14643), .I2(n14642), .O(n14648) );
  NAND_GATE U14886 ( .I1(n14644), .I2(n14648), .O(n14652) );
  NAND_GATE U14887 ( .I1(n14646), .I2(n14645), .O(n14647) );
  NAND_GATE U14888 ( .I1(n14648), .I2(n14647), .O(n14649) );
  NAND_GATE U14889 ( .I1(n14650), .I2(n14649), .O(n14651) );
  NAND_GATE U14890 ( .I1(n14652), .I2(n14651), .O(n14653) );
  NAND_GATE U14891 ( .I1(n14654), .I2(n14653), .O(n15143) );
  OR_GATE U14892 ( .I1(n14655), .I2(n14660), .O(n14658) );
  OR_GATE U14893 ( .I1(n14656), .I2(n14659), .O(n14657) );
  AND_GATE U14894 ( .I1(n14658), .I2(n14657), .O(n14665) );
  NAND_GATE U14895 ( .I1(n14659), .I2(n1025), .O(n14663) );
  NAND3_GATE U14896 ( .I1(n14663), .I2(n14662), .I3(n14661), .O(n14664) );
  NAND_GATE U14897 ( .I1(n14665), .I2(n14664), .O(n15156) );
  INV_GATE U14898 ( .I1(n15156), .O(n15149) );
  OR_GATE U14899 ( .I1(n14666), .I2(n14668), .O(n14679) );
  NAND_GATE U14900 ( .I1(n14668), .I2(n14667), .O(n14673) );
  NAND_GATE U14901 ( .I1(n14669), .I2(n14673), .O(n14677) );
  NAND_GATE U14902 ( .I1(n14671), .I2(n14670), .O(n14672) );
  NAND_GATE U14903 ( .I1(n14673), .I2(n14672), .O(n14674) );
  NAND_GATE U14904 ( .I1(n14675), .I2(n14674), .O(n14676) );
  NAND_GATE U14905 ( .I1(n14677), .I2(n14676), .O(n14678) );
  NAND_GATE U14906 ( .I1(n14679), .I2(n14678), .O(n15172) );
  OR_GATE U14907 ( .I1(n14680), .I2(n14684), .O(n14683) );
  OR_GATE U14908 ( .I1(n14681), .I2(n14685), .O(n14682) );
  AND_GATE U14909 ( .I1(n14683), .I2(n14682), .O(n14690) );
  NAND_GATE U14910 ( .I1(n14684), .I2(n1029), .O(n14688) );
  NAND3_GATE U14911 ( .I1(n14688), .I2(n14687), .I3(n14686), .O(n14689) );
  NAND_GATE U14912 ( .I1(n14690), .I2(n14689), .O(n15185) );
  INV_GATE U14913 ( .I1(n15185), .O(n15178) );
  OR_GATE U14914 ( .I1(n14691), .I2(n14693), .O(n14704) );
  NAND_GATE U14915 ( .I1(n14693), .I2(n14692), .O(n14698) );
  NAND_GATE U14916 ( .I1(n14694), .I2(n14698), .O(n14702) );
  NAND_GATE U14917 ( .I1(n14696), .I2(n14695), .O(n14697) );
  NAND_GATE U14918 ( .I1(n14698), .I2(n14697), .O(n14699) );
  NAND_GATE U14919 ( .I1(n14700), .I2(n14699), .O(n14701) );
  NAND_GATE U14920 ( .I1(n14702), .I2(n14701), .O(n14703) );
  NAND_GATE U14921 ( .I1(n14704), .I2(n14703), .O(n15201) );
  OR_GATE U14922 ( .I1(n14705), .I2(n14709), .O(n14708) );
  OR_GATE U14923 ( .I1(n14706), .I2(n14710), .O(n14707) );
  AND_GATE U14924 ( .I1(n14708), .I2(n14707), .O(n14715) );
  NAND_GATE U14925 ( .I1(n14709), .I2(n1031), .O(n14713) );
  NAND3_GATE U14926 ( .I1(n14713), .I2(n14712), .I3(n14711), .O(n14714) );
  NAND_GATE U14927 ( .I1(n14715), .I2(n14714), .O(n15214) );
  INV_GATE U14928 ( .I1(n15214), .O(n15207) );
  OR_GATE U14929 ( .I1(n14716), .I2(n14718), .O(n14729) );
  NAND_GATE U14930 ( .I1(n14718), .I2(n14717), .O(n14723) );
  NAND_GATE U14931 ( .I1(n14719), .I2(n14723), .O(n14727) );
  NAND_GATE U14932 ( .I1(n14721), .I2(n14720), .O(n14722) );
  NAND_GATE U14933 ( .I1(n14723), .I2(n14722), .O(n14724) );
  NAND_GATE U14934 ( .I1(n14725), .I2(n14724), .O(n14726) );
  NAND_GATE U14935 ( .I1(n14727), .I2(n14726), .O(n14728) );
  NAND_GATE U14936 ( .I1(n14729), .I2(n14728), .O(n15230) );
  OR_GATE U14937 ( .I1(n14730), .I2(n14734), .O(n14733) );
  OR_GATE U14938 ( .I1(n14731), .I2(n14735), .O(n14732) );
  AND_GATE U14939 ( .I1(n14733), .I2(n14732), .O(n14740) );
  NAND_GATE U14940 ( .I1(n14734), .I2(n1124), .O(n14738) );
  NAND3_GATE U14941 ( .I1(n14738), .I2(n14737), .I3(n14736), .O(n14739) );
  NAND_GATE U14942 ( .I1(n14740), .I2(n14739), .O(n15243) );
  INV_GATE U14943 ( .I1(n15243), .O(n15236) );
  OR_GATE U14944 ( .I1(n14741), .I2(n14743), .O(n14754) );
  NAND_GATE U14945 ( .I1(n14743), .I2(n14742), .O(n14748) );
  NAND_GATE U14946 ( .I1(n14744), .I2(n14748), .O(n14752) );
  NAND_GATE U14947 ( .I1(n14746), .I2(n14745), .O(n14747) );
  NAND_GATE U14948 ( .I1(n14748), .I2(n14747), .O(n14749) );
  NAND_GATE U14949 ( .I1(n14750), .I2(n14749), .O(n14751) );
  NAND_GATE U14950 ( .I1(n14752), .I2(n14751), .O(n14753) );
  NAND_GATE U14951 ( .I1(n14754), .I2(n14753), .O(n15259) );
  OR_GATE U14952 ( .I1(n14755), .I2(n14759), .O(n14758) );
  OR_GATE U14953 ( .I1(n14756), .I2(n14760), .O(n14757) );
  AND_GATE U14954 ( .I1(n14758), .I2(n14757), .O(n14765) );
  NAND_GATE U14955 ( .I1(n14759), .I2(n1191), .O(n14763) );
  NAND3_GATE U14956 ( .I1(n14763), .I2(n14762), .I3(n14761), .O(n14764) );
  NAND_GATE U14957 ( .I1(n14765), .I2(n14764), .O(n15272) );
  INV_GATE U14958 ( .I1(n15272), .O(n15265) );
  INV_GATE U14959 ( .I1(n14766), .O(n14767) );
  NAND_GATE U14960 ( .I1(n14771), .I2(n14767), .O(n14779) );
  NAND_GATE U14961 ( .I1(n14769), .I2(n14773), .O(n14777) );
  NAND_GATE U14962 ( .I1(n14771), .I2(n14770), .O(n14772) );
  NAND_GATE U14963 ( .I1(n14773), .I2(n14772), .O(n14774) );
  NAND_GATE U14964 ( .I1(n14775), .I2(n14774), .O(n14776) );
  NAND_GATE U14965 ( .I1(n14777), .I2(n14776), .O(n14778) );
  NAND_GATE U14966 ( .I1(n14779), .I2(n14778), .O(n15288) );
  NAND3_GATE U14967 ( .I1(B[1]), .I2(B[0]), .I3(n1196), .O(n15301) );
  INV_GATE U14968 ( .I1(n15301), .O(n15294) );
  NAND_GATE U14969 ( .I1(n1364), .I2(A[0]), .O(n14780) );
  NAND_GATE U14970 ( .I1(n14781), .I2(n14780), .O(n14782) );
  NAND_GATE U14971 ( .I1(n1365), .I2(n14782), .O(n14787) );
  NAND_GATE U14972 ( .I1(n1366), .I2(A[1]), .O(n14783) );
  NAND_GATE U14973 ( .I1(n14784), .I2(n14783), .O(n14785) );
  NAND_GATE U14974 ( .I1(B[1]), .I2(n14785), .O(n14786) );
  NAND_GATE U14975 ( .I1(n14787), .I2(n14786), .O(n15293) );
  INV_GATE U14976 ( .I1(n15293), .O(n15291) );
  NAND_GATE U14977 ( .I1(A[2]), .I2(B[0]), .O(n15298) );
  NAND_GATE U14978 ( .I1(n15291), .I2(n15298), .O(n14788) );
  NAND_GATE U14979 ( .I1(n15294), .I2(n14788), .O(n14789) );
  INV_GATE U14980 ( .I1(n15298), .O(n15292) );
  NAND_GATE U14981 ( .I1(n15293), .I2(n15292), .O(n15302) );
  NAND_GATE U14982 ( .I1(n14789), .I2(n15302), .O(n15278) );
  INV_GATE U14983 ( .I1(n15278), .O(n15280) );
  NAND_GATE U14984 ( .I1(A[3]), .I2(B[0]), .O(n15283) );
  NAND_GATE U14985 ( .I1(n15280), .I2(n15283), .O(n14790) );
  NAND_GATE U14986 ( .I1(n15288), .I2(n14790), .O(n14791) );
  INV_GATE U14987 ( .I1(n15283), .O(n15277) );
  NAND_GATE U14988 ( .I1(n15278), .I2(n15277), .O(n15286) );
  NAND_GATE U14989 ( .I1(n14791), .I2(n15286), .O(n15264) );
  INV_GATE U14990 ( .I1(n15264), .O(n15262) );
  NAND_GATE U14991 ( .I1(A[4]), .I2(B[0]), .O(n15269) );
  NAND_GATE U14992 ( .I1(n15262), .I2(n15269), .O(n14792) );
  NAND_GATE U14993 ( .I1(n15265), .I2(n14792), .O(n14793) );
  INV_GATE U14994 ( .I1(n15269), .O(n15263) );
  NAND_GATE U14995 ( .I1(n15264), .I2(n15263), .O(n15273) );
  NAND_GATE U14996 ( .I1(n14793), .I2(n15273), .O(n15249) );
  INV_GATE U14997 ( .I1(n15249), .O(n15251) );
  NAND_GATE U14998 ( .I1(A[5]), .I2(B[0]), .O(n15254) );
  NAND_GATE U14999 ( .I1(n15251), .I2(n15254), .O(n14794) );
  NAND_GATE U15000 ( .I1(n15259), .I2(n14794), .O(n14795) );
  INV_GATE U15001 ( .I1(n15254), .O(n15248) );
  NAND_GATE U15002 ( .I1(n15249), .I2(n15248), .O(n15257) );
  NAND_GATE U15003 ( .I1(n14795), .I2(n15257), .O(n15235) );
  INV_GATE U15004 ( .I1(n15235), .O(n15233) );
  NAND_GATE U15005 ( .I1(A[6]), .I2(B[0]), .O(n15240) );
  NAND_GATE U15006 ( .I1(n15233), .I2(n15240), .O(n14796) );
  NAND_GATE U15007 ( .I1(n15236), .I2(n14796), .O(n14797) );
  INV_GATE U15008 ( .I1(n15240), .O(n15234) );
  NAND_GATE U15009 ( .I1(n15235), .I2(n15234), .O(n15244) );
  NAND_GATE U15010 ( .I1(n14797), .I2(n15244), .O(n15220) );
  INV_GATE U15011 ( .I1(n15220), .O(n15222) );
  NAND_GATE U15012 ( .I1(A[7]), .I2(B[0]), .O(n15225) );
  NAND_GATE U15013 ( .I1(n15222), .I2(n15225), .O(n14798) );
  NAND_GATE U15014 ( .I1(n15230), .I2(n14798), .O(n14799) );
  INV_GATE U15015 ( .I1(n15225), .O(n15219) );
  NAND_GATE U15016 ( .I1(n15220), .I2(n15219), .O(n15228) );
  NAND_GATE U15017 ( .I1(n14799), .I2(n15228), .O(n15206) );
  INV_GATE U15018 ( .I1(n15206), .O(n15204) );
  NAND_GATE U15019 ( .I1(A[8]), .I2(B[0]), .O(n15211) );
  NAND_GATE U15020 ( .I1(n15204), .I2(n15211), .O(n14800) );
  NAND_GATE U15021 ( .I1(n15207), .I2(n14800), .O(n14801) );
  INV_GATE U15022 ( .I1(n15211), .O(n15205) );
  NAND_GATE U15023 ( .I1(n15206), .I2(n15205), .O(n15215) );
  NAND_GATE U15024 ( .I1(n14801), .I2(n15215), .O(n15191) );
  INV_GATE U15025 ( .I1(n15191), .O(n15193) );
  NAND_GATE U15026 ( .I1(A[9]), .I2(B[0]), .O(n15196) );
  NAND_GATE U15027 ( .I1(n15193), .I2(n15196), .O(n14802) );
  NAND_GATE U15028 ( .I1(n15201), .I2(n14802), .O(n14803) );
  INV_GATE U15029 ( .I1(n15196), .O(n15190) );
  NAND_GATE U15030 ( .I1(n15191), .I2(n15190), .O(n15199) );
  NAND_GATE U15031 ( .I1(n14803), .I2(n15199), .O(n15177) );
  INV_GATE U15032 ( .I1(n15177), .O(n15175) );
  NAND_GATE U15033 ( .I1(A[10]), .I2(B[0]), .O(n15182) );
  NAND_GATE U15034 ( .I1(n15175), .I2(n15182), .O(n14804) );
  NAND_GATE U15035 ( .I1(n15178), .I2(n14804), .O(n14805) );
  INV_GATE U15036 ( .I1(n15182), .O(n15176) );
  NAND_GATE U15037 ( .I1(n15177), .I2(n15176), .O(n15186) );
  NAND_GATE U15038 ( .I1(n14805), .I2(n15186), .O(n15162) );
  INV_GATE U15039 ( .I1(n15162), .O(n15164) );
  NAND_GATE U15040 ( .I1(A[11]), .I2(B[0]), .O(n15167) );
  NAND_GATE U15041 ( .I1(n15164), .I2(n15167), .O(n14806) );
  NAND_GATE U15042 ( .I1(n15172), .I2(n14806), .O(n14807) );
  INV_GATE U15043 ( .I1(n15167), .O(n15161) );
  NAND_GATE U15044 ( .I1(n15162), .I2(n15161), .O(n15170) );
  NAND_GATE U15045 ( .I1(n14807), .I2(n15170), .O(n15148) );
  INV_GATE U15046 ( .I1(n15148), .O(n15146) );
  NAND_GATE U15047 ( .I1(A[12]), .I2(B[0]), .O(n15153) );
  NAND_GATE U15048 ( .I1(n15146), .I2(n15153), .O(n14808) );
  NAND_GATE U15049 ( .I1(n15149), .I2(n14808), .O(n14809) );
  INV_GATE U15050 ( .I1(n15153), .O(n15147) );
  NAND_GATE U15051 ( .I1(n15148), .I2(n15147), .O(n15157) );
  NAND_GATE U15052 ( .I1(n14809), .I2(n15157), .O(n15133) );
  INV_GATE U15053 ( .I1(n15133), .O(n15135) );
  NAND_GATE U15054 ( .I1(n15135), .I2(n15138), .O(n14810) );
  NAND_GATE U15055 ( .I1(n15143), .I2(n14810), .O(n14811) );
  INV_GATE U15056 ( .I1(n15138), .O(n15132) );
  NAND_GATE U15057 ( .I1(n15133), .I2(n15132), .O(n15141) );
  NAND_GATE U15058 ( .I1(n14811), .I2(n15141), .O(n15119) );
  INV_GATE U15059 ( .I1(n15119), .O(n15117) );
  NAND_GATE U15060 ( .I1(A[14]), .I2(B[0]), .O(n15124) );
  NAND_GATE U15061 ( .I1(n15117), .I2(n15124), .O(n14812) );
  NAND_GATE U15062 ( .I1(n15120), .I2(n14812), .O(n14813) );
  INV_GATE U15063 ( .I1(n15124), .O(n15118) );
  NAND_GATE U15064 ( .I1(n15119), .I2(n15118), .O(n15128) );
  NAND_GATE U15065 ( .I1(n14813), .I2(n15128), .O(n15104) );
  INV_GATE U15066 ( .I1(n15104), .O(n15106) );
  NAND_GATE U15067 ( .I1(A[15]), .I2(B[0]), .O(n15109) );
  NAND_GATE U15068 ( .I1(n15106), .I2(n15109), .O(n14814) );
  NAND_GATE U15069 ( .I1(n15114), .I2(n14814), .O(n14815) );
  INV_GATE U15070 ( .I1(n15109), .O(n15103) );
  NAND_GATE U15071 ( .I1(n15104), .I2(n15103), .O(n15112) );
  NAND_GATE U15072 ( .I1(n14815), .I2(n15112), .O(n15090) );
  INV_GATE U15073 ( .I1(n15090), .O(n15088) );
  NAND_GATE U15074 ( .I1(A[16]), .I2(B[0]), .O(n15095) );
  NAND_GATE U15075 ( .I1(n15088), .I2(n15095), .O(n14816) );
  NAND_GATE U15076 ( .I1(n15091), .I2(n14816), .O(n14817) );
  INV_GATE U15077 ( .I1(n15095), .O(n15089) );
  NAND_GATE U15078 ( .I1(n15090), .I2(n15089), .O(n15099) );
  NAND_GATE U15079 ( .I1(n14817), .I2(n15099), .O(n15075) );
  NAND_GATE U15080 ( .I1(n15077), .I2(n15080), .O(n14818) );
  NAND_GATE U15081 ( .I1(n15085), .I2(n14818), .O(n14819) );
  INV_GATE U15082 ( .I1(n15080), .O(n15074) );
  NAND_GATE U15083 ( .I1(n15075), .I2(n15074), .O(n15083) );
  NAND_GATE U15084 ( .I1(n14819), .I2(n15083), .O(n15061) );
  INV_GATE U15085 ( .I1(n15061), .O(n15059) );
  NAND_GATE U15086 ( .I1(A[18]), .I2(B[0]), .O(n15066) );
  NAND_GATE U15087 ( .I1(n15059), .I2(n15066), .O(n14820) );
  NAND_GATE U15088 ( .I1(n15062), .I2(n14820), .O(n14821) );
  INV_GATE U15089 ( .I1(n15066), .O(n15060) );
  NAND_GATE U15090 ( .I1(n15061), .I2(n15060), .O(n15070) );
  NAND_GATE U15091 ( .I1(n14821), .I2(n15070), .O(n15047) );
  NAND_GATE U15092 ( .I1(A[19]), .I2(B[0]), .O(n15051) );
  NAND_GATE U15093 ( .I1(n15048), .I2(n15051), .O(n14822) );
  NAND_GATE U15094 ( .I1(n15056), .I2(n14822), .O(n14823) );
  INV_GATE U15095 ( .I1(n15051), .O(n15046) );
  NAND_GATE U15096 ( .I1(n15047), .I2(n15046), .O(n15054) );
  NAND_GATE U15097 ( .I1(A[20]), .I2(B[0]), .O(n15038) );
  NAND_GATE U15098 ( .I1(n787), .I2(n15038), .O(n14824) );
  NAND_GATE U15099 ( .I1(n15034), .I2(n14824), .O(n14825) );
  INV_GATE U15100 ( .I1(n15038), .O(n15032) );
  NAND_GATE U15101 ( .I1(n15033), .I2(n15032), .O(n15042) );
  NAND_GATE U15102 ( .I1(n14825), .I2(n15042), .O(n15020) );
  NAND_GATE U15103 ( .I1(A[21]), .I2(B[0]), .O(n15024) );
  NAND_GATE U15104 ( .I1(n22), .I2(n14825), .O(n14826) );
  NAND_GATE U15105 ( .I1(n15029), .I2(n14826), .O(n14827) );
  INV_GATE U15106 ( .I1(n15024), .O(n15019) );
  NAND_GATE U15107 ( .I1(n15020), .I2(n15019), .O(n15027) );
  NAND_GATE U15108 ( .I1(n14827), .I2(n15027), .O(n15007) );
  NAND_GATE U15109 ( .I1(A[22]), .I2(B[0]), .O(n15011) );
  NAND_GATE U15110 ( .I1(n1281), .I2(n15011), .O(n14828) );
  NAND_GATE U15111 ( .I1(n1362), .I2(n14828), .O(n14829) );
  INV_GATE U15112 ( .I1(n15011), .O(n15006) );
  NAND_GATE U15113 ( .I1(n15007), .I2(n15006), .O(n15015) );
  NAND_GATE U15114 ( .I1(A[23]), .I2(B[0]), .O(n14998) );
  NAND_GATE U15115 ( .I1(n828), .I2(n14998), .O(n14830) );
  NAND_GATE U15116 ( .I1(n15003), .I2(n14830), .O(n14831) );
  INV_GATE U15117 ( .I1(n14998), .O(n14993) );
  NAND_GATE U15118 ( .I1(n14831), .I2(n15001), .O(n14980) );
  NAND_GATE U15119 ( .I1(A[24]), .I2(B[0]), .O(n14985) );
  NAND_GATE U15120 ( .I1(n14981), .I2(n14832), .O(n14833) );
  INV_GATE U15121 ( .I1(n14985), .O(n14979) );
  INV_GATE U15122 ( .I1(n14834), .O(n14835) );
  NAND_GATE U15123 ( .I1(n14840), .I2(n14835), .O(n14847) );
  NAND_GATE U15124 ( .I1(n14837), .I2(n14836), .O(n14845) );
  NAND_GATE U15125 ( .I1(n14840), .I2(n14839), .O(n14841) );
  NAND_GATE U15126 ( .I1(n14836), .I2(n14841), .O(n14842) );
  NAND_GATE U15127 ( .I1(n14843), .I2(n14842), .O(n14844) );
  NAND_GATE U15128 ( .I1(n14845), .I2(n14844), .O(n14846) );
  NAND_GATE U15129 ( .I1(n14847), .I2(n14846), .O(n14976) );
  NAND_GATE U15130 ( .I1(n14833), .I2(n1349), .O(n14848) );
  NAND_GATE U15131 ( .I1(n14976), .I2(n14848), .O(n14849) );
  NAND_GATE U15132 ( .I1(n14975), .I2(n14849), .O(n14955) );
  INV_GATE U15133 ( .I1(n14955), .O(n14954) );
  NAND_GATE U15134 ( .I1(A[26]), .I2(B[0]), .O(n14960) );
  NAND_GATE U15135 ( .I1(n14956), .I2(n14850), .O(n14851) );
  NAND_GATE U15136 ( .I1(n14955), .I2(n1298), .O(n14964) );
  NAND_GATE U15137 ( .I1(n14851), .I2(n14964), .O(n14943) );
  NAND_GATE U15138 ( .I1(n14942), .I2(n14943), .O(n14949) );
  NAND_GATE U15139 ( .I1(n14855), .I2(n1319), .O(n14853) );
  NAND_GATE U15140 ( .I1(n14854), .I2(n14853), .O(n14859) );
  NAND_GATE U15141 ( .I1(n14856), .I2(n1357), .O(n14857) );
  NAND_GATE U15142 ( .I1(n14861), .I2(n14860), .O(n14950) );
  NAND_GATE U15143 ( .I1(n14950), .I2(n14862), .O(n14863) );
  NAND_GATE U15144 ( .I1(n14949), .I2(n14863), .O(n14933) );
  NAND_GATE U15145 ( .I1(n14869), .I2(n441), .O(n14866) );
  NAND3_GATE U15146 ( .I1(n14866), .I2(n14865), .I3(n14864), .O(n14873) );
  OR_GATE U15147 ( .I1(n14868), .I2(n14867), .O(n14872) );
  OR_GATE U15148 ( .I1(n14870), .I2(n14869), .O(n14871) );
  NAND3_GATE U15149 ( .I1(n14873), .I2(n14872), .I3(n14871), .O(n14939) );
  NAND_GATE U15150 ( .I1(n14932), .I2(n14874), .O(n14876) );
  NAND3_GATE U15151 ( .I1(n14924), .I2(n14938), .I3(n14876), .O(n14875) );
  NAND_GATE U15152 ( .I1(n14929), .I2(n14875), .O(n14877) );
  INV_GATE U15153 ( .I1(n14924), .O(n14919) );
  NAND_GATE U15154 ( .I1(n14938), .I2(n14876), .O(n14920) );
  NAND_GATE U15155 ( .I1(n14919), .I2(n14920), .O(n14927) );
  NAND_GATE U15156 ( .I1(n14877), .I2(n14927), .O(n14910) );
  OR_GATE U15157 ( .I1(n14878), .I2(n14884), .O(n14881) );
  OR_GATE U15158 ( .I1(n14879), .I2(n14883), .O(n14880) );
  AND_GATE U15159 ( .I1(n14881), .I2(n14880), .O(n14890) );
  INV_GATE U15160 ( .I1(n14884), .O(n14882) );
  NAND_GATE U15161 ( .I1(n14883), .I2(n14882), .O(n14888) );
  INV_GATE U15162 ( .I1(n14883), .O(n14885) );
  NAND_GATE U15163 ( .I1(n14885), .I2(n14884), .O(n14887) );
  NAND3_GATE U15164 ( .I1(n14888), .I2(n14887), .I3(n14886), .O(n14889) );
  NAND_GATE U15165 ( .I1(n348), .I2(n14891), .O(n14893) );
  NAND_GATE U15166 ( .I1(n14907), .I2(n14892), .O(n14894) );
  NAND_GATE U15167 ( .I1(n14916), .I2(n14893), .O(n14898) );
  NAND_GATE U15168 ( .I1(n425), .I2(n14898), .O(n14905) );
  NAND_GATE U15169 ( .I1(n14894), .I2(n14905), .O(n15366) );
  NAND_GATE U15170 ( .I1(n290), .I2(n15366), .O(n14896) );
  AND_GATE U15171 ( .I1(n14896), .I2(n14895), .O(\A1[30] ) );
  INV_GATE U15172 ( .I1(n14898), .O(n14899) );
  NAND_GATE U15173 ( .I1(n384), .I2(n14899), .O(n14897) );
  NAND_GATE U15174 ( .I1(n425), .I2(n14897), .O(n14904) );
  NAND_GATE U15175 ( .I1(n384), .I2(n14898), .O(n14901) );
  NAND_GATE U15176 ( .I1(n14907), .I2(n14899), .O(n14900) );
  NAND3_GATE U15177 ( .I1(n14902), .I2(n14901), .I3(n14900), .O(n14903) );
  NAND_GATE U15178 ( .I1(n14904), .I2(n14903), .O(n14909) );
  INV_GATE U15179 ( .I1(n14905), .O(n14906) );
  NAND_GATE U15180 ( .I1(n14907), .I2(n14906), .O(n14908) );
  NAND_GATE U15181 ( .I1(n14909), .I2(n14908), .O(\A1[29] ) );
  NAND_GATE U15182 ( .I1(n1342), .I2(n14912), .O(n14915) );
  NAND_GATE U15183 ( .I1(n14910), .I2(n348), .O(n14911) );
  NAND_GATE U15184 ( .I1(n14912), .I2(n14911), .O(n14913) );
  OR_GATE U15185 ( .I1(n305), .I2(n14916), .O(n14917) );
  INV_GATE U15186 ( .I1(n14920), .O(n14921) );
  NAND_GATE U15187 ( .I1(n628), .I2(n14921), .O(n14918) );
  NAND_GATE U15188 ( .I1(n14919), .I2(n14918), .O(n14926) );
  NAND_GATE U15189 ( .I1(n628), .I2(n14920), .O(n14923) );
  NAND_GATE U15190 ( .I1(n14929), .I2(n14921), .O(n14922) );
  NAND3_GATE U15191 ( .I1(n14924), .I2(n14923), .I3(n14922), .O(n14925) );
  NAND_GATE U15192 ( .I1(n14926), .I2(n14925), .O(n14931) );
  INV_GATE U15193 ( .I1(n14927), .O(n14928) );
  NAND_GATE U15194 ( .I1(n14929), .I2(n14928), .O(n14930) );
  NAND_GATE U15195 ( .I1(n14931), .I2(n14930), .O(\A1[27] ) );
  NAND_GATE U15196 ( .I1(n14933), .I2(n14932), .O(n14934) );
  NAND_GATE U15197 ( .I1(n14935), .I2(n14934), .O(n14936) );
  OR_GATE U15198 ( .I1(n14939), .I2(n14938), .O(n14940) );
  NAND_GATE U15199 ( .I1(n292), .I2(n1323), .O(n14941) );
  NAND_GATE U15200 ( .I1(n14942), .I2(n14941), .O(n14948) );
  NAND_GATE U15201 ( .I1(n14943), .I2(n1323), .O(n14945) );
  NAND_GATE U15202 ( .I1(n292), .I2(n14950), .O(n14944) );
  NAND3_GATE U15203 ( .I1(n14946), .I2(n14945), .I3(n14944), .O(n14947) );
  NAND_GATE U15204 ( .I1(n14948), .I2(n14947), .O(n14953) );
  INV_GATE U15205 ( .I1(n14949), .O(n14951) );
  NAND_GATE U15206 ( .I1(n14951), .I2(n14950), .O(n14952) );
  NAND_GATE U15207 ( .I1(n14953), .I2(n14952), .O(\A1[25] ) );
  NAND_GATE U15208 ( .I1(n14963), .I2(n14954), .O(n14958) );
  NAND_GATE U15209 ( .I1(n1298), .I2(n14958), .O(n14962) );
  NAND_GATE U15210 ( .I1(n14956), .I2(n14955), .O(n14957) );
  NAND_GATE U15211 ( .I1(n14958), .I2(n14957), .O(n14959) );
  NAND_GATE U15212 ( .I1(n14960), .I2(n14959), .O(n14961) );
  NAND_GATE U15213 ( .I1(n14962), .I2(n14961), .O(n14966) );
  OR_GATE U15214 ( .I1(n14964), .I2(n14963), .O(n14965) );
  NAND_GATE U15215 ( .I1(n14966), .I2(n14965), .O(\A1[24] ) );
  INV_GATE U15216 ( .I1(n14976), .O(n14969) );
  NAND_GATE U15217 ( .I1(n1280), .I2(n14969), .O(n14967) );
  NAND_GATE U15218 ( .I1(n14968), .I2(n14967), .O(n14974) );
  NAND_GATE U15219 ( .I1(n1350), .I2(n14969), .O(n14971) );
  NAND_GATE U15220 ( .I1(n1280), .I2(n14976), .O(n14970) );
  NAND3_GATE U15221 ( .I1(n14972), .I2(n14971), .I3(n14970), .O(n14973) );
  NAND_GATE U15222 ( .I1(n14974), .I2(n14973), .O(n14978) );
  NAND_GATE U15223 ( .I1(n1272), .I2(n14976), .O(n14977) );
  NAND_GATE U15224 ( .I1(n14978), .I2(n14977), .O(\A1[23] ) );
  NAND_GATE U15225 ( .I1(n14988), .I2(n647), .O(n14983) );
  NAND_GATE U15226 ( .I1(n14979), .I2(n14983), .O(n14987) );
  NAND_GATE U15227 ( .I1(n14981), .I2(n14980), .O(n14982) );
  NAND_GATE U15228 ( .I1(n14983), .I2(n14982), .O(n14984) );
  NAND_GATE U15229 ( .I1(n14985), .I2(n14984), .O(n14986) );
  NAND_GATE U15230 ( .I1(n14987), .I2(n14986), .O(n14991) );
  OR_GATE U15231 ( .I1(n14989), .I2(n14988), .O(n14990) );
  NAND_GATE U15232 ( .I1(n14991), .I2(n14990), .O(\A1[22] ) );
  INV_GATE U15233 ( .I1(n15003), .O(n14995) );
  NAND_GATE U15234 ( .I1(n14995), .I2(n828), .O(n14992) );
  NAND_GATE U15235 ( .I1(n14993), .I2(n14992), .O(n15000) );
  NAND_GATE U15236 ( .I1(n14995), .I2(n14994), .O(n14997) );
  NAND_GATE U15237 ( .I1(n15003), .I2(n828), .O(n14996) );
  NAND3_GATE U15238 ( .I1(n14998), .I2(n14997), .I3(n14996), .O(n14999) );
  NAND_GATE U15239 ( .I1(n15000), .I2(n14999), .O(n15005) );
  INV_GATE U15240 ( .I1(n15001), .O(n15002) );
  NAND_GATE U15241 ( .I1(n15003), .I2(n15002), .O(n15004) );
  NAND_GATE U15242 ( .I1(n15005), .I2(n15004), .O(\A1[21] ) );
  NAND_GATE U15243 ( .I1(n15014), .I2(n1281), .O(n15009) );
  NAND_GATE U15244 ( .I1(n15006), .I2(n15009), .O(n15013) );
  NAND_GATE U15245 ( .I1(n1362), .I2(n15007), .O(n15008) );
  NAND_GATE U15246 ( .I1(n15009), .I2(n15008), .O(n15010) );
  NAND_GATE U15247 ( .I1(n15011), .I2(n15010), .O(n15012) );
  NAND_GATE U15248 ( .I1(n15013), .I2(n15012), .O(n15017) );
  OR_GATE U15249 ( .I1(n15015), .I2(n15014), .O(n15016) );
  NAND_GATE U15250 ( .I1(n15017), .I2(n15016), .O(\A1[20] ) );
  NAND_GATE U15251 ( .I1(n1282), .I2(n15021), .O(n15018) );
  NAND_GATE U15252 ( .I1(n15019), .I2(n15018), .O(n15026) );
  NAND_GATE U15253 ( .I1(n1282), .I2(n15020), .O(n15023) );
  NAND_GATE U15254 ( .I1(n15029), .I2(n15021), .O(n15022) );
  NAND3_GATE U15255 ( .I1(n15024), .I2(n15023), .I3(n15022), .O(n15025) );
  NAND_GATE U15256 ( .I1(n15026), .I2(n15025), .O(n15031) );
  INV_GATE U15257 ( .I1(n15027), .O(n15028) );
  NAND_GATE U15258 ( .I1(n15029), .I2(n15028), .O(n15030) );
  NAND_GATE U15259 ( .I1(n15031), .I2(n15030), .O(\A1[19] ) );
  NAND_GATE U15260 ( .I1(n15041), .I2(n787), .O(n15036) );
  NAND_GATE U15261 ( .I1(n15032), .I2(n15036), .O(n15040) );
  NAND_GATE U15262 ( .I1(n15034), .I2(n15033), .O(n15035) );
  NAND_GATE U15263 ( .I1(n15036), .I2(n15035), .O(n15037) );
  NAND_GATE U15264 ( .I1(n15038), .I2(n15037), .O(n15039) );
  NAND_GATE U15265 ( .I1(n15040), .I2(n15039), .O(n15044) );
  OR_GATE U15266 ( .I1(n15042), .I2(n15041), .O(n15043) );
  NAND_GATE U15267 ( .I1(n15044), .I2(n15043), .O(\A1[18] ) );
  NAND_GATE U15268 ( .I1(n648), .I2(n15048), .O(n15045) );
  NAND_GATE U15269 ( .I1(n15046), .I2(n15045), .O(n15053) );
  NAND_GATE U15270 ( .I1(n648), .I2(n15047), .O(n15050) );
  NAND_GATE U15271 ( .I1(n15056), .I2(n15048), .O(n15049) );
  NAND3_GATE U15272 ( .I1(n15051), .I2(n15050), .I3(n15049), .O(n15052) );
  NAND_GATE U15273 ( .I1(n15053), .I2(n15052), .O(n15058) );
  INV_GATE U15274 ( .I1(n15054), .O(n15055) );
  NAND_GATE U15275 ( .I1(n15056), .I2(n15055), .O(n15057) );
  NAND_GATE U15276 ( .I1(n15058), .I2(n15057), .O(\A1[17] ) );
  NAND_GATE U15277 ( .I1(n15069), .I2(n15059), .O(n15064) );
  NAND_GATE U15278 ( .I1(n15060), .I2(n15064), .O(n15068) );
  NAND_GATE U15279 ( .I1(n15062), .I2(n15061), .O(n15063) );
  NAND_GATE U15280 ( .I1(n15064), .I2(n15063), .O(n15065) );
  NAND_GATE U15281 ( .I1(n15066), .I2(n15065), .O(n15067) );
  NAND_GATE U15282 ( .I1(n15068), .I2(n15067), .O(n15072) );
  OR_GATE U15283 ( .I1(n15070), .I2(n15069), .O(n15071) );
  NAND_GATE U15284 ( .I1(n15072), .I2(n15071), .O(\A1[16] ) );
  INV_GATE U15285 ( .I1(n15085), .O(n15076) );
  NAND_GATE U15286 ( .I1(n15076), .I2(n15077), .O(n15073) );
  NAND_GATE U15287 ( .I1(n15074), .I2(n15073), .O(n15082) );
  NAND_GATE U15288 ( .I1(n15076), .I2(n15075), .O(n15079) );
  NAND_GATE U15289 ( .I1(n15085), .I2(n15077), .O(n15078) );
  NAND3_GATE U15290 ( .I1(n15080), .I2(n15079), .I3(n15078), .O(n15081) );
  NAND_GATE U15291 ( .I1(n15082), .I2(n15081), .O(n15087) );
  INV_GATE U15292 ( .I1(n15083), .O(n15084) );
  NAND_GATE U15293 ( .I1(n15085), .I2(n15084), .O(n15086) );
  NAND_GATE U15294 ( .I1(n15087), .I2(n15086), .O(\A1[15] ) );
  NAND_GATE U15295 ( .I1(n15098), .I2(n15088), .O(n15093) );
  NAND_GATE U15296 ( .I1(n15089), .I2(n15093), .O(n15097) );
  NAND_GATE U15297 ( .I1(n15091), .I2(n15090), .O(n15092) );
  NAND_GATE U15298 ( .I1(n15093), .I2(n15092), .O(n15094) );
  NAND_GATE U15299 ( .I1(n15095), .I2(n15094), .O(n15096) );
  NAND_GATE U15300 ( .I1(n15097), .I2(n15096), .O(n15101) );
  OR_GATE U15301 ( .I1(n15099), .I2(n15098), .O(n15100) );
  NAND_GATE U15302 ( .I1(n15101), .I2(n15100), .O(\A1[14] ) );
  INV_GATE U15303 ( .I1(n15114), .O(n15105) );
  NAND_GATE U15304 ( .I1(n15105), .I2(n15106), .O(n15102) );
  NAND_GATE U15305 ( .I1(n15103), .I2(n15102), .O(n15111) );
  NAND_GATE U15306 ( .I1(n15105), .I2(n15104), .O(n15108) );
  NAND_GATE U15307 ( .I1(n15114), .I2(n15106), .O(n15107) );
  NAND3_GATE U15308 ( .I1(n15109), .I2(n15108), .I3(n15107), .O(n15110) );
  NAND_GATE U15309 ( .I1(n15111), .I2(n15110), .O(n15116) );
  INV_GATE U15310 ( .I1(n15112), .O(n15113) );
  NAND_GATE U15311 ( .I1(n15114), .I2(n15113), .O(n15115) );
  NAND_GATE U15312 ( .I1(n15116), .I2(n15115), .O(\A1[13] ) );
  NAND_GATE U15313 ( .I1(n15127), .I2(n15117), .O(n15122) );
  NAND_GATE U15314 ( .I1(n15118), .I2(n15122), .O(n15126) );
  NAND_GATE U15315 ( .I1(n15120), .I2(n15119), .O(n15121) );
  NAND_GATE U15316 ( .I1(n15122), .I2(n15121), .O(n15123) );
  NAND_GATE U15317 ( .I1(n15124), .I2(n15123), .O(n15125) );
  NAND_GATE U15318 ( .I1(n15126), .I2(n15125), .O(n15130) );
  OR_GATE U15319 ( .I1(n15128), .I2(n15127), .O(n15129) );
  NAND_GATE U15320 ( .I1(n15130), .I2(n15129), .O(\A1[12] ) );
  INV_GATE U15321 ( .I1(n15143), .O(n15134) );
  NAND_GATE U15322 ( .I1(n15134), .I2(n15135), .O(n15131) );
  NAND_GATE U15323 ( .I1(n15132), .I2(n15131), .O(n15140) );
  NAND_GATE U15324 ( .I1(n15134), .I2(n15133), .O(n15137) );
  NAND_GATE U15325 ( .I1(n15143), .I2(n15135), .O(n15136) );
  NAND3_GATE U15326 ( .I1(n15138), .I2(n15137), .I3(n15136), .O(n15139) );
  NAND_GATE U15327 ( .I1(n15140), .I2(n15139), .O(n15145) );
  INV_GATE U15328 ( .I1(n15141), .O(n15142) );
  NAND_GATE U15329 ( .I1(n15143), .I2(n15142), .O(n15144) );
  NAND_GATE U15330 ( .I1(n15145), .I2(n15144), .O(\A1[11] ) );
  NAND_GATE U15331 ( .I1(n15156), .I2(n15146), .O(n15151) );
  NAND_GATE U15332 ( .I1(n15147), .I2(n15151), .O(n15155) );
  NAND_GATE U15333 ( .I1(n15149), .I2(n15148), .O(n15150) );
  NAND_GATE U15334 ( .I1(n15151), .I2(n15150), .O(n15152) );
  NAND_GATE U15335 ( .I1(n15153), .I2(n15152), .O(n15154) );
  NAND_GATE U15336 ( .I1(n15155), .I2(n15154), .O(n15159) );
  OR_GATE U15337 ( .I1(n15157), .I2(n15156), .O(n15158) );
  NAND_GATE U15338 ( .I1(n15159), .I2(n15158), .O(\A1[10] ) );
  INV_GATE U15339 ( .I1(n15172), .O(n15163) );
  NAND_GATE U15340 ( .I1(n15163), .I2(n15164), .O(n15160) );
  NAND_GATE U15341 ( .I1(n15161), .I2(n15160), .O(n15169) );
  NAND_GATE U15342 ( .I1(n15163), .I2(n15162), .O(n15166) );
  NAND_GATE U15343 ( .I1(n15172), .I2(n15164), .O(n15165) );
  NAND3_GATE U15344 ( .I1(n15167), .I2(n15166), .I3(n15165), .O(n15168) );
  NAND_GATE U15345 ( .I1(n15169), .I2(n15168), .O(n15174) );
  INV_GATE U15346 ( .I1(n15170), .O(n15171) );
  NAND_GATE U15347 ( .I1(n15172), .I2(n15171), .O(n15173) );
  NAND_GATE U15348 ( .I1(n15174), .I2(n15173), .O(\A1[9] ) );
  NAND_GATE U15349 ( .I1(n15185), .I2(n15175), .O(n15180) );
  NAND_GATE U15350 ( .I1(n15176), .I2(n15180), .O(n15184) );
  NAND_GATE U15351 ( .I1(n15178), .I2(n15177), .O(n15179) );
  NAND_GATE U15352 ( .I1(n15180), .I2(n15179), .O(n15181) );
  NAND_GATE U15353 ( .I1(n15182), .I2(n15181), .O(n15183) );
  NAND_GATE U15354 ( .I1(n15184), .I2(n15183), .O(n15188) );
  OR_GATE U15355 ( .I1(n15186), .I2(n15185), .O(n15187) );
  NAND_GATE U15356 ( .I1(n15188), .I2(n15187), .O(\A1[8] ) );
  INV_GATE U15357 ( .I1(n15201), .O(n15192) );
  NAND_GATE U15358 ( .I1(n15192), .I2(n15193), .O(n15189) );
  NAND_GATE U15359 ( .I1(n15190), .I2(n15189), .O(n15198) );
  NAND_GATE U15360 ( .I1(n15192), .I2(n15191), .O(n15195) );
  NAND_GATE U15361 ( .I1(n15201), .I2(n15193), .O(n15194) );
  NAND3_GATE U15362 ( .I1(n15196), .I2(n15195), .I3(n15194), .O(n15197) );
  NAND_GATE U15363 ( .I1(n15198), .I2(n15197), .O(n15203) );
  INV_GATE U15364 ( .I1(n15199), .O(n15200) );
  NAND_GATE U15365 ( .I1(n15201), .I2(n15200), .O(n15202) );
  NAND_GATE U15366 ( .I1(n15203), .I2(n15202), .O(\A1[7] ) );
  NAND_GATE U15367 ( .I1(n15214), .I2(n15204), .O(n15209) );
  NAND_GATE U15368 ( .I1(n15205), .I2(n15209), .O(n15213) );
  NAND_GATE U15369 ( .I1(n15207), .I2(n15206), .O(n15208) );
  NAND_GATE U15370 ( .I1(n15209), .I2(n15208), .O(n15210) );
  NAND_GATE U15371 ( .I1(n15211), .I2(n15210), .O(n15212) );
  NAND_GATE U15372 ( .I1(n15213), .I2(n15212), .O(n15217) );
  OR_GATE U15373 ( .I1(n15215), .I2(n15214), .O(n15216) );
  NAND_GATE U15374 ( .I1(n15217), .I2(n15216), .O(\A1[6] ) );
  INV_GATE U15375 ( .I1(n15230), .O(n15221) );
  NAND_GATE U15376 ( .I1(n15221), .I2(n15222), .O(n15218) );
  NAND_GATE U15377 ( .I1(n15219), .I2(n15218), .O(n15227) );
  NAND_GATE U15378 ( .I1(n15221), .I2(n15220), .O(n15224) );
  NAND_GATE U15379 ( .I1(n15230), .I2(n15222), .O(n15223) );
  NAND3_GATE U15380 ( .I1(n15225), .I2(n15224), .I3(n15223), .O(n15226) );
  NAND_GATE U15381 ( .I1(n15227), .I2(n15226), .O(n15232) );
  INV_GATE U15382 ( .I1(n15228), .O(n15229) );
  NAND_GATE U15383 ( .I1(n15230), .I2(n15229), .O(n15231) );
  NAND_GATE U15384 ( .I1(n15232), .I2(n15231), .O(\A1[5] ) );
  NAND_GATE U15385 ( .I1(n15243), .I2(n15233), .O(n15238) );
  NAND_GATE U15386 ( .I1(n15234), .I2(n15238), .O(n15242) );
  NAND_GATE U15387 ( .I1(n15236), .I2(n15235), .O(n15237) );
  NAND_GATE U15388 ( .I1(n15238), .I2(n15237), .O(n15239) );
  NAND_GATE U15389 ( .I1(n15240), .I2(n15239), .O(n15241) );
  NAND_GATE U15390 ( .I1(n15242), .I2(n15241), .O(n15246) );
  OR_GATE U15391 ( .I1(n15244), .I2(n15243), .O(n15245) );
  NAND_GATE U15392 ( .I1(n15246), .I2(n15245), .O(\A1[4] ) );
  INV_GATE U15393 ( .I1(n15259), .O(n15250) );
  NAND_GATE U15394 ( .I1(n15250), .I2(n15251), .O(n15247) );
  NAND_GATE U15395 ( .I1(n15248), .I2(n15247), .O(n15256) );
  NAND_GATE U15396 ( .I1(n15250), .I2(n15249), .O(n15253) );
  NAND_GATE U15397 ( .I1(n15259), .I2(n15251), .O(n15252) );
  NAND3_GATE U15398 ( .I1(n15254), .I2(n15253), .I3(n15252), .O(n15255) );
  NAND_GATE U15399 ( .I1(n15256), .I2(n15255), .O(n15261) );
  INV_GATE U15400 ( .I1(n15257), .O(n15258) );
  NAND_GATE U15401 ( .I1(n15259), .I2(n15258), .O(n15260) );
  NAND_GATE U15402 ( .I1(n15261), .I2(n15260), .O(\A1[3] ) );
  NAND_GATE U15403 ( .I1(n15272), .I2(n15262), .O(n15267) );
  NAND_GATE U15404 ( .I1(n15263), .I2(n15267), .O(n15271) );
  NAND_GATE U15405 ( .I1(n15265), .I2(n15264), .O(n15266) );
  NAND_GATE U15406 ( .I1(n15267), .I2(n15266), .O(n15268) );
  NAND_GATE U15407 ( .I1(n15269), .I2(n15268), .O(n15270) );
  NAND_GATE U15408 ( .I1(n15271), .I2(n15270), .O(n15275) );
  OR_GATE U15409 ( .I1(n15273), .I2(n15272), .O(n15274) );
  NAND_GATE U15410 ( .I1(n15275), .I2(n15274), .O(\A1[2] ) );
  INV_GATE U15411 ( .I1(n15288), .O(n15279) );
  NAND_GATE U15412 ( .I1(n15279), .I2(n15280), .O(n15276) );
  NAND_GATE U15413 ( .I1(n15277), .I2(n15276), .O(n15285) );
  NAND_GATE U15414 ( .I1(n15279), .I2(n15278), .O(n15282) );
  NAND_GATE U15415 ( .I1(n15288), .I2(n15280), .O(n15281) );
  NAND3_GATE U15416 ( .I1(n15283), .I2(n15282), .I3(n15281), .O(n15284) );
  NAND_GATE U15417 ( .I1(n15285), .I2(n15284), .O(n15290) );
  INV_GATE U15418 ( .I1(n15286), .O(n15287) );
  NAND_GATE U15419 ( .I1(n15288), .I2(n15287), .O(n15289) );
  NAND_GATE U15420 ( .I1(n15290), .I2(n15289), .O(\A1[1] ) );
  NAND_GATE U15421 ( .I1(n15301), .I2(n15291), .O(n15296) );
  NAND_GATE U15422 ( .I1(n15292), .I2(n15296), .O(n15300) );
  NAND_GATE U15423 ( .I1(n15294), .I2(n15293), .O(n15295) );
  NAND_GATE U15424 ( .I1(n15296), .I2(n15295), .O(n15297) );
  NAND_GATE U15425 ( .I1(n15298), .I2(n15297), .O(n15299) );
  NAND_GATE U15426 ( .I1(n15300), .I2(n15299), .O(n15304) );
  OR_GATE U15427 ( .I1(n15302), .I2(n15301), .O(n15303) );
  NAND_GATE U15428 ( .I1(n15304), .I2(n15303), .O(\A1[0] ) );
  AND_GATE U15429 ( .I1(A[31]), .I2(n15305), .O(\A2[61] ) );
  AND_GATE U15430 ( .I1(n15307), .I2(n15306), .O(\A2[60] ) );
  AND_GATE U15431 ( .I1(n15309), .I2(n15308), .O(\A2[59] ) );
  INV_GATE U15432 ( .I1(n15310), .O(n15376) );
  AND_GATE U15433 ( .I1(n15312), .I2(n15311), .O(\A2[57] ) );
  INV_GATE U15434 ( .I1(n15313), .O(n15373) );
  AND_GATE U15435 ( .I1(n15315), .I2(n15314), .O(\A2[55] ) );
  INV_GATE U15436 ( .I1(n15316), .O(n15374) );
  AND_GATE U15437 ( .I1(n15318), .I2(n15317), .O(\A2[53] ) );
  INV_GATE U15438 ( .I1(n15319), .O(n15372) );
  AND_GATE U15439 ( .I1(n15321), .I2(n15320), .O(\A2[51] ) );
  INV_GATE U15440 ( .I1(n15322), .O(n15370) );
  AND_GATE U15441 ( .I1(n15324), .I2(n15323), .O(\A2[49] ) );
  AND_GATE U15442 ( .I1(n15327), .I2(n15326), .O(\A2[47] ) );
  INV_GATE U15443 ( .I1(n15328), .O(n15375) );
  AND_GATE U15444 ( .I1(n15330), .I2(n15329), .O(\A2[45] ) );
  INV_GATE U15445 ( .I1(n15331), .O(n15369) );
  AND_GATE U15446 ( .I1(n15333), .I2(n15332), .O(\A2[43] ) );
  INV_GATE U15447 ( .I1(n15334), .O(n15368) );
  AND_GATE U15448 ( .I1(n15340), .I2(n15339), .O(\A2[41] ) );
  INV_GATE U15449 ( .I1(n15341), .O(n15367) );
  NAND_GATE U15450 ( .I1(n15343), .I2(n15342), .O(n15344) );
  NAND_GATE U15451 ( .I1(n15345), .I2(n15344), .O(n15346) );
  NAND_GATE U15452 ( .I1(n15347), .I2(n15346), .O(n15348) );
  AND_GATE U15453 ( .I1(n15349), .I2(n15348), .O(\A2[39] ) );
  NAND_GATE U15454 ( .I1(n1220), .I2(n15350), .O(n15353) );
  AND_GATE U15455 ( .I1(n15358), .I2(n15357), .O(\A2[35] ) );
  AND4_GATE U15456 ( .I1(n15362), .I2(n15361), .I3(n15360), .I4(n15359), .O(
        \A2[34] ) );
  AND_GATE U15457 ( .I1(n15364), .I2(n15363), .O(\A2[33] ) );
  AND_GATE U15458 ( .I1(n290), .I2(n15366), .O(\A2[31] ) );
  NAND_GATE U15461 ( .I1(B[1]), .I2(A[0]), .O(n15379) );
  AND_GATE U15462 ( .I1(A[0]), .I2(B[0]), .O(PRODUCT[0]) );
endmodule


module alu_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] ,
         \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] ,
         \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] ,
         \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] ,
         \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] ,
         \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] ,
         \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] ,
         \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] ,
         \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[61] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14839;

  alu_DW01_add_10 FS_1 ( .A({\A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , 
        \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , 
        \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , 
        \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , 
        \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , 
        \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , 
        \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , 
        \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , 
        \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[61] , n14835, n14836, \A2[58] , \A2[57] , \A2[56] , \A2[55] , 
        \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , 
        \A2[47] , \A2[46] , \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , 
        \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , 
        \A2[33] , \A2[32] , \A2[31] , n14834, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2]) );
  AND_GATE U2 ( .I1(n9684), .I2(n9688), .O(n3) );
  AND3_GATE U3 ( .I1(n7238), .I2(n7237), .I3(n7094), .O(n4) );
  NAND3_GATE U4 ( .I1(n6204), .I2(n5600), .I3(n5599), .O(n5) );
  AND3_GATE U5 ( .I1(n10267), .I2(n10266), .I3(n10072), .O(n6) );
  AND3_GATE U6 ( .I1(n5588), .I2(n5587), .I3(n6184), .O(n7) );
  INV_GATE U7 ( .I1(n7), .O(n6199) );
  NAND_GATE U8 ( .I1(n10607), .I2(n11), .O(n8) );
  AND_GATE U9 ( .I1(n8), .I2(n9), .O(n10548) );
  OR_GATE U10 ( .I1(n10), .I2(n10606), .O(n9) );
  INV_GATE U11 ( .I1(n10614), .O(n10) );
  AND_GATE U12 ( .I1(n10605), .I2(n10614), .O(n11) );
  OR_GATE U13 ( .I1(n11092), .I2(n11091), .O(n11096) );
  NAND_GATE U14 ( .I1(n9468), .I2(n15), .O(n12) );
  AND_GATE U15 ( .I1(n12), .I2(n13), .O(n10016) );
  OR_GATE U16 ( .I1(n14), .I2(n9471), .O(n13) );
  INV_GATE U17 ( .I1(n9472), .O(n14) );
  AND_GATE U18 ( .I1(n9469), .I2(n9472), .O(n15) );
  NAND_GATE U19 ( .I1(n10670), .I2(n19), .O(n16) );
  AND_GATE U20 ( .I1(n16), .I2(n17), .O(n11273) );
  OR_GATE U21 ( .I1(n18), .I2(n10672), .O(n17) );
  INV_GATE U22 ( .I1(n10673), .O(n18) );
  AND_GATE U23 ( .I1(n10671), .I2(n10673), .O(n19) );
  OR_GATE U24 ( .I1(n97), .I2(n10027), .O(n9655) );
  AND_GATE U25 ( .I1(n9658), .I2(n640), .O(n20) );
  INV_GATE U26 ( .I1(n20), .O(n9795) );
  NOR_GATE U27 ( .I1(n20), .I2(n9794), .O(n21) );
  OR_GATE U28 ( .I1(n11685), .I2(n11687), .O(n11293) );
  NAND_GATE U29 ( .I1(n11293), .I2(n25), .O(n22) );
  AND_GATE U30 ( .I1(n22), .I2(n23), .O(n11466) );
  OR_GATE U31 ( .I1(n24), .I2(n11682), .O(n23) );
  INV_GATE U32 ( .I1(n11306), .O(n24) );
  AND_GATE U33 ( .I1(n11686), .I2(n11306), .O(n25) );
  NAND3_GATE U34 ( .I1(n10484), .I2(n10485), .I3(n10491), .O(n26) );
  NAND_GATE U35 ( .I1(n10658), .I2(n30), .O(n27) );
  AND_GATE U36 ( .I1(n27), .I2(n28), .O(n11287) );
  OR_GATE U37 ( .I1(n29), .I2(n10661), .O(n28) );
  INV_GATE U38 ( .I1(n10662), .O(n29) );
  AND_GATE U39 ( .I1(n10659), .I2(n10662), .O(n30) );
  NAND_GATE U40 ( .I1(n10660), .I2(n34), .O(n31) );
  AND_GATE U41 ( .I1(n31), .I2(n32), .O(n11284) );
  OR_GATE U42 ( .I1(n33), .I2(n10662), .O(n32) );
  INV_GATE U43 ( .I1(n10840), .O(n33) );
  AND_GATE U44 ( .I1(n10661), .I2(n10840), .O(n34) );
  AND3_GATE U45 ( .I1(n11284), .I2(n10841), .I3(n11283), .O(n35) );
  OR_GATE U46 ( .I1(n7318), .I2(n7317), .O(n7320) );
  NAND_GATE U47 ( .I1(n14286), .I2(n14503), .O(n36) );
  AND_GATE U48 ( .I1(n14487), .I2(n14503), .O(n37) );
  NAND_GATE U49 ( .I1(n14288), .I2(n41), .O(n38) );
  NAND_GATE U50 ( .I1(n38), .I2(n39), .O(n439) );
  OR_GATE U51 ( .I1(n40), .I2(n14468), .O(n39) );
  INV_GATE U52 ( .I1(n14460), .O(n40) );
  AND_GATE U53 ( .I1(n14491), .I2(n14460), .O(n41) );
  NAND_GATE U54 ( .I1(n1368), .I2(n42), .O(n486) );
  NOR_GATE U55 ( .I1(n14425), .I2(n14436), .O(n42) );
  NOR_GATE U56 ( .I1(n8980), .I2(n8979), .O(n43) );
  NAND_GATE U57 ( .I1(n63), .I2(n44), .O(n9138) );
  AND_GATE U58 ( .I1(n64), .I2(n9635), .O(n44) );
  OR_GATE U59 ( .I1(n11325), .I2(n52), .O(n10891) );
  NAND_GATE U60 ( .I1(n12346), .I2(n48), .O(n45) );
  AND_GATE U61 ( .I1(n45), .I2(n46), .O(n13002) );
  OR_GATE U62 ( .I1(n47), .I2(n12348), .O(n46) );
  INV_GATE U63 ( .I1(n12349), .O(n47) );
  AND_GATE U64 ( .I1(n12347), .I2(n12349), .O(n48) );
  OR_GATE U65 ( .I1(n13583), .I2(n13582), .O(n13587) );
  AND3_GATE U66 ( .I1(n12997), .I2(n13404), .I3(n13403), .O(n49) );
  NAND_GATE U67 ( .I1(n11323), .I2(n53), .O(n50) );
  AND_GATE U68 ( .I1(n50), .I2(n51), .O(n11332) );
  OR_GATE U69 ( .I1(n52), .I2(n11325), .O(n51) );
  INV_GATE U70 ( .I1(n11326), .O(n52) );
  AND_GATE U71 ( .I1(n11324), .I2(n11326), .O(n53) );
  NAND_GATE U72 ( .I1(n11336), .I2(n57), .O(n54) );
  AND_GATE U73 ( .I1(n54), .I2(n55), .O(n11447) );
  OR_GATE U74 ( .I1(n56), .I2(n11337), .O(n55) );
  INV_GATE U75 ( .I1(n11446), .O(n56) );
  AND_GATE U76 ( .I1(n11719), .I2(n11446), .O(n57) );
  AND_GATE U77 ( .I1(n10855), .I2(n10506), .O(n58) );
  OR_GATE U78 ( .I1(n1138), .I2(n62), .O(n59) );
  AND_GATE U79 ( .I1(n59), .I2(n60), .O(n10869) );
  OR_GATE U80 ( .I1(n61), .I2(n10855), .O(n60) );
  INV_GATE U81 ( .I1(n10520), .O(n61) );
  OR_GATE U82 ( .I1(n10858), .I2(n61), .O(n62) );
  NAND_GATE U83 ( .I1(n8974), .I2(n65), .O(n63) );
  AND_GATE U84 ( .I1(n63), .I2(n64), .O(n9636) );
  OR_GATE U85 ( .I1(n43), .I2(n8977), .O(n64) );
  AND_GATE U86 ( .I1(n8975), .I2(n8981), .O(n65) );
  NAND_GATE U87 ( .I1(n8978), .I2(n69), .O(n66) );
  AND_GATE U88 ( .I1(n66), .I2(n67), .O(n9634) );
  OR_GATE U89 ( .I1(n68), .I2(n8981), .O(n67) );
  INV_GATE U90 ( .I1(n9137), .O(n68) );
  AND_GATE U91 ( .I1(n8977), .I2(n9137), .O(n69) );
  AND3_GATE U92 ( .I1(n13011), .I2(n13419), .I3(n13418), .O(n70) );
  NAND_GATE U93 ( .I1(n10027), .I2(n71), .O(n96) );
  NOR_GATE U94 ( .I1(n10035), .I2(n97), .O(n71) );
  AND_GATE U95 ( .I1(n9795), .I2(n9666), .O(n72) );
  NAND_GATE U96 ( .I1(n9816), .I2(n76), .O(n73) );
  AND_GATE U97 ( .I1(n73), .I2(n74), .O(n10497) );
  OR_GATE U98 ( .I1(n75), .I2(n9818), .O(n74) );
  INV_GATE U99 ( .I1(n9821), .O(n75) );
  AND_GATE U100 ( .I1(n9817), .I2(n9821), .O(n76) );
  AND_GATE U101 ( .I1(n11338), .I2(n11337), .O(n77) );
  AND3_GATE U102 ( .I1(n12288), .I2(n12211), .I3(n12289), .O(n78) );
  NAND_GATE U103 ( .I1(n11718), .I2(n82), .O(n79) );
  AND_GATE U104 ( .I1(n79), .I2(n80), .O(n11914) );
  OR_GATE U105 ( .I1(n81), .I2(n11716), .O(n80) );
  INV_GATE U106 ( .I1(n11920), .O(n81) );
  AND_GATE U107 ( .I1(n11719), .I2(n11920), .O(n82) );
  AND_GATE U108 ( .I1(n11717), .I2(n11716), .O(n83) );
  INV_GATE U109 ( .I1(n83), .O(n11915) );
  AND3_GATE U110 ( .I1(n11464), .I2(n11463), .I3(n11462), .O(n84) );
  AND_GATE U111 ( .I1(n11951), .I2(n11950), .O(n85) );
  AND3_GATE U112 ( .I1(n13014), .I2(n13015), .I3(n13021), .O(n86) );
  NOR_GATE U113 ( .I1(n70), .I2(n13153), .O(n87) );
  INV_GATE U114 ( .I1(n87), .O(n13162) );
  NAND_GATE U115 ( .I1(n13159), .I2(n90), .O(n88) );
  AND_GATE U116 ( .I1(n88), .I2(n89), .O(n13871) );
  OR_GATE U117 ( .I1(n87), .I2(n13161), .O(n89) );
  AND_GATE U118 ( .I1(n13160), .I2(n13162), .O(n90) );
  NAND_GATE U119 ( .I1(n10028), .I2(n94), .O(n91) );
  NAND_GATE U120 ( .I1(n91), .I2(n92), .O(n645) );
  OR_GATE U121 ( .I1(n93), .I2(n10025), .O(n92) );
  INV_GATE U122 ( .I1(n10037), .O(n93) );
  AND_GATE U123 ( .I1(n10035), .I2(n10037), .O(n94) );
  NAND_GATE U124 ( .I1(n10028), .I2(n98), .O(n95) );
  AND_GATE U125 ( .I1(n95), .I2(n96), .O(n10032) );
  INV_GATE U126 ( .I1(n10031), .O(n97) );
  AND_GATE U127 ( .I1(n10035), .I2(n10031), .O(n98) );
  OR_GATE U128 ( .I1(n9804), .I2(n9799), .O(n99) );
  NAND_GATE U129 ( .I1(n10857), .I2(n10861), .O(n109) );
  NAND_GATE U130 ( .I1(n10030), .I2(n103), .O(n100) );
  AND_GATE U131 ( .I1(n100), .I2(n101), .O(n10297) );
  OR_GATE U132 ( .I1(n102), .I2(n10033), .O(n101) );
  INV_GATE U133 ( .I1(n10036), .O(n102) );
  AND_GATE U134 ( .I1(n10031), .I2(n10036), .O(n103) );
  NAND_GATE U135 ( .I1(n11729), .I2(n104), .O(n154) );
  AND_GATE U136 ( .I1(n11890), .I2(n11728), .O(n104) );
  NAND_GATE U137 ( .I1(n10858), .I2(n105), .O(n107) );
  NOR_GATE U138 ( .I1(n10857), .I2(n108), .O(n105) );
  OR_GATE U139 ( .I1(n10858), .I2(n109), .O(n106) );
  AND_GATE U140 ( .I1(n106), .I2(n107), .O(n10862) );
  INV_GATE U141 ( .I1(n10861), .O(n108) );
  AND_GATE U142 ( .I1(n11682), .I2(n11294), .O(n110) );
  OR_GATE U143 ( .I1(n12182), .I2(n12181), .O(n12185) );
  OR_GATE U144 ( .I1(n11960), .I2(n11953), .O(n111) );
  NAND_GATE U145 ( .I1(n11959), .I2(n115), .O(n112) );
  AND_GATE U146 ( .I1(n112), .I2(n113), .O(n12566) );
  OR_GATE U147 ( .I1(n114), .I2(n11961), .O(n113) );
  INV_GATE U148 ( .I1(n11962), .O(n114) );
  AND_GATE U149 ( .I1(n11960), .I2(n11962), .O(n115) );
  NAND_GATE U150 ( .I1(n11690), .I2(n119), .O(n116) );
  AND_GATE U151 ( .I1(n116), .I2(n117), .O(n11945) );
  OR_GATE U152 ( .I1(n118), .I2(n11693), .O(n117) );
  INV_GATE U153 ( .I1(n11694), .O(n118) );
  AND_GATE U154 ( .I1(n11691), .I2(n11694), .O(n119) );
  NAND_GATE U155 ( .I1(n12576), .I2(n123), .O(n120) );
  AND_GATE U156 ( .I1(n120), .I2(n121), .O(n12738) );
  OR_GATE U157 ( .I1(n122), .I2(n12747), .O(n121) );
  INV_GATE U158 ( .I1(n12591), .O(n122) );
  AND_GATE U159 ( .I1(n12750), .I2(n12591), .O(n123) );
  AND_GATE U160 ( .I1(n13142), .I2(n13027), .O(n124) );
  OR_GATE U161 ( .I1(n13146), .I2(n125), .O(n559) );
  OR_GATE U162 ( .I1(n1282), .I2(n126), .O(n125) );
  INV_GATE U163 ( .I1(n13148), .O(n126) );
  NAND_GATE U164 ( .I1(n14327), .I2(n127), .O(n766) );
  NOR_GATE U165 ( .I1(n14324), .I2(n14326), .O(n127) );
  AND_GATE U166 ( .I1(n14333), .I2(n14332), .O(n128) );
  AND_GATE U167 ( .I1(n11295), .I2(n10854), .O(n129) );
  NAND_GATE U168 ( .I1(n11302), .I2(n133), .O(n130) );
  AND_GATE U169 ( .I1(n130), .I2(n131), .O(n11469) );
  OR_GATE U170 ( .I1(n132), .I2(n11304), .O(n131) );
  INV_GATE U171 ( .I1(n11305), .O(n132) );
  AND_GATE U172 ( .I1(n11303), .I2(n11305), .O(n133) );
  AND_GATE U173 ( .I1(n12578), .I2(n12195), .O(n134) );
  AND_GATE U174 ( .I1(n14349), .I2(n14348), .O(n135) );
  AND3_GATE U175 ( .I1(n13000), .I2(n13001), .I3(n13007), .O(n136) );
  NAND_GATE U176 ( .I1(n13980), .I2(n140), .O(n137) );
  AND_GATE U177 ( .I1(n137), .I2(n138), .O(n13984) );
  OR_GATE U178 ( .I1(n139), .I2(n13982), .O(n138) );
  INV_GATE U179 ( .I1(n13983), .O(n139) );
  AND_GATE U180 ( .I1(n13981), .I2(n13983), .O(n140) );
  AND_GATE U181 ( .I1(n14290), .I2(n14477), .O(n141) );
  NAND_GATE U182 ( .I1(n440), .I2(n142), .O(n443) );
  NOR_GATE U183 ( .I1(n14460), .I2(n14447), .O(n142) );
  NAND_GATE U184 ( .I1(n12623), .I2(n143), .O(n146) );
  AND_GATE U185 ( .I1(n494), .I2(n144), .O(n143) );
  INV_GATE U186 ( .I1(n147), .O(n144) );
  NAND_GATE U187 ( .I1(n12620), .I2(n148), .O(n145) );
  AND_GATE U188 ( .I1(n145), .I2(n146), .O(n12690) );
  INV_GATE U189 ( .I1(n12689), .O(n147) );
  AND_GATE U190 ( .I1(n748), .I2(n12689), .O(n148) );
  NOR_GATE U191 ( .I1(n14464), .I2(n14447), .O(n444) );
  NAND_GATE U192 ( .I1(n628), .I2(n152), .O(n149) );
  AND_GATE U193 ( .I1(n149), .I2(n150), .O(n632) );
  OR_GATE U194 ( .I1(n151), .I2(n14351), .O(n150) );
  INV_GATE U195 ( .I1(n631), .O(n151) );
  AND_GATE U196 ( .I1(n629), .I2(n631), .O(n152) );
  NOR_GATE U197 ( .I1(n11347), .I2(n11340), .O(n467) );
  NAND_GATE U198 ( .I1(n11890), .I2(n153), .O(n155) );
  NOR_GATE U199 ( .I1(n11729), .I2(n11728), .O(n153) );
  AND_GATE U200 ( .I1(n154), .I2(n155), .O(n11732) );
  OR_GATE U201 ( .I1(n11900), .I2(n156), .O(n12284) );
  OR_GATE U202 ( .I1(n11901), .I2(n157), .O(n156) );
  INV_GATE U203 ( .I1(n12283), .O(n157) );
  AND3_GATE U204 ( .I1(n11895), .I2(n11735), .I3(n11734), .O(n158) );
  NAND_GATE U205 ( .I1(n12604), .I2(n159), .O(n1260) );
  NOR_GATE U206 ( .I1(n913), .I2(n12608), .O(n159) );
  AND_GATE U207 ( .I1(n1262), .I2(n12616), .O(n160) );
  OR3_GATE U208 ( .I1(n3591), .I2(n3590), .I3(n3605), .O(n3595) );
  OR3_GATE U209 ( .I1(n161), .I2(n3825), .I3(n731), .O(n3827) );
  INV_GATE U210 ( .I1(n338), .O(n161) );
  OR3_GATE U211 ( .I1(n4721), .I2(n4722), .I3(n4727), .O(n4726) );
  AND_GATE U212 ( .I1(n9254), .I2(n9233), .O(n162) );
  NAND_GATE U213 ( .I1(n8863), .I2(n166), .O(n163) );
  NAND_GATE U214 ( .I1(n163), .I2(n164), .O(n276) );
  OR_GATE U215 ( .I1(n165), .I2(n9233), .O(n164) );
  INV_GATE U216 ( .I1(n9254), .O(n165) );
  AND_GATE U217 ( .I1(n9236), .I2(n9254), .O(n166) );
  NOR_GATE U218 ( .I1(n666), .I2(n510), .O(n511) );
  OR_GATE U219 ( .I1(n731), .I2(n167), .O(n3612) );
  AND_GATE U220 ( .I1(n3731), .I2(n3732), .O(n167) );
  NAND_GATE U221 ( .I1(n3524), .I2(n168), .O(n3525) );
  AND_GATE U222 ( .I1(n2928), .I2(n2927), .O(n168) );
  OR_GATE U223 ( .I1(n3524), .I2(n168), .O(n3526) );
  AND3_GATE U224 ( .I1(n10190), .I2(n10129), .I3(n10128), .O(n169) );
  NAND_GATE U225 ( .I1(n10125), .I2(n9702), .O(n170) );
  NAND_GATE U226 ( .I1(n9749), .I2(n174), .O(n171) );
  AND_GATE U227 ( .I1(n171), .I2(n172), .O(n9752) );
  OR_GATE U228 ( .I1(n173), .I2(n9747), .O(n172) );
  INV_GATE U229 ( .I1(n9751), .O(n173) );
  AND_GATE U230 ( .I1(n742), .I2(n9751), .O(n174) );
  AND3_GATE U231 ( .I1(n3614), .I2(n2961), .I3(n2960), .O(n175) );
  NAND_GATE U232 ( .I1(n5660), .I2(n179), .O(n176) );
  AND_GATE U233 ( .I1(n176), .I2(n177), .O(n5662) );
  OR_GATE U234 ( .I1(n178), .I2(n5658), .O(n177) );
  INV_GATE U235 ( .I1(n5661), .O(n178) );
  AND_GATE U236 ( .I1(n935), .I2(n5661), .O(n179) );
  AND3_GATE U237 ( .I1(n5963), .I2(n5962), .I3(n5667), .O(n180) );
  NAND_GATE U238 ( .I1(n5662), .I2(n184), .O(n181) );
  AND_GATE U239 ( .I1(n181), .I2(n182), .O(n5962) );
  OR_GATE U240 ( .I1(n183), .I2(n5665), .O(n182) );
  INV_GATE U241 ( .I1(n5666), .O(n183) );
  AND_GATE U242 ( .I1(n5663), .I2(n5666), .O(n184) );
  OR_GATE U243 ( .I1(n6328), .I2(n6325), .O(n6331) );
  NAND_GATE U244 ( .I1(n6244), .I2(n6319), .O(n185) );
  NAND_GATE U245 ( .I1(n185), .I2(n186), .O(n188) );
  AND_GATE U246 ( .I1(n187), .I2(n6318), .O(n186) );
  INV_GATE U247 ( .I1(n192), .O(n187) );
  OR_GATE U248 ( .I1(n347), .I2(n188), .O(n191) );
  AND_GATE U249 ( .I1(n6559), .I2(n5971), .O(n189) );
  NAND_GATE U250 ( .I1(n6557), .I2(n193), .O(n190) );
  AND_GATE U251 ( .I1(n190), .I2(n191), .O(n6560) );
  INV_GATE U252 ( .I1(n6559), .O(n192) );
  AND_GATE U253 ( .I1(n189), .I2(n5972), .O(n193) );
  AND_GATE U254 ( .I1(n6847), .I2(n7468), .O(n194) );
  NAND_GATE U255 ( .I1(n7467), .I2(n198), .O(n195) );
  AND_GATE U256 ( .I1(n195), .I2(n196), .O(n7469) );
  OR_GATE U257 ( .I1(n197), .I2(n7465), .O(n196) );
  INV_GATE U258 ( .I1(n7468), .O(n197) );
  AND_GATE U259 ( .I1(n194), .I2(n6846), .O(n198) );
  AND3_GATE U260 ( .I1(n7682), .I2(n7681), .I3(n7474), .O(n199) );
  NAND_GATE U261 ( .I1(n6582), .I2(n203), .O(n200) );
  AND_GATE U262 ( .I1(n200), .I2(n201), .O(n204) );
  OR_GATE U263 ( .I1(n202), .I2(n6584), .O(n201) );
  INV_GATE U264 ( .I1(n6592), .O(n202) );
  AND_GATE U265 ( .I1(n6583), .I2(n6592), .O(n203) );
  NAND_GATE U266 ( .I1(n847), .I2(n204), .O(n206) );
  NAND_GATE U267 ( .I1(n6588), .I2(n207), .O(n205) );
  NAND_GATE U268 ( .I1(n205), .I2(n206), .O(n6815) );
  AND_GATE U269 ( .I1(n6589), .I2(n847), .O(n207) );
  NAND_GATE U270 ( .I1(n10961), .I2(n208), .O(n617) );
  NOR_GATE U271 ( .I1(n10962), .I2(n10959), .O(n208) );
  AND3_GATE U272 ( .I1(n10984), .I2(n10983), .I3(n10982), .O(n209) );
  NAND_GATE U273 ( .I1(n10992), .I2(n213), .O(n210) );
  AND_GATE U274 ( .I1(n210), .I2(n211), .O(n10953) );
  OR_GATE U275 ( .I1(n212), .I2(n10996), .O(n211) );
  INV_GATE U276 ( .I1(n10995), .O(n212) );
  AND_GATE U277 ( .I1(n10952), .I2(n10995), .O(n213) );
  OR_GATE U278 ( .I1(n10978), .I2(n214), .O(n10986) );
  INV_GATE U279 ( .I1(n10980), .O(n214) );
  NAND_GATE U280 ( .I1(n6588), .I2(n218), .O(n215) );
  AND_GATE U281 ( .I1(n215), .I2(n216), .O(n6819) );
  OR_GATE U282 ( .I1(n217), .I2(n6590), .O(n216) );
  INV_GATE U283 ( .I1(n6591), .O(n217) );
  AND_GATE U284 ( .I1(n6589), .I2(n6591), .O(n218) );
  AND_GATE U285 ( .I1(n10979), .I2(n10980), .O(n219) );
  NOR_GATE U286 ( .I1(n4797), .I2(n4800), .O(n220) );
  INV_GATE U287 ( .I1(n220), .O(n4792) );
  AND_GATE U288 ( .I1(n8038), .I2(n8037), .O(n221) );
  NAND_GATE U289 ( .I1(n726), .I2(n222), .O(n225) );
  AND_GATE U290 ( .I1(n8899), .I2(n223), .O(n222) );
  INV_GATE U291 ( .I1(n226), .O(n223) );
  OR_GATE U292 ( .I1(n726), .I2(n227), .O(n224) );
  AND_GATE U293 ( .I1(n224), .I2(n225), .O(n8902) );
  INV_GATE U294 ( .I1(n8901), .O(n226) );
  OR_GATE U295 ( .I1(n8899), .I2(n226), .O(n227) );
  NAND_GATE U296 ( .I1(n4799), .I2(n231), .O(n228) );
  AND_GATE U297 ( .I1(n228), .I2(n229), .O(n5128) );
  OR_GATE U298 ( .I1(n230), .I2(n4801), .O(n229) );
  INV_GATE U299 ( .I1(n4802), .O(n230) );
  AND_GATE U300 ( .I1(n4800), .I2(n4802), .O(n231) );
  OR_GATE U301 ( .I1(n935), .I2(n5659), .O(n5361) );
  OR_GATE U302 ( .I1(n8451), .I2(n8450), .O(n232) );
  OR3_GATE U303 ( .I1(n8440), .I2(n233), .I3(n234), .O(n8443) );
  INV_GATE U304 ( .I1(n8442), .O(n233) );
  INV_GATE U305 ( .I1(n8441), .O(n234) );
  NAND_GATE U306 ( .I1(n8383), .I2(n238), .O(n235) );
  NAND_GATE U307 ( .I1(n235), .I2(n236), .O(n1336) );
  OR_GATE U308 ( .I1(n237), .I2(n8386), .O(n236) );
  INV_GATE U309 ( .I1(n8388), .O(n237) );
  AND_GATE U310 ( .I1(n8384), .I2(n8388), .O(n238) );
  INV_GATE U311 ( .I1(n8364), .O(n239) );
  OR_GATE U312 ( .I1(n8368), .I2(n240), .O(n582) );
  NAND_GATE U313 ( .I1(n8365), .I2(n239), .O(n240) );
  OR_GATE U314 ( .I1(n14812), .I2(n8444), .O(n8438) );
  NAND_GATE U315 ( .I1(n9283), .I2(n244), .O(n241) );
  AND_GATE U316 ( .I1(n241), .I2(n242), .O(n9317) );
  OR_GATE U317 ( .I1(n243), .I2(n9286), .O(n242) );
  INV_GATE U318 ( .I1(n9287), .O(n243) );
  AND_GATE U319 ( .I1(n9284), .I2(n9287), .O(n244) );
  NAND_GATE U320 ( .I1(n9283), .I2(n248), .O(n245) );
  NAND_GATE U321 ( .I1(n245), .I2(n246), .O(n835) );
  OR_GATE U322 ( .I1(n247), .I2(n9286), .O(n246) );
  INV_GATE U323 ( .I1(n9287), .O(n247) );
  AND_GATE U324 ( .I1(n9284), .I2(n9287), .O(n248) );
  NAND_GATE U325 ( .I1(n8872), .I2(n8895), .O(n249) );
  NAND_GATE U326 ( .I1(n249), .I2(n250), .O(n257) );
  AND_GATE U327 ( .I1(n251), .I2(n799), .O(n250) );
  INV_GATE U328 ( .I1(n258), .O(n251) );
  OR_GATE U329 ( .I1(n763), .I2(n8408), .O(n7994) );
  OR_GATE U330 ( .I1(n8424), .I2(n255), .O(n252) );
  AND_GATE U331 ( .I1(n252), .I2(n253), .O(n8428) );
  OR_GATE U332 ( .I1(n254), .I2(n8425), .O(n253) );
  INV_GATE U333 ( .I1(n8427), .O(n254) );
  OR_GATE U334 ( .I1(n824), .I2(n254), .O(n255) );
  OR_GATE U335 ( .I1(n8888), .I2(n259), .O(n256) );
  AND_GATE U336 ( .I1(n256), .I2(n257), .O(n8891) );
  INV_GATE U337 ( .I1(n8890), .O(n258) );
  OR_GATE U338 ( .I1(n799), .I2(n258), .O(n259) );
  NAND_GATE U339 ( .I1(n9720), .I2(n263), .O(n260) );
  AND_GATE U340 ( .I1(n260), .I2(n261), .O(n9727) );
  OR_GATE U341 ( .I1(n262), .I2(n9724), .O(n261) );
  INV_GATE U342 ( .I1(n9726), .O(n262) );
  AND_GATE U343 ( .I1(n9721), .I2(n9726), .O(n263) );
  NAND_GATE U344 ( .I1(n270), .I2(n271), .O(n264) );
  INV_GATE U345 ( .I1(n264), .O(n12601) );
  NAND_GATE U346 ( .I1(n14319), .I2(n268), .O(n265) );
  NAND_GATE U347 ( .I1(n265), .I2(n266), .O(n682) );
  OR_GATE U348 ( .I1(n267), .I2(n448), .O(n266) );
  INV_GATE U349 ( .I1(n14425), .O(n267) );
  AND_GATE U350 ( .I1(n14450), .I2(n14425), .O(n268) );
  AND_GATE U351 ( .I1(n12297), .I2(n12209), .O(n269) );
  OR_GATE U352 ( .I1(n12288), .I2(n273), .O(n270) );
  OR_GATE U353 ( .I1(n272), .I2(n12290), .O(n271) );
  INV_GATE U354 ( .I1(n13046), .O(n272) );
  OR_GATE U355 ( .I1(n12292), .I2(n272), .O(n273) );
  OR_GATE U356 ( .I1(n1374), .I2(n12285), .O(n12287) );
  OR_GATE U357 ( .I1(n12293), .I2(n269), .O(n12295) );
  AND3_GATE U358 ( .I1(n13538), .I2(n13537), .I3(n13536), .O(n274) );
  AND_GATE U359 ( .I1(n162), .I2(n8864), .O(n275) );
  NAND_GATE U360 ( .I1(n7215), .I2(n278), .O(n277) );
  NOR_GATE U361 ( .I1(n7212), .I2(n7218), .O(n278) );
  NOR_GATE U362 ( .I1(n10899), .I2(n10898), .O(n279) );
  INV_GATE U363 ( .I1(n279), .O(n10902) );
  AND_GATE U364 ( .I1(n12639), .I2(n12638), .O(n280) );
  NAND_GATE U365 ( .I1(n5594), .I2(n284), .O(n281) );
  AND_GATE U366 ( .I1(n281), .I2(n282), .O(n6208) );
  OR_GATE U367 ( .I1(n283), .I2(n5597), .O(n282) );
  INV_GATE U368 ( .I1(n6207), .O(n283) );
  AND_GATE U369 ( .I1(n5595), .I2(n6207), .O(n284) );
  NAND_GATE U370 ( .I1(n2907), .I2(n2908), .O(n285) );
  AND3_GATE U371 ( .I1(n11840), .I2(n11772), .I3(n11771), .O(n286) );
  NAND_GATE U372 ( .I1(n10914), .I2(n10913), .O(n287) );
  NAND_GATE U373 ( .I1(n10056), .I2(n291), .O(n288) );
  AND_GATE U374 ( .I1(n288), .I2(n289), .O(n10267) );
  OR_GATE U375 ( .I1(n290), .I2(n10529), .O(n289) );
  INV_GATE U376 ( .I1(n10068), .O(n290) );
  AND_GATE U377 ( .I1(n10532), .I2(n10068), .O(n291) );
  AND_GATE U378 ( .I1(n8294), .I2(n8293), .O(n292) );
  AND3_GATE U379 ( .I1(n7242), .I2(n7241), .I3(n7240), .O(n293) );
  AND_GATE U380 ( .I1(n7395), .I2(n7078), .O(n294) );
  NAND_GATE U381 ( .I1(n8561), .I2(n298), .O(n295) );
  AND_GATE U382 ( .I1(n295), .I2(n296), .O(n8554) );
  OR_GATE U383 ( .I1(n297), .I2(n8557), .O(n296) );
  INV_GATE U384 ( .I1(n8303), .O(n297) );
  AND_GATE U385 ( .I1(n8555), .I2(n8303), .O(n298) );
  AND_GATE U386 ( .I1(n5318), .I2(n5317), .O(n299) );
  AND3_GATE U387 ( .I1(n11453), .I2(n11321), .I3(n11452), .O(n300) );
  INV_GATE U388 ( .I1(n300), .O(n11719) );
  AND_GATE U389 ( .I1(n1487), .I2(n1486), .O(n301) );
  INV_GATE U390 ( .I1(n301), .O(n1845) );
  AND_GATE U391 ( .I1(n5172), .I2(n5171), .O(n302) );
  AND_GATE U392 ( .I1(n3823), .I2(n3822), .O(n303) );
  AND3_GATE U393 ( .I1(n2899), .I2(n2898), .I3(n3573), .O(n304) );
  AND_GATE U394 ( .I1(n8339), .I2(n7985), .O(n305) );
  AND_GATE U395 ( .I1(n7456), .I2(n7455), .O(n306) );
  AND3_GATE U396 ( .I1(n7122), .I2(n7121), .I3(n7120), .O(n307) );
  NAND_GATE U397 ( .I1(n4446), .I2(n4445), .O(n308) );
  AND3_GATE U398 ( .I1(n7726), .I2(n7725), .I3(n7458), .O(n309) );
  AND3_GATE U399 ( .I1(n6015), .I2(n6014), .I3(n6013), .O(n310) );
  AND_GATE U400 ( .I1(n4469), .I2(n4468), .O(n311) );
  AND3_GATE U401 ( .I1(n3534), .I2(n3533), .I3(n3532), .O(n312) );
  OR_GATE U402 ( .I1(n313), .I2(n4809), .O(n4811) );
  INV_GATE U403 ( .I1(n4807), .O(n313) );
  NAND_GATE U404 ( .I1(n6631), .I2(n317), .O(n314) );
  AND_GATE U405 ( .I1(n314), .I2(n315), .O(n6787) );
  OR_GATE U406 ( .I1(n316), .I2(n6634), .O(n315) );
  INV_GATE U407 ( .I1(n6635), .O(n316) );
  AND_GATE U408 ( .I1(n6632), .I2(n6635), .O(n317) );
  AND_GATE U409 ( .I1(n6793), .I2(n6792), .O(n318) );
  AND_GATE U410 ( .I1(n2073), .I2(n2072), .O(n319) );
  AND_GATE U411 ( .I1(n1836), .I2(n1835), .O(n320) );
  AND3_GATE U412 ( .I1(n3462), .I2(n3461), .I3(n3022), .O(n321) );
  AND3_GATE U413 ( .I1(n3496), .I2(n2977), .I3(n3499), .O(n322) );
  NAND_GATE U414 ( .I1(n3919), .I2(n325), .O(n323) );
  AND_GATE U415 ( .I1(n323), .I2(n324), .O(n4275) );
  OR_GATE U416 ( .I1(n4281), .I2(n3922), .O(n324) );
  AND_GATE U417 ( .I1(n3920), .I2(n3923), .O(n325) );
  AND_GATE U418 ( .I1(n2732), .I2(n2731), .O(n326) );
  NAND_GATE U419 ( .I1(n6553), .I2(n6247), .O(n327) );
  AND3_GATE U420 ( .I1(n3519), .I2(n2959), .I3(n2958), .O(n328) );
  OR_GATE U421 ( .I1(n934), .I2(n329), .O(n3632) );
  INV_GATE U422 ( .I1(n3887), .O(n329) );
  AND3_GATE U423 ( .I1(n5150), .I2(n5149), .I3(n5148), .O(n330) );
  AND_GATE U424 ( .I1(n2703), .I2(n2702), .O(n331) );
  AND_GATE U425 ( .I1(n5653), .I2(n5652), .O(n332) );
  AND3_GATE U426 ( .I1(n4334), .I2(n4333), .I3(n3855), .O(n333) );
  NAND_GATE U427 ( .I1(n4472), .I2(n337), .O(n334) );
  NAND_GATE U428 ( .I1(n334), .I2(n335), .O(n900) );
  OR_GATE U429 ( .I1(n336), .I2(n4768), .O(n335) );
  INV_GATE U430 ( .I1(n4569), .O(n336) );
  AND_GATE U431 ( .I1(n4769), .I2(n4569), .O(n337) );
  AND3_GATE U432 ( .I1(n3523), .I2(n3522), .I3(n3521), .O(n338) );
  AND_GATE U433 ( .I1(n3589), .I2(n2938), .O(n339) );
  OR_GATE U434 ( .I1(n5143), .I2(n909), .O(n5145) );
  AND_GATE U435 ( .I1(n1847), .I2(n1846), .O(n340) );
  INV_GATE U436 ( .I1(n340), .O(n1984) );
  OR_GATE U437 ( .I1(n1375), .I2(n341), .O(n2747) );
  AND_GATE U438 ( .I1(n2867), .I2(n2866), .O(n341) );
  NAND_GATE U439 ( .I1(n5647), .I2(n345), .O(n342) );
  AND_GATE U440 ( .I1(n342), .I2(n343), .O(n5973) );
  OR_GATE U441 ( .I1(n344), .I2(n5652), .O(n343) );
  INV_GATE U442 ( .I1(n5654), .O(n344) );
  AND_GATE U443 ( .I1(n5648), .I2(n5654), .O(n345) );
  INV_GATE U444 ( .I1(n1400), .O(n346) );
  AND_GATE U445 ( .I1(n5972), .I2(n5971), .O(n347) );
  AND_GATE U446 ( .I1(n2940), .I2(n2939), .O(n348) );
  AND_GATE U447 ( .I1(n1867), .I2(n1866), .O(n349) );
  AND_GATE U448 ( .I1(n12236), .I2(n12235), .O(n350) );
  AND3_GATE U449 ( .I1(n8851), .I2(n8852), .I3(n8853), .O(n351) );
  AND3_GATE U450 ( .I1(n8855), .I2(n8854), .I3(n9204), .O(n352) );
  INV_GATE U451 ( .I1(n352), .O(n8919) );
  AND3_GATE U452 ( .I1(n6897), .I2(n6896), .I3(n6895), .O(n353) );
  AND_GATE U453 ( .I1(n7442), .I2(n7441), .O(n354) );
  AND_GATE U454 ( .I1(n5473), .I2(n5472), .O(n355) );
  AND_GATE U455 ( .I1(n4699), .I2(n4698), .O(n356) );
  NAND_GATE U456 ( .I1(n11409), .I2(n11408), .O(n357) );
  AND3_GATE U457 ( .I1(n9394), .I2(n9213), .I3(n9397), .O(n358) );
  AND3_GATE U458 ( .I1(n9369), .I2(n9370), .I3(n9382), .O(n359) );
  NAND_GATE U459 ( .I1(n6535), .I2(n6534), .O(n360) );
  AND_GATE U460 ( .I1(n5338), .I2(n5337), .O(n361) );
  OR_GATE U461 ( .I1(n1303), .I2(n4736), .O(n4734) );
  AND3_GATE U462 ( .I1(n9634), .I2(n9138), .I3(n9637), .O(n362) );
  NAND_GATE U463 ( .I1(n1425), .I2(A[9]), .O(n363) );
  NAND_GATE U464 ( .I1(n8745), .I2(n364), .O(n8749) );
  INV_GATE U465 ( .I1(n363), .O(n364) );
  OR_GATE U466 ( .I1(n365), .I2(n10242), .O(n10246) );
  INV_GATE U467 ( .I1(n10243), .O(n365) );
  AND_GATE U468 ( .I1(n5701), .I2(n5370), .O(n366) );
  NAND_GATE U469 ( .I1(n5099), .I2(n5098), .O(n367) );
  AND_GATE U470 ( .I1(n2631), .I2(n2630), .O(n368) );
  AND3_GATE U471 ( .I1(n6749), .I2(n6748), .I3(n6684), .O(n369) );
  AND3_GATE U472 ( .I1(n3482), .I2(n3483), .I3(n2991), .O(n370) );
  INV_GATE U473 ( .I1(n370), .O(n3477) );
  OR3_GATE U474 ( .I1(n21), .I2(n371), .I3(n9799), .O(n9802) );
  INV_GATE U475 ( .I1(n9800), .O(n371) );
  AND3_GATE U476 ( .I1(n11419), .I2(n11382), .I3(n11381), .O(n372) );
  INV_GATE U477 ( .I1(n372), .O(n11849) );
  OR_GATE U478 ( .I1(n11857), .I2(n376), .O(n373) );
  AND_GATE U479 ( .I1(n373), .I2(n374), .O(n12224) );
  OR_GATE U480 ( .I1(n375), .I2(n11865), .O(n374) );
  INV_GATE U481 ( .I1(n12258), .O(n375) );
  OR_GATE U482 ( .I1(n11858), .I2(n375), .O(n376) );
  NAND_GATE U483 ( .I1(n9761), .I2(n380), .O(n377) );
  AND_GATE U484 ( .I1(n377), .I2(n378), .O(n9768) );
  OR_GATE U485 ( .I1(n379), .I2(n9759), .O(n378) );
  INV_GATE U486 ( .I1(n9691), .O(n379) );
  AND_GATE U487 ( .I1(n9758), .I2(n9691), .O(n380) );
  OR_GATE U488 ( .I1(n1108), .I2(n384), .O(n381) );
  AND_GATE U489 ( .I1(n381), .I2(n382), .O(n8603) );
  OR_GATE U490 ( .I1(n383), .I2(n8595), .O(n382) );
  INV_GATE U491 ( .I1(n8297), .O(n383) );
  OR_GATE U492 ( .I1(n1362), .I2(n383), .O(n384) );
  AND_GATE U493 ( .I1(n4706), .I2(n4710), .O(n385) );
  AND_GATE U494 ( .I1(n3809), .I2(n3808), .O(n386) );
  NAND3_GATE U495 ( .I1(n4701), .I2(n4702), .I3(n4700), .O(n387) );
  OR_GATE U496 ( .I1(n5287), .I2(n5289), .O(n388) );
  AND3_GATE U497 ( .I1(n3794), .I2(n3792), .I3(n3793), .O(n389) );
  AND3_GATE U498 ( .I1(n11430), .I2(n11429), .I3(n11428), .O(n390) );
  AND_GATE U499 ( .I1(n10546), .I2(n10545), .O(n391) );
  AND3_GATE U500 ( .I1(n10619), .I2(n10618), .I3(n10617), .O(n392) );
  AND3_GATE U501 ( .I1(n9792), .I2(n9791), .I3(n9790), .O(n393) );
  AND_GATE U502 ( .I1(n8957), .I2(n8956), .O(n394) );
  NAND3_GATE U503 ( .I1(n8280), .I2(n8279), .I3(n8814), .O(n395) );
  NAND3_GATE U504 ( .I1(n7258), .I2(n7257), .I3(n7256), .O(n396) );
  AND_GATE U505 ( .I1(n10529), .I2(n10057), .O(n397) );
  AND3_GATE U506 ( .I1(n4632), .I2(n4631), .I3(n4630), .O(n398) );
  AND3_GATE U507 ( .I1(n12282), .I2(n12281), .I3(n12280), .O(n399) );
  OR3_GATE U508 ( .I1(n400), .I2(n401), .I3(n6372), .O(n6375) );
  INV_GATE U509 ( .I1(n6370), .O(n400) );
  INV_GATE U510 ( .I1(n6225), .O(n401) );
  NOR_GATE U511 ( .I1(n5863), .I2(n5871), .O(n402) );
  AND_GATE U512 ( .I1(n5851), .I2(n5850), .O(n403) );
  AND_GATE U513 ( .I1(n7606), .I2(n7605), .O(n404) );
  AND3_GATE U514 ( .I1(n5407), .I2(n5400), .I3(n5399), .O(n405) );
  AND_GATE U515 ( .I1(n4140), .I2(n4139), .O(n406) );
  AND3_GATE U516 ( .I1(n3688), .I2(n3681), .I3(n3680), .O(n407) );
  AND_GATE U517 ( .I1(n2434), .I2(n2433), .O(n408) );
  AND_GATE U518 ( .I1(n2416), .I2(n2415), .O(n409) );
  AND3_GATE U519 ( .I1(n1936), .I2(n1935), .I3(n1934), .O(n410) );
  AND3_GATE U520 ( .I1(n11836), .I2(n715), .I3(n11768), .O(n411) );
  AND_GATE U521 ( .I1(n13484), .I2(n13485), .O(n412) );
  AND_GATE U522 ( .I1(n3598), .I2(n3597), .O(n413) );
  AND3_GATE U523 ( .I1(B[24]), .I2(B[25]), .I3(n1254), .O(n414) );
  AND3_GATE U524 ( .I1(n6734), .I2(n6733), .I3(n6732), .O(n415) );
  OR_GATE U525 ( .I1(n683), .I2(n14429), .O(n14421) );
  OR_GATE U526 ( .I1(n683), .I2(n128), .O(n14423) );
  NAND_GATE U527 ( .I1(n13897), .I2(n419), .O(n416) );
  AND_GATE U528 ( .I1(n416), .I2(n417), .O(n13962) );
  OR_GATE U529 ( .I1(n418), .I2(n13898), .O(n417) );
  INV_GATE U530 ( .I1(n13961), .O(n418) );
  AND_GATE U531 ( .I1(n13896), .I2(n13961), .O(n419) );
  OR_GATE U532 ( .I1(n13894), .I2(n13961), .O(n13895) );
  OR_GATE U533 ( .I1(n14322), .I2(n420), .O(n14333) );
  INV_GATE U534 ( .I1(n14327), .O(n420) );
  NAND_GATE U535 ( .I1(n13550), .I2(n421), .O(n544) );
  NOR_GATE U536 ( .I1(n13553), .I2(n13551), .O(n421) );
  OR_GATE U537 ( .I1(n422), .I2(n13953), .O(n13958) );
  INV_GATE U538 ( .I1(n13954), .O(n422) );
  NAND_GATE U539 ( .I1(n13550), .I2(n961), .O(n13554) );
  AND_GATE U540 ( .I1(n14329), .I2(n14325), .O(n423) );
  NAND_GATE U541 ( .I1(n14326), .I2(n423), .O(n767) );
  NAND_GATE U542 ( .I1(n14334), .I2(n426), .O(n424) );
  AND_GATE U543 ( .I1(n424), .I2(n425), .O(n14418) );
  OR_GATE U544 ( .I1(n14416), .I2(n14428), .O(n425) );
  AND_GATE U545 ( .I1(n14429), .I2(n14411), .O(n426) );
  NAND_GATE U546 ( .I1(n14415), .I2(n430), .O(n427) );
  AND_GATE U547 ( .I1(n427), .I2(n428), .O(\A1[26] ) );
  OR_GATE U548 ( .I1(n429), .I2(n14417), .O(n428) );
  INV_GATE U549 ( .I1(n14420), .O(n429) );
  AND_GATE U550 ( .I1(n14416), .I2(n14420), .O(n430) );
  NAND_GATE U551 ( .I1(n84), .I2(n431), .O(n433) );
  AND_GATE U552 ( .I1(n12199), .I2(n12201), .O(n431) );
  OR_GATE U553 ( .I1(n84), .I2(n435), .O(n432) );
  AND_GATE U554 ( .I1(n432), .I2(n433), .O(n12202) );
  INV_GATE U555 ( .I1(n12201), .O(n434) );
  OR_GATE U556 ( .I1(n12199), .I2(n434), .O(n435) );
  OR_GATE U557 ( .I1(n13466), .I2(n436), .O(n13478) );
  INV_GATE U558 ( .I1(n13469), .O(n436) );
  OR_GATE U559 ( .I1(n14538), .I2(n14537), .O(n14279) );
  OR_GATE U560 ( .I1(n14002), .I2(n14001), .O(n14006) );
  AND_GATE U561 ( .I1(n14013), .I2(n14012), .O(n437) );
  AND3_GATE U562 ( .I1(n11930), .I2(n11929), .I3(n11928), .O(n438) );
  NAND_GATE U563 ( .I1(n14290), .I2(n14477), .O(n440) );
  OR_GATE U564 ( .I1(n13573), .I2(n441), .O(n541) );
  NAND_GATE U565 ( .I1(n13571), .I2(n13575), .O(n441) );
  OR_GATE U566 ( .I1(n13573), .I2(n13572), .O(n13574) );
  NAND_GATE U567 ( .I1(n14301), .I2(n444), .O(n442) );
  AND_GATE U568 ( .I1(n442), .I2(n443), .O(n14450) );
  AND_GATE U569 ( .I1(n14463), .I2(n14302), .O(n445) );
  NAND_GATE U570 ( .I1(n14302), .I2(n449), .O(n446) );
  NAND_GATE U571 ( .I1(n446), .I2(n447), .O(n1353) );
  OR_GATE U572 ( .I1(n448), .I2(n529), .O(n447) );
  INV_GATE U573 ( .I1(n14436), .O(n448) );
  AND_GATE U574 ( .I1(n14463), .I2(n14436), .O(n449) );
  NAND_GATE U575 ( .I1(n14320), .I2(n450), .O(n485) );
  AND_GATE U576 ( .I1(n14422), .I2(n484), .O(n450) );
  NOR_GATE U577 ( .I1(n12749), .I2(n12752), .O(n451) );
  INV_GATE U578 ( .I1(n451), .O(n12747) );
  OR_GATE U579 ( .I1(n936), .I2(n14395), .O(n14389) );
  NAND_GATE U580 ( .I1(n14391), .I2(n455), .O(n452) );
  AND_GATE U581 ( .I1(n452), .I2(n453), .O(\A1[28] ) );
  OR_GATE U582 ( .I1(n454), .I2(n14393), .O(n453) );
  INV_GATE U583 ( .I1(n14396), .O(n454) );
  AND_GATE U584 ( .I1(n14392), .I2(n14396), .O(n455) );
  OR3_GATE U585 ( .I1(n456), .I2(n457), .I3(n13921), .O(n13927) );
  AND3_GATE U586 ( .I1(n13925), .I2(n13926), .I3(n970), .O(n456) );
  AND3_GATE U587 ( .I1(n727), .I2(n13926), .I3(n970), .O(n457) );
  NAND_GATE U588 ( .I1(n12330), .I2(n458), .O(n460) );
  NOR_GATE U589 ( .I1(n12331), .I2(n461), .O(n458) );
  NAND_GATE U590 ( .I1(n85), .I2(n462), .O(n459) );
  AND_GATE U591 ( .I1(n459), .I2(n460), .O(n12334) );
  INV_GATE U592 ( .I1(n12333), .O(n461) );
  AND_GATE U593 ( .I1(n12331), .I2(n12333), .O(n462) );
  OR_GATE U594 ( .I1(n12749), .I2(n463), .O(n555) );
  NAND_GATE U595 ( .I1(n12750), .I2(n12752), .O(n463) );
  AND_GATE U596 ( .I1(n11343), .I2(n11347), .O(n464) );
  NAND_GATE U597 ( .I1(n638), .I2(n464), .O(n466) );
  NAND_GATE U598 ( .I1(n11342), .I2(n467), .O(n465) );
  AND_GATE U599 ( .I1(n465), .I2(n466), .O(n11344) );
  OR_GATE U600 ( .I1(n10898), .I2(n468), .O(n859) );
  NAND_GATE U601 ( .I1(n10903), .I2(n10899), .O(n468) );
  AND_GATE U602 ( .I1(n11346), .I2(n10895), .O(n469) );
  NOR_GATE U603 ( .I1(n1383), .I2(n1099), .O(n470) );
  AND_GATE U604 ( .I1(n11723), .I2(n473), .O(n471) );
  NOR_GATE U605 ( .I1(n471), .I2(n472), .O(n11895) );
  AND_GATE U606 ( .I1(n11896), .I2(n1383), .O(n472) );
  AND_GATE U607 ( .I1(n11911), .I2(n11896), .O(n473) );
  AND_GATE U608 ( .I1(n12585), .I2(n12586), .O(n474) );
  NAND_GATE U609 ( .I1(n12584), .I2(n474), .O(n477) );
  AND_GATE U610 ( .I1(n11704), .I2(n11707), .O(n475) );
  NAND_GATE U611 ( .I1(n11703), .I2(n475), .O(n1341) );
  NAND_GATE U612 ( .I1(n12582), .I2(n478), .O(n476) );
  AND_GATE U613 ( .I1(n476), .I2(n477), .O(n12587) );
  AND_GATE U614 ( .I1(n12583), .I2(n12586), .O(n478) );
  AND_GATE U615 ( .I1(n12747), .I2(n12577), .O(n479) );
  NAND_GATE U616 ( .I1(n13146), .I2(n480), .O(n558) );
  AND_GATE U617 ( .I1(n13148), .I2(n1282), .O(n480) );
  NAND_GATE U618 ( .I1(n10898), .I2(n481), .O(n860) );
  NOR_GATE U619 ( .I1(n10903), .I2(n482), .O(n481) );
  INV_GATE U620 ( .I1(n10899), .O(n482) );
  AND_GATE U621 ( .I1(n12284), .I2(n12214), .O(n483) );
  AND_GATE U622 ( .I1(n13975), .I2(n13974), .O(n484) );
  AND_GATE U623 ( .I1(n485), .I2(n486), .O(n14428) );
  AND_GATE U624 ( .I1(n13028), .I2(n12594), .O(n487) );
  OR_GATE U625 ( .I1(n13454), .I2(n13042), .O(n785) );
  OR_GATE U626 ( .I1(n488), .I2(n13454), .O(n13451) );
  INV_GATE U627 ( .I1(n13453), .O(n488) );
  OR_GATE U628 ( .I1(n438), .I2(n12300), .O(n12298) );
  AND3_GATE U629 ( .I1(n12730), .I2(n12596), .I3(n12733), .O(n489) );
  AND_GATE U630 ( .I1(n13455), .I2(n13456), .O(n490) );
  NAND_GATE U631 ( .I1(n13454), .I2(n490), .O(n786) );
  AND_GATE U632 ( .I1(n13444), .I2(n13569), .O(n491) );
  NAND_GATE U633 ( .I1(n13573), .I2(n492), .O(n542) );
  NOR_GATE U634 ( .I1(n13571), .I2(n493), .O(n492) );
  INV_GATE U635 ( .I1(n13575), .O(n493) );
  NAND3_GATE U636 ( .I1(n12216), .I2(n12215), .I3(n12609), .O(n494) );
  AND_GATE U637 ( .I1(n11755), .I2(n11754), .O(n495) );
  OR_GATE U638 ( .I1(n11874), .I2(n495), .O(n11884) );
  NAND_GATE U639 ( .I1(n11888), .I2(n498), .O(n496) );
  AND_GATE U640 ( .I1(n496), .I2(n497), .O(n12611) );
  OR_GATE U641 ( .I1(n11886), .I2(n11889), .O(n497) );
  AND_GATE U642 ( .I1(n158), .I2(n12607), .O(n498) );
  NAND_GATE U643 ( .I1(n5630), .I2(n499), .O(n501) );
  AND_GATE U644 ( .I1(n5635), .I2(n5631), .O(n499) );
  OR_GATE U645 ( .I1(n5630), .I2(n503), .O(n500) );
  AND_GATE U646 ( .I1(n500), .I2(n501), .O(n5632) );
  INV_GATE U647 ( .I1(n5631), .O(n502) );
  OR_GATE U648 ( .I1(n5635), .I2(n502), .O(n503) );
  OR_GATE U649 ( .I1(n8314), .I2(n8309), .O(n8316) );
  AND_GATE U650 ( .I1(n703), .I2(n7188), .O(n504) );
  NAND_GATE U651 ( .I1(n7192), .I2(n504), .O(n585) );
  AND3_GATE U652 ( .I1(n6863), .I2(n6862), .I3(n6550), .O(n505) );
  AND_GATE U653 ( .I1(n6315), .I2(n6331), .O(n506) );
  NAND_GATE U654 ( .I1(n6314), .I2(n507), .O(n1377) );
  AND_GATE U655 ( .I1(n506), .I2(n6243), .O(n507) );
  NAND_GATE U656 ( .I1(n6242), .I2(n511), .O(n508) );
  NAND_GATE U657 ( .I1(n508), .I2(n509), .O(n1378) );
  OR_GATE U658 ( .I1(n510), .I2(n6331), .O(n509) );
  INV_GATE U659 ( .I1(n6315), .O(n510) );
  NAND_GATE U660 ( .I1(n7469), .I2(n514), .O(n512) );
  AND_GATE U661 ( .I1(n512), .I2(n513), .O(n7681) );
  OR_GATE U662 ( .I1(n7687), .I2(n7472), .O(n513) );
  AND_GATE U663 ( .I1(n7470), .I2(n7473), .O(n514) );
  NAND_GATE U664 ( .I1(n8902), .I2(n517), .O(n515) );
  AND_GATE U665 ( .I1(n515), .I2(n516), .O(n9301) );
  OR_GATE U666 ( .I1(n9307), .I2(n8905), .O(n516) );
  AND_GATE U667 ( .I1(n8903), .I2(n9290), .O(n517) );
  OR3_GATE U668 ( .I1(n9296), .I2(n518), .I3(n519), .O(n9299) );
  INV_GATE U669 ( .I1(n9298), .O(n518) );
  INV_GATE U670 ( .I1(n9297), .O(n519) );
  NAND_GATE U671 ( .I1(n9366), .I2(n520), .O(n9369) );
  NOR_GATE U672 ( .I1(n9379), .I2(n9378), .O(n520) );
  AND3_GATE U673 ( .I1(n571), .I2(n10112), .I3(n10200), .O(n521) );
  NOR4_GATE U674 ( .I1(n219), .I2(n522), .I3(n209), .I4(n775), .O(n1390) );
  INV_GATE U675 ( .I1(n10987), .O(n522) );
  NAND_GATE U676 ( .I1(n7), .I2(n759), .O(n6195) );
  OR_GATE U677 ( .I1(n414), .I2(n4393), .O(n4662) );
  AND_GATE U678 ( .I1(n11867), .I2(n11871), .O(n523) );
  INV_GATE U679 ( .I1(n523), .O(n12267) );
  OR_GATE U680 ( .I1(n13103), .I2(n524), .O(n13104) );
  AND_GATE U681 ( .I1(n13102), .I2(n13101), .O(n524) );
  OR3_GATE U682 ( .I1(n1399), .I2(n525), .I3(n526), .O(n13932) );
  AND_GATE U683 ( .I1(n1406), .I2(A[31]), .O(n525) );
  AND_GATE U684 ( .I1(n13930), .I2(n13515), .O(n526) );
  NAND_GATE U685 ( .I1(n14290), .I2(n530), .O(n527) );
  NAND_GATE U686 ( .I1(n527), .I2(n528), .O(n539) );
  OR_GATE U687 ( .I1(n529), .I2(n14455), .O(n528) );
  INV_GATE U688 ( .I1(n14447), .O(n529) );
  AND_GATE U689 ( .I1(n14477), .I2(n14447), .O(n530) );
  NAND_GATE U690 ( .I1(n10602), .I2(n531), .O(n534) );
  NOR_GATE U691 ( .I1(n10600), .I2(n532), .O(n531) );
  INV_GATE U692 ( .I1(n11385), .O(n532) );
  NAND_GATE U693 ( .I1(n681), .I2(n535), .O(n533) );
  AND_GATE U694 ( .I1(n533), .I2(n534), .O(n11386) );
  AND_GATE U695 ( .I1(n10600), .I2(n11385), .O(n535) );
  NOR_GATE U696 ( .I1(n11777), .I2(n11774), .O(n580) );
  OR3_GATE U697 ( .I1(n536), .I2(n537), .I3(n11802), .O(n11805) );
  INV_GATE U698 ( .I1(n11800), .O(n536) );
  INV_GATE U699 ( .I1(n11799), .O(n537) );
  NOR_GATE U700 ( .I1(n13548), .I2(n13540), .O(n1023) );
  NAND_GATE U701 ( .I1(n14301), .I2(n14456), .O(n538) );
  NAND_GATE U702 ( .I1(n538), .I2(n539), .O(n14318) );
  NAND_GATE U703 ( .I1(n12749), .I2(n540), .O(n556) );
  NOR_GATE U704 ( .I1(n12750), .I2(n557), .O(n540) );
  AND_GATE U705 ( .I1(n541), .I2(n542), .O(n13576) );
  OR_GATE U706 ( .I1(n13550), .I2(n543), .O(n545) );
  NAND_GATE U707 ( .I1(n13553), .I2(n13555), .O(n543) );
  AND_GATE U708 ( .I1(n544), .I2(n545), .O(n13556) );
  OR_GATE U709 ( .I1(n546), .I2(n13956), .O(n13951) );
  NAND_GATE U710 ( .I1(n13557), .I2(n13556), .O(n546) );
  OR3_GATE U711 ( .I1(n547), .I2(n913), .I3(n12609), .O(n12615) );
  AND_GATE U712 ( .I1(n12608), .I2(n12611), .O(n547) );
  OR4_GATE U713 ( .I1(n11882), .I2(n548), .I3(n549), .I4(n11874), .O(n11878)
         );
  INV_GATE U714 ( .I1(n11876), .O(n548) );
  INV_GATE U715 ( .I1(n11875), .O(n549) );
  AND_GATE U716 ( .I1(n12689), .I2(n12688), .O(n550) );
  OR3_GATE U717 ( .I1(n550), .I2(n551), .I3(n12684), .O(n12686) );
  INV_GATE U718 ( .I1(n12682), .O(n551) );
  NAND_GATE U719 ( .I1(n14354), .I2(n554), .O(n552) );
  AND_GATE U720 ( .I1(n552), .I2(n553), .O(n14361) );
  OR_GATE U721 ( .I1(n978), .I2(n14356), .O(n553) );
  AND_GATE U722 ( .I1(n14355), .I2(n14357), .O(n554) );
  AND_GATE U723 ( .I1(n555), .I2(n556), .O(n12753) );
  INV_GATE U724 ( .I1(n12752), .O(n557) );
  AND_GATE U725 ( .I1(n558), .I2(n559), .O(n13149) );
  AND_GATE U726 ( .I1(n14317), .I2(n14316), .O(n560) );
  OR_GATE U727 ( .I1(n8876), .I2(n14813), .O(n8878) );
  OR_GATE U728 ( .I1(n9293), .I2(n14814), .O(n9295) );
  OR_GATE U729 ( .I1(n561), .I2(n11819), .O(n11830) );
  INV_GATE U730 ( .I1(n11826), .O(n561) );
  NAND_GATE U731 ( .I1(n11415), .I2(n564), .O(n562) );
  AND_GATE U732 ( .I1(n562), .I2(n563), .O(n11799) );
  OR_GATE U733 ( .I1(n11807), .I2(n11418), .O(n563) );
  AND_GATE U734 ( .I1(n11416), .I2(n11809), .O(n564) );
  NAND_GATE U735 ( .I1(n11808), .I2(n568), .O(n565) );
  AND_GATE U736 ( .I1(n565), .I2(n566), .O(n11815) );
  OR_GATE U737 ( .I1(n567), .I2(n11810), .O(n566) );
  INV_GATE U738 ( .I1(n11811), .O(n567) );
  AND_GATE U739 ( .I1(n11809), .I2(n11811), .O(n568) );
  NOR_GATE U740 ( .I1(n8876), .I2(n8883), .O(\A2[44] ) );
  AND_GATE U741 ( .I1(n10559), .I2(n10558), .O(n569) );
  NAND_GATE U742 ( .I1(n10114), .I2(n570), .O(n753) );
  NOR_GATE U743 ( .I1(n10113), .I2(n571), .O(n570) );
  INV_GATE U744 ( .I1(n10201), .O(n571) );
  NAND_GATE U745 ( .I1(n752), .I2(n753), .O(n572) );
  AND3_GATE U746 ( .I1(n13498), .I2(n13497), .I3(n13496), .O(n573) );
  OR3_GATE U747 ( .I1(n13943), .I2(n13942), .I3(n274), .O(n13945) );
  NAND_GATE U748 ( .I1(n8367), .I2(n576), .O(n574) );
  NAND_GATE U749 ( .I1(n574), .I2(n575), .O(n817) );
  OR_GATE U750 ( .I1(n8504), .I2(n8364), .O(n575) );
  AND_GATE U751 ( .I1(n8368), .I2(n8374), .O(n576) );
  AND_GATE U752 ( .I1(n11827), .I2(n11777), .O(n577) );
  NAND_GATE U753 ( .I1(n11778), .I2(n577), .O(n579) );
  NAND_GATE U754 ( .I1(n11776), .I2(n580), .O(n578) );
  AND_GATE U755 ( .I1(n578), .I2(n579), .O(n11779) );
  NAND_GATE U756 ( .I1(n8367), .I2(n583), .O(n581) );
  AND_GATE U757 ( .I1(n581), .I2(n582), .O(n8370) );
  AND_GATE U758 ( .I1(n8368), .I2(n8369), .O(n583) );
  NAND_GATE U759 ( .I1(n7186), .I2(n586), .O(n584) );
  AND_GATE U760 ( .I1(n584), .I2(n585), .O(n7189) );
  AND_GATE U761 ( .I1(n7187), .I2(n7188), .O(n586) );
  NAND_GATE U762 ( .I1(n7714), .I2(n589), .O(n587) );
  AND_GATE U763 ( .I1(n587), .I2(n588), .O(n7460) );
  OR_GATE U764 ( .I1(n309), .I2(n7710), .O(n588) );
  AND_GATE U765 ( .I1(n7708), .I2(n7716), .O(n589) );
  AND_GATE U766 ( .I1(n7702), .I2(n7701), .O(n590) );
  NAND_GATE U767 ( .I1(n8355), .I2(n593), .O(n591) );
  AND_GATE U768 ( .I1(n591), .I2(n592), .O(n8509) );
  OR_GATE U769 ( .I1(n8515), .I2(n8358), .O(n592) );
  AND_GATE U770 ( .I1(n8356), .I2(n8359), .O(n593) );
  AND3_GATE U771 ( .I1(n8510), .I2(n8509), .I3(n8360), .O(n594) );
  OR_GATE U772 ( .I1(n10571), .I2(n1323), .O(n10573) );
  NAND_GATE U773 ( .I1(n9253), .I2(n275), .O(n596) );
  NAND_GATE U774 ( .I1(n807), .I2(n276), .O(n595) );
  AND_GATE U775 ( .I1(n595), .I2(n596), .O(n9255) );
  AND_GATE U776 ( .I1(n9258), .I2(n9337), .O(n597) );
  OR3_GATE U777 ( .I1(n521), .I2(n10205), .I3(n572), .O(n10207) );
  AND_GATE U778 ( .I1(n9240), .I2(n9226), .O(n598) );
  NAND_GATE U779 ( .I1(n8861), .I2(n602), .O(n599) );
  NAND_GATE U780 ( .I1(n599), .I2(n600), .O(n608) );
  OR_GATE U781 ( .I1(n601), .I2(n9226), .O(n600) );
  INV_GATE U782 ( .I1(n9240), .O(n601) );
  AND_GATE U783 ( .I1(n9227), .I2(n9240), .O(n602) );
  AND3_GATE U784 ( .I1(n9355), .I2(n9356), .I3(n9232), .O(n603) );
  OR_GATE U785 ( .I1(n1320), .I2(n10976), .O(n10969) );
  AND_GATE U786 ( .I1(n13073), .I2(n13072), .O(n604) );
  AND_GATE U787 ( .I1(n8862), .I2(n598), .O(n605) );
  NAND_GATE U788 ( .I1(n9239), .I2(n605), .O(n607) );
  NAND_GATE U789 ( .I1(n9237), .I2(n608), .O(n606) );
  AND_GATE U790 ( .I1(n606), .I2(n607), .O(n9241) );
  AND_GATE U791 ( .I1(n10169), .I2(n609), .O(n612) );
  AND_GATE U792 ( .I1(n10168), .I2(n10580), .O(n609) );
  NAND_GATE U793 ( .I1(n10176), .I2(n612), .O(n610) );
  AND_GATE U794 ( .I1(n610), .I2(n611), .O(n10581) );
  OR_GATE U795 ( .I1(n10577), .I2(n926), .O(n611) );
  NOR_GATE U796 ( .I1(n13097), .I2(n604), .O(n613) );
  AND_GATE U797 ( .I1(n13932), .I2(n13931), .O(n614) );
  AND3_GATE U798 ( .I1(n13060), .I2(n13059), .I3(n13493), .O(n615) );
  INV_GATE U799 ( .I1(n615), .O(n13511) );
  OR_GATE U800 ( .I1(n9712), .I2(n14816), .O(n9714) );
  NAND_GATE U801 ( .I1(n10963), .I2(n618), .O(n616) );
  AND_GATE U802 ( .I1(n616), .I2(n617), .O(n10967) );
  AND_GATE U803 ( .I1(n10962), .I2(n10964), .O(n618) );
  AND_GATE U804 ( .I1(n9311), .I2(n9310), .O(n619) );
  AND_GATE U805 ( .I1(n752), .I2(n753), .O(n10202) );
  AND_GATE U806 ( .I1(n10113), .I2(n10201), .O(n620) );
  AND3_GATE U807 ( .I1(n10215), .I2(n10214), .I3(n10213), .O(n621) );
  OR3_GATE U808 ( .I1(n11790), .I2(n622), .I3(n623), .O(n11793) );
  AND_GATE U809 ( .I1(n11786), .I2(n911), .O(n622) );
  AND3_GATE U810 ( .I1(n11788), .I2(n11787), .I3(n911), .O(n623) );
  NAND_GATE U811 ( .I1(n14321), .I2(n627), .O(n624) );
  NAND_GATE U812 ( .I1(n624), .I2(n625), .O(n630) );
  OR_GATE U813 ( .I1(n626), .I2(n14422), .O(n625) );
  INV_GATE U814 ( .I1(n14392), .O(n626) );
  AND_GATE U815 ( .I1(n14440), .I2(n14392), .O(n627) );
  NAND_GATE U816 ( .I1(n14336), .I2(n630), .O(n628) );
  OR_GATE U817 ( .I1(n626), .I2(n14411), .O(n629) );
  OR_GATE U818 ( .I1(n11837), .I2(n411), .O(n11847) );
  OR_GATE U819 ( .I1(n626), .I2(n14398), .O(n631) );
  NAND_GATE U820 ( .I1(n14352), .I2(n14406), .O(n633) );
  INV_GATE U821 ( .I1(n633), .O(n936) );
  NAND3_GATE U822 ( .I1(n571), .I2(n10112), .I3(n10200), .O(n10203) );
  NAND3_GATE U823 ( .I1(n10101), .I2(n10105), .I3(n10219), .O(n10220) );
  NAND3_GATE U824 ( .I1(n11774), .I2(n11773), .I3(n11826), .O(n11820) );
  NAND3_GATE U825 ( .I1(n9576), .I2(n9577), .I3(n9583), .O(n9864) );
  AND_GATE U826 ( .I1(n6707), .I2(n6706), .O(n14802) );
  NAND4_GATE U827 ( .I1(n7159), .I2(n6742), .I3(n6746), .I4(n6743), .O(n7155)
         );
  AND3_GATE U828 ( .I1(n10942), .I2(n10943), .I3(n11030), .O(n11012) );
  AND_GATE U829 ( .I1(n6721), .I2(n6720), .O(n14804) );
  AND3_GATE U830 ( .I1(n6732), .I2(n6733), .I3(n6734), .O(n14805) );
  NAND_GATE U831 ( .I1(A[3]), .I2(B[30]), .O(n1850) );
  NAND3_GATE U832 ( .I1(n12622), .I2(n12621), .I3(n12693), .O(n12682) );
  AND_GATE U833 ( .I1(n10302), .I2(n10301), .O(n10885) );
  AND_GATE U834 ( .I1(n14576), .I2(n14276), .O(n14554) );
  AND_GATE U835 ( .I1(n10852), .I2(n10851), .O(n11297) );
  NAND3_GATE U836 ( .I1(n418), .I2(n13898), .I3(n13965), .O(n13900) );
  NAND5_GATE U837 ( .I1(n6925), .I2(n6216), .I3(n6215), .I4(n6513), .I5(n6217), 
        .O(n1360) );
  AND3_GATE U838 ( .I1(n8806), .I2(n8253), .I3(n8803), .O(n8617) );
  AND3_GATE U839 ( .I1(n12718), .I2(n12713), .I3(n12603), .O(n12703) );
  NAND4_GATE U840 ( .I1(n12606), .I2(n1261), .I3(n1260), .I4(n12605), .O(
        n12616) );
  NAND3_GATE U841 ( .I1(n8169), .I2(n8170), .I3(n8176), .O(n8663) );
  AND3_GATE U842 ( .I1(n13537), .I2(n13536), .I3(n13538), .O(n13939) );
  NAND4_GATE U843 ( .I1(n7223), .I2(n7095), .I3(n7230), .I4(n7096), .O(n7231)
         );
  AND_GATE U844 ( .I1(n13949), .I2(n13948), .O(n14830) );
  AND3_GATE U845 ( .I1(n11933), .I2(n11934), .I3(n11940), .O(n12585) );
  AND3_GATE U846 ( .I1(n12317), .I2(n12193), .I3(n12318), .O(n12582) );
  AND3_GATE U847 ( .I1(n12734), .I2(n12735), .I3(n12736), .O(n13455) );
  AND3_GATE U848 ( .I1(n13118), .I2(n13054), .I3(n13055), .O(n13472) );
  NAND3_GATE U849 ( .I1(n12290), .I2(n12291), .I3(n12597), .O(n13048) );
  NAND3_GATE U850 ( .I1(n9093), .I2(n9094), .I3(n9100), .O(n9494) );
  NAND3_GATE U851 ( .I1(n8717), .I2(n8718), .I3(n8724), .O(n9011) );
  NAND3_GATE U852 ( .I1(n6511), .I2(n6925), .I3(n6510), .O(n1361) );
  AND_GATE U853 ( .I1(n2006), .I2(n2007), .O(n2689) );
  NAND4_GATE U854 ( .I1(n13988), .I2(n13989), .I3(n13866), .I4(n13978), .O(
        n13982) );
  NAND3_GATE U855 ( .I1(n12564), .I2(n12565), .I3(n12571), .O(n12759) );
  AND3_GATE U856 ( .I1(n10627), .I2(n10543), .I3(n10628), .O(n10621) );
  NAND3_GATE U857 ( .I1(n11142), .I2(n11143), .I3(n11149), .O(n11524) );
  AND3_GATE U858 ( .I1(n11816), .I2(n11817), .I3(n11818), .O(n12640) );
  AND3_GATE U859 ( .I1(n11035), .I2(n11034), .I3(n11036), .O(n11778) );
  NAND5_GATE U860 ( .I1(n11774), .I2(n11035), .I3(n11777), .I4(n11034), .I5(
        n11036), .O(n11826) );
  AND_GATE U861 ( .I1(n1490), .I2(n1491), .O(n1819) );
  NAND_GATE U862 ( .I1(n9182), .I2(n9672), .O(n9442) );
  AND_GATE U863 ( .I1(n12237), .I2(n12238), .O(n14820) );
  NAND_GATE U864 ( .I1(n3625), .I2(n3626), .O(n3850) );
  AND3_GATE U865 ( .I1(n5129), .I2(n5130), .I3(n5131), .O(n5673) );
  AND_GATE U866 ( .I1(n8864), .I2(n9233), .O(n9252) );
  AND_GATE U867 ( .I1(n1823), .I2(n1824), .O(n2066) );
  AND_GATE U868 ( .I1(n1858), .I2(n1857), .O(n940) );
  NAND4_GATE U869 ( .I1(n13943), .I2(n13537), .I3(n13536), .I4(n13538), .O(
        n14372) );
  NAND3_GATE U870 ( .I1(n6019), .I2(n6020), .I3(n6033), .O(n6339) );
  NAND3_GATE U871 ( .I1(n11514), .I2(n11515), .I3(n11521), .O(n12000) );
  AND3_GATE U872 ( .I1(n13966), .I2(n13901), .I3(n13960), .O(n14325) );
  NAND3_GATE U873 ( .I1(n7967), .I2(n7231), .I3(n7232), .O(n7962) );
  NAND3_GATE U874 ( .I1(n6364), .I2(n6365), .I3(n6376), .O(n7083) );
  NAND3_GATE U875 ( .I1(n7410), .I2(n7952), .I3(n7964), .O(n7963) );
  NAND4_GATE U876 ( .I1(n10923), .I2(n10926), .I3(n10924), .I4(n10925), .O(
        n10929) );
  AND_GATE U877 ( .I1(n8862), .I2(n9226), .O(n9238) );
  AND_GATE U878 ( .I1(n8529), .I2(n8528), .O(n9217) );
  NAND3_GATE U879 ( .I1(n4471), .I2(n4753), .I3(n4762), .O(n4760) );
  NAND3_GATE U880 ( .I1(n5362), .I2(n5656), .I3(n5674), .O(n5670) );
  NAND3_GATE U881 ( .I1(n8532), .I2(n8533), .I3(n8539), .O(n8910) );
  AND_GATE U882 ( .I1(n14375), .I2(n14374), .O(n14826) );
  NAND3_GATE U883 ( .I1(n12352), .I2(n12353), .I3(n12359), .O(n12773) );
  NAND3_GATE U884 ( .I1(n11990), .I2(n11991), .I3(n11997), .O(n12362) );
  AND3_GATE U885 ( .I1(n8511), .I2(n8512), .I3(n8518), .O(n9237) );
  AND_GATE U886 ( .I1(n10586), .I2(n10587), .O(n10591) );
  AND_GATE U887 ( .I1(n6243), .I2(n6331), .O(n6313) );
  NAND3_GATE U888 ( .I1(n11082), .I2(n11083), .I3(n11089), .O(n11704) );
  AND3_GATE U889 ( .I1(n8765), .I2(n8231), .I3(n8774), .O(n8783) );
  AND3_GATE U890 ( .I1(n10496), .I2(n10010), .I3(n10501), .O(n10510) );
  AND3_GATE U891 ( .I1(n11437), .I2(n11739), .I3(n11438), .O(n1395) );
  NAND4_GATE U892 ( .I1(n12737), .I2(n12592), .I3(n12738), .I4(n13032), .O(
        n13030) );
  AND_GATE U893 ( .I1(n13448), .I2(n13895), .O(n13558) );
  AND_GATE U894 ( .I1(n13478), .I2(n13477), .O(n13544) );
  NAND3_GATE U895 ( .I1(n7706), .I2(n7707), .I3(n7720), .O(n8322) );
  AND3_GATE U896 ( .I1(n11439), .I2(n11366), .I3(n11435), .O(n11750) );
  NAND3_GATE U897 ( .I1(n13869), .I2(n13870), .I3(n13876), .O(n13978) );
  NAND3_GATE U898 ( .I1(n13420), .I2(n13421), .I3(n13427), .O(n13582) );
  NAND3_GATE U899 ( .I1(n13000), .I2(n13001), .I3(n13007), .O(n13165) );
  NAND3_GATE U900 ( .I1(n14293), .I2(n14294), .I3(n14300), .O(n14464) );
  NAND3_GATE U901 ( .I1(n9311), .I2(n9715), .I3(n9310), .O(n9717) );
  NAND4_GATE U902 ( .I1(n8447), .I2(n8448), .I3(n8879), .I4(n8454), .O(n8883)
         );
  AND3_GATE U903 ( .I1(n11351), .I2(n11352), .I3(n11447), .O(n11728) );
  AND3_GATE U904 ( .I1(n14291), .I2(n14292), .I3(n13880), .O(n14308) );
  NAND3_GATE U905 ( .I1(n13014), .I2(n13015), .I3(n13021), .O(n13154) );
  AND3_GATE U906 ( .I1(n6796), .I2(n6797), .I3(n6803), .O(n938) );
  NAND3_GATE U907 ( .I1(n2634), .I2(n2635), .I3(n2641), .O(n2999) );
  AND3_GATE U908 ( .I1(n4599), .I2(n4590), .I3(n4589), .O(n5343) );
  NAND3_GATE U909 ( .I1(n5345), .I2(n5342), .I3(n5456), .O(n5468) );
  AND_GATE U910 ( .I1(n12628), .I2(n13063), .O(n887) );
  NAND5_GATE U911 ( .I1(n634), .I2(n12281), .I3(n13100), .I4(n12280), .I5(
        n12282), .O(n13107) );
  INV_GATE U912 ( .I1(n13103), .O(n634) );
  AND3_GATE U913 ( .I1(n3752), .I2(n3754), .I3(n3753), .O(n4426) );
  NAND3_GATE U914 ( .I1(n6356), .I2(n6355), .I3(n6907), .O(n6914) );
  NAND4_GATE U915 ( .I1(n7433), .I2(n6886), .I3(n6884), .I4(n6885), .O(n7430)
         );
  AND_GATE U916 ( .I1(n13107), .I2(n13106), .O(n13112) );
  NAND3_GATE U917 ( .I1(n10359), .I2(n10360), .I3(n10366), .O(n10700) );
  AND_GATE U918 ( .I1(n13933), .I2(n13934), .O(n14823) );
  AND3_GATE U919 ( .I1(n6167), .I2(n6409), .I3(n6408), .O(n6946) );
  NAND4_GATE U920 ( .I1(n13551), .I2(n13129), .I3(n13124), .I4(n13130), .O(
        n13549) );
  AND3_GATE U921 ( .I1(n6353), .I2(n6352), .I3(n6354), .O(n6902) );
  AND3_GATE U922 ( .I1(n10484), .I2(n10485), .I3(n10491), .O(n779) );
  AND3_GATE U923 ( .I1(n6393), .I2(n6394), .I3(n6395), .O(n7070) );
  AND3_GATE U924 ( .I1(n8254), .I2(n7935), .I3(n8259), .O(n8268) );
  NAND3_GATE U925 ( .I1(n13545), .I2(n13549), .I3(n13465), .O(n13546) );
  NAND3_GATE U926 ( .I1(n635), .I2(n170), .I3(n9750), .O(n9747) );
  INV_GATE U927 ( .I1(n1284), .O(n635) );
  NAND3_GATE U928 ( .I1(n8866), .I2(n9247), .I3(n9264), .O(n9268) );
  AND_GATE U929 ( .I1(n1494), .I2(n1495), .O(n1796) );
  NAND3_GATE U930 ( .I1(n2769), .I2(n3102), .I3(n3120), .O(n3125) );
  NAND3_GATE U931 ( .I1(n3647), .I2(n3988), .I3(n4006), .O(n4011) );
  NAND3_GATE U932 ( .I1(n4508), .I2(n4917), .I3(n4935), .O(n4940) );
  NAND3_GATE U933 ( .I1(n5393), .I2(n5794), .I3(n5813), .O(n5818) );
  NAND3_GATE U934 ( .I1(n6686), .I2(n6290), .I3(n6279), .O(n6295) );
  NAND3_GATE U935 ( .I1(n8067), .I2(n7974), .I3(n8068), .O(n8051) );
  AND3_GATE U936 ( .I1(n9154), .I2(n8813), .I3(n9153), .O(n9167) );
  NAND3_GATE U937 ( .I1(n13904), .I2(n13556), .I3(n13557), .O(n13955) );
  NAND3_GATE U938 ( .I1(n13956), .I2(n13556), .I3(n13557), .O(n13905) );
  NAND3_GATE U939 ( .I1(n12319), .I2(n12320), .I3(n12326), .O(n12749) );
  NAND_GATE U940 ( .I1(n13556), .I2(n13557), .O(n13954) );
  NAND3_GATE U941 ( .I1(n10959), .I2(n10188), .I3(n10187), .O(n10956) );
  NAND3_GATE U942 ( .I1(n8841), .I2(n8840), .I3(n8846), .O(n8591) );
  NAND3_GATE U943 ( .I1(n9704), .I2(n9745), .I3(n10137), .O(n10134) );
  NAND3_GATE U944 ( .I1(n7132), .I2(n7475), .I3(n7491), .O(n7495) );
  NAND3_GATE U945 ( .I1(n5038), .I2(n5039), .I3(n5045), .O(n5797) );
  NAND3_GATE U946 ( .I1(n5048), .I2(n5049), .I3(n5055), .O(n5780) );
  NAND3_GATE U947 ( .I1(n6291), .I2(n6293), .I3(n6292), .O(n6712) );
  NAND3_GATE U948 ( .I1(n2547), .I2(n2548), .I3(n2554), .O(n3120) );
  NAND3_GATE U949 ( .I1(n5028), .I2(n5029), .I3(n5035), .O(n5813) );
  NAND3_GATE U950 ( .I1(n10255), .I2(n10084), .I3(n10253), .O(n10925) );
  AND_GATE U951 ( .I1(n12262), .I2(n12226), .O(n12652) );
  AND3_GATE U952 ( .I1(n12696), .I2(n12625), .I3(n12626), .O(n13101) );
  NAND4_GATE U953 ( .I1(n13506), .I2(n12698), .I3(n12699), .I4(n12700), .O(
        n13510) );
  NAND3_GATE U954 ( .I1(n13883), .I2(n13884), .I3(n13890), .O(n14307) );
  NAND3_GATE U955 ( .I1(n12739), .I2(n12740), .I3(n12746), .O(n13146) );
  NAND3_GATE U956 ( .I1(n13134), .I2(n13135), .I3(n13141), .O(n13894) );
  AND_GATE U957 ( .I1(n7104), .I2(n7430), .O(n7446) );
  AND3_GATE U958 ( .I1(n10270), .I2(n10271), .I3(n10272), .O(n10624) );
  NAND4_GATE U959 ( .I1(n1096), .I2(n12290), .I3(n12291), .I4(n12597), .O(
        n13044) );
  AND_GATE U960 ( .I1(n14547), .I2(n14280), .O(n14525) );
  AND3_GATE U961 ( .I1(n1993), .I2(n1994), .I3(n1995), .O(n897) );
  AND3_GATE U962 ( .I1(n3474), .I2(n3475), .I3(n3481), .O(n934) );
  AND3_GATE U963 ( .I1(n6050), .I2(n6049), .I3(n6051), .O(n6527) );
  NAND3_GATE U964 ( .I1(n7217), .I2(n7216), .I3(n7100), .O(n7424) );
  OR3_GATE U965 ( .I1(n7108), .I2(n747), .I3(n6543), .O(n7106) );
  NAND4_GATE U966 ( .I1(n14341), .I2(n13542), .I3(n13543), .I4(n13541), .O(
        n14345) );
  NAND3_GATE U967 ( .I1(n14368), .I2(n14367), .I3(n14366), .O(n14379) );
  NAND3_GATE U968 ( .I1(n9079), .I2(n9080), .I3(n9086), .O(n9508) );
  NAND3_GATE U969 ( .I1(n6548), .I2(n7118), .I3(n7117), .O(n6864) );
  AND3_GATE U970 ( .I1(n7752), .I2(n7751), .I3(n7753), .O(n8050) );
  NAND3_GATE U971 ( .I1(n5608), .I2(n5613), .I3(n6046), .O(n6036) );
  NAND3_GATE U972 ( .I1(n9961), .I2(n9962), .I3(n9968), .O(n10330) );
  NAND3_GATE U973 ( .I1(n9590), .I2(n9591), .I3(n9597), .O(n9850) );
  AND3_GATE U974 ( .I1(n9617), .I2(n9119), .I3(n9622), .O(n9477) );
  NAND3_GATE U975 ( .I1(n9947), .I2(n9948), .I3(n9954), .O(n10344) );
  AND3_GATE U976 ( .I1(n9331), .I2(n9332), .I3(n9333), .O(n9736) );
  NAND3_GATE U977 ( .I1(n9706), .I2(n10132), .I3(n9733), .O(n9738) );
  AND_GATE U978 ( .I1(B[29]), .I2(A[2]), .O(n2031) );
  AND3_GATE U979 ( .I1(n7651), .I2(n7652), .I3(n7658), .O(n857) );
  AND3_GATE U980 ( .I1(n7641), .I2(n7642), .I3(n7648), .O(n763) );
  NAND3_GATE U981 ( .I1(n11864), .I2(n11865), .I3(n12255), .O(n12256) );
  NAND3_GATE U982 ( .I1(n10815), .I2(n10816), .I3(n10822), .O(n11103) );
  NAND3_GATE U983 ( .I1(n10455), .I2(n10456), .I3(n10462), .O(n10675) );
  NAND3_GATE U984 ( .I1(n532), .I2(n10599), .I3(n11384), .O(n11392) );
  NAND3_GATE U985 ( .I1(n9604), .I2(n9605), .I3(n9612), .O(n9836) );
  NAND3_GATE U986 ( .I1(n7924), .I2(n7925), .I3(n7931), .O(n8089) );
  NAND3_GATE U987 ( .I1(n7958), .I2(n1357), .I3(n1358), .O(n8287) );
  NAND3_GATE U988 ( .I1(n9184), .I2(n9185), .I3(n9193), .O(n9194) );
  NAND3_GATE U989 ( .I1(n12283), .I2(n12287), .I3(n12719), .O(n12708) );
  AND_GATE U990 ( .I1(n2023), .I2(n2024), .O(n1225) );
  AND3_GATE U991 ( .I1(n5185), .I2(n5186), .I3(n5187), .O(n829) );
  NAND3_GATE U992 ( .I1(n11672), .I2(n11673), .I3(n11679), .O(n11953) );
  NAND3_GATE U993 ( .I1(n11271), .I2(n11272), .I3(n11278), .O(n11476) );
  AND_GATE U994 ( .I1(n11318), .I2(n11319), .O(n11457) );
  AND_GATE U995 ( .I1(n14518), .I2(n14284), .O(n14497) );
  NAND3_GATE U996 ( .I1(n3615), .I2(n3622), .I3(n3616), .O(n3836) );
  AND3_GATE U997 ( .I1(n7631), .I2(n7632), .I3(n7638), .O(n824) );
  AND3_GATE U998 ( .I1(n3429), .I2(n3430), .I3(n3436), .O(n822) );
  NAND3_GATE U999 ( .I1(n9369), .I2(n9370), .I3(n9382), .O(n10114) );
  AND3_GATE U1000 ( .I1(n7740), .I2(n7741), .I3(n7739), .O(n8041) );
  AND_GATE U1001 ( .I1(n8551), .I2(n8550), .O(n8918) );
  NAND3_GATE U1002 ( .I1(n4422), .I2(n4428), .I3(n4607), .O(n4605) );
  NAND3_GATE U1003 ( .I1(n6340), .I2(n6336), .I3(n6872), .O(n6879) );
  NAND3_GATE U1004 ( .I1(n10690), .I2(n10691), .I3(n10697), .O(n11128) );
  NAND3_GATE U1005 ( .I1(n10629), .I2(n10630), .I3(n10636), .O(n11357) );
  NAND3_GATE U1006 ( .I1(n10626), .I2(n10623), .I3(n10912), .O(n11058) );
  AND3_GATE U1007 ( .I1(n4315), .I2(n4316), .I3(n4317), .O(n903) );
  NOR_GATE U1008 ( .I1(n11881), .I2(n11880), .O(n12623) );
  AND3_GATE U1009 ( .I1(n8458), .I2(n8459), .I3(n8465), .O(n799) );
  AND3_GATE U1010 ( .I1(n8468), .I2(n8469), .I3(n8475), .O(n726) );
  NAND3_GATE U1011 ( .I1(n11118), .I2(n11119), .I3(n11125), .O(n11500) );
  NAND3_GATE U1012 ( .I1(n10919), .I2(n10918), .I3(n11040), .O(n11048) );
  NAND3_GATE U1013 ( .I1(n9451), .I2(n9452), .I3(n9458), .O(n10043) );
  NAND3_GATE U1014 ( .I1(n11490), .I2(n11491), .I3(n11497), .O(n11976) );
  OR_GATE U1015 ( .I1(B[30]), .I2(n1443), .O(n1400) );
  AND3_GATE U1016 ( .I1(n5920), .I2(n5921), .I3(n5927), .O(n750) );
  NAND3_GATE U1017 ( .I1(n8183), .I2(n8184), .I3(n8190), .O(n8649) );
  NAND3_GATE U1018 ( .I1(n11933), .I2(n11934), .I3(n11940), .O(n12583) );
  NAND3_GATE U1019 ( .I1(n11467), .I2(n11468), .I3(n11474), .O(n12182) );
  NAND3_GATE U1020 ( .I1(n11285), .I2(n11286), .I3(n11292), .O(n11683) );
  NAND3_GATE U1021 ( .I1(n11072), .I2(n11073), .I3(n11079), .O(n11729) );
  NAND3_GATE U1022 ( .I1(n8511), .I2(n8512), .I3(n8518), .O(n9239) );
  NOR_GATE U1023 ( .I1(n1275), .I2(n1158), .O(n636) );
  AND_GATE U1024 ( .I1(n13510), .I2(n13062), .O(n637) );
  AND_GATE U1025 ( .I1(n10651), .I2(n10650), .O(n638) );
  AND_GATE U1026 ( .I1(n14825), .I2(n14824), .O(n639) );
  AND_GATE U1027 ( .I1(n9163), .I2(n9162), .O(n640) );
  AND_GATE U1028 ( .I1(n13466), .I2(n13057), .O(n641) );
  AND_GATE U1029 ( .I1(n13501), .I2(n13500), .O(n642) );
  NAND_GATE U1030 ( .I1(n10032), .I2(n645), .O(n643) );
  AND_GATE U1031 ( .I1(n643), .I2(n644), .O(n10292) );
  OR_GATE U1032 ( .I1(n10300), .I2(n10036), .O(n644) );
  OR_GATE U1033 ( .I1(n13097), .I2(n604), .O(n13094) );
  OR_GATE U1034 ( .I1(n11860), .I2(n11859), .O(n11862) );
  AND_GATE U1035 ( .I1(n10071), .I2(n10067), .O(n646) );
  AND_GATE U1036 ( .I1(n11744), .I2(n11368), .O(n647) );
  INV_GATE U1037 ( .I1(n647), .O(n11423) );
  NAND_GATE U1038 ( .I1(n5740), .I2(n650), .O(n648) );
  AND_GATE U1039 ( .I1(n648), .I2(n649), .O(n5907) );
  OR_GATE U1040 ( .I1(n5913), .I2(n5743), .O(n649) );
  AND_GATE U1041 ( .I1(n5741), .I2(n5744), .O(n650) );
  NAND_GATE U1042 ( .I1(n6663), .I2(n653), .O(n651) );
  AND_GATE U1043 ( .I1(n651), .I2(n652), .O(n6761) );
  OR_GATE U1044 ( .I1(n6767), .I2(n6666), .O(n652) );
  AND_GATE U1045 ( .I1(n6664), .I2(n6667), .O(n653) );
  AND_GATE U1046 ( .I1(n9420), .I2(n9419), .O(n654) );
  NOR_GATE U1047 ( .I1(n1356), .I2(n1107), .O(n655) );
  AND_GATE U1048 ( .I1(n10477), .I2(n10476), .O(n656) );
  AND_GATE U1049 ( .I1(n9672), .I2(n9182), .O(n657) );
  AND_GATE U1050 ( .I1(n12220), .I2(n12219), .O(n658) );
  NAND_GATE U1051 ( .I1(n914), .I2(n659), .O(n12262) );
  AND_GATE U1052 ( .I1(n12255), .I2(n660), .O(n659) );
  INV_GATE U1053 ( .I1(n12258), .O(n660) );
  NAND_GATE U1054 ( .I1(n8644), .I2(n663), .O(n661) );
  AND_GATE U1055 ( .I1(n661), .I2(n662), .O(n9106) );
  OR_GATE U1056 ( .I1(n9111), .I2(n8647), .O(n662) );
  AND_GATE U1057 ( .I1(n8645), .I2(n8742), .O(n663) );
  AND_GATE U1058 ( .I1(n9480), .I2(n9117), .O(n664) );
  AND3_GATE U1059 ( .I1(n7118), .I2(n7117), .I3(n6548), .O(n665) );
  AND_GATE U1060 ( .I1(n6540), .I2(n6241), .O(n666) );
  INV_GATE U1061 ( .I1(n666), .O(n6332) );
  NAND_GATE U1062 ( .I1(n11692), .I2(n669), .O(n667) );
  AND_GATE U1063 ( .I1(n667), .I2(n668), .O(n11941) );
  OR_GATE U1064 ( .I1(n11947), .I2(n11694), .O(n668) );
  AND_GATE U1065 ( .I1(n11693), .I2(n11695), .O(n669) );
  NAND_GATE U1066 ( .I1(n12753), .I2(n672), .O(n670) );
  AND_GATE U1067 ( .I1(n670), .I2(n671), .O(n13432) );
  OR_GATE U1068 ( .I1(n13438), .I2(n12756), .O(n671) );
  AND_GATE U1069 ( .I1(n12754), .I2(n13024), .O(n672) );
  NAND_GATE U1070 ( .I1(n13620), .I2(n675), .O(n673) );
  AND_GATE U1071 ( .I1(n673), .I2(n674), .O(n14040) );
  OR_GATE U1072 ( .I1(n14046), .I2(n13623), .O(n674) );
  AND_GATE U1073 ( .I1(n13621), .I2(n13835), .O(n675) );
  AND_GATE U1074 ( .I1(n5262), .I2(n5263), .O(n676) );
  AND3_GATE U1075 ( .I1(n10232), .I2(n10231), .I3(n10230), .O(n677) );
  AND_GATE U1076 ( .I1(n10098), .I2(n10097), .O(n678) );
  AND_GATE U1077 ( .I1(n9134), .I2(n9133), .O(n679) );
  AND_GATE U1078 ( .I1(n4717), .I2(n4716), .O(n680) );
  AND3_GATE U1079 ( .I1(n10553), .I2(n10552), .I3(n10551), .O(n681) );
  NAND_GATE U1080 ( .I1(n14321), .I2(n14440), .O(n683) );
  AND3_GATE U1081 ( .I1(n13905), .I2(n13953), .I3(n13955), .O(n684) );
  NAND_GATE U1082 ( .I1(n10312), .I2(n687), .O(n685) );
  AND_GATE U1083 ( .I1(n685), .I2(n686), .O(n10843) );
  OR_GATE U1084 ( .I1(n10848), .I2(n10315), .O(n686) );
  AND_GATE U1085 ( .I1(n10313), .I2(n10494), .O(n687) );
  NAND_GATE U1086 ( .I1(n6475), .I2(n688), .O(n6966) );
  NOR_GATE U1087 ( .I1(n689), .I2(n1364), .O(n688) );
  INV_GATE U1088 ( .I1(n6474), .O(n689) );
  AND3_GATE U1089 ( .I1(n9122), .I2(n8763), .I3(n9121), .O(n690) );
  NAND_GATE U1090 ( .I1(n7323), .I2(n693), .O(n691) );
  AND_GATE U1091 ( .I1(n691), .I2(n692), .O(n7852) );
  OR_GATE U1092 ( .I1(n7858), .I2(n7326), .O(n692) );
  AND_GATE U1093 ( .I1(n7324), .I2(n7327), .O(n693) );
  AND_GATE U1094 ( .I1(n6491), .I2(n6490), .O(n694) );
  AND_GATE U1095 ( .I1(n10883), .I2(n10523), .O(n695) );
  AND_GATE U1096 ( .I1(n7304), .I2(n7303), .O(n696) );
  NAND_GATE U1097 ( .I1(n3888), .I2(n699), .O(n697) );
  AND_GATE U1098 ( .I1(n697), .I2(n698), .O(n4297) );
  OR_GATE U1099 ( .I1(n4303), .I2(n3891), .O(n698) );
  AND_GATE U1100 ( .I1(n3889), .I2(n3892), .O(n699) );
  AND3_GATE U1101 ( .I1(n6249), .I2(n6248), .I3(n5683), .O(n700) );
  AND_GATE U1102 ( .I1(n7691), .I2(n7690), .O(n701) );
  AND_GATE U1103 ( .I1(n3730), .I2(n3612), .O(n702) );
  AND3_GATE U1104 ( .I1(n6857), .I2(n6856), .I3(n6855), .O(n703) );
  AND3_GATE U1105 ( .I1(n5162), .I2(n5161), .I3(n4759), .O(n704) );
  AND_GATE U1106 ( .I1(n8317), .I2(n8316), .O(n705) );
  AND_GATE U1107 ( .I1(n6052), .I2(n5607), .O(n706) );
  NAND_GATE U1108 ( .I1(n4845), .I2(n709), .O(n707) );
  AND_GATE U1109 ( .I1(n707), .I2(n708), .O(n5089) );
  OR_GATE U1110 ( .I1(n5095), .I2(n4848), .O(n708) );
  AND_GATE U1111 ( .I1(n4846), .I2(n4849), .O(n709) );
  NAND_GATE U1112 ( .I1(n3903), .I2(n712), .O(n710) );
  AND_GATE U1113 ( .I1(n710), .I2(n711), .O(n4286) );
  OR_GATE U1114 ( .I1(n4292), .I2(n3906), .O(n711) );
  AND_GATE U1115 ( .I1(n3904), .I2(n3907), .O(n712) );
  AND_GATE U1116 ( .I1(n5917), .I2(n5916), .O(n713) );
  INV_GATE U1117 ( .I1(n713), .O(n6640) );
  AND_GATE U1118 ( .I1(n7427), .I2(n7426), .O(n714) );
  AND3_GATE U1119 ( .I1(n11400), .I2(n11399), .I3(n11398), .O(n715) );
  AND3_GATE U1120 ( .I1(n11834), .I2(n11833), .I3(n11832), .O(n716) );
  AND3_GATE U1121 ( .I1(n9400), .I2(n9399), .I3(n9398), .O(n717) );
  AND3_GATE U1122 ( .I1(n9438), .I2(n9437), .I3(n9436), .O(n718) );
  AND_GATE U1123 ( .I1(n10177), .I2(n10176), .O(n719) );
  NAND_GATE U1124 ( .I1(n6633), .I2(n722), .O(n720) );
  AND_GATE U1125 ( .I1(n720), .I2(n721), .O(n6783) );
  OR_GATE U1126 ( .I1(n6789), .I2(n6635), .O(n721) );
  AND_GATE U1127 ( .I1(n6634), .I2(n6636), .O(n722) );
  AND3_GATE U1128 ( .I1(n4276), .I2(n4275), .I3(n3924), .O(n723) );
  NAND_GATE U1129 ( .I1(n1444), .I2(A[1]), .O(n724) );
  OR_GATE U1130 ( .I1(n12762), .I2(n12761), .O(n12764) );
  OR_GATE U1131 ( .I1(n1444), .I2(A[1]), .O(n14241) );
  NAND_GATE U1132 ( .I1(n7003), .I2(n725), .O(n769) );
  AND_GATE U1133 ( .I1(n7001), .I2(n7000), .O(n725) );
  INV_GATE U1134 ( .I1(n726), .O(n8897) );
  OR_GATE U1135 ( .I1(n13103), .I2(n13102), .O(n13063) );
  AND3_GATE U1136 ( .I1(n13116), .I2(n13115), .I3(n13114), .O(n727) );
  OR3_GATE U1137 ( .I1(n5298), .I2(n728), .I3(n4688), .O(n5301) );
  INV_GATE U1138 ( .I1(n4689), .O(n728) );
  NOR3_GATE U1139 ( .I1(n5593), .I2(n6207), .I3(n5592), .O(n729) );
  OR_GATE U1140 ( .I1(n713), .I2(n6642), .O(n6644) );
  AND_GATE U1141 ( .I1(n4738), .I2(n4735), .O(n730) );
  INV_GATE U1142 ( .I1(n730), .O(n4740) );
  AND3_GATE U1143 ( .I1(n3611), .I2(n3610), .I3(n3734), .O(n731) );
  NAND_GATE U1144 ( .I1(n8333), .I2(n734), .O(n732) );
  AND_GATE U1145 ( .I1(n732), .I2(n733), .O(n8337) );
  OR_GATE U1146 ( .I1(n8332), .I2(n8335), .O(n733) );
  AND_GATE U1147 ( .I1(n8334), .I2(n8336), .O(n734) );
  NAND_GATE U1148 ( .I1(n6017), .I2(n735), .O(n6020) );
  NOR_GATE U1149 ( .I1(n6030), .I2(n6029), .O(n735) );
  NAND_GATE U1150 ( .I1(n7714), .I2(n738), .O(n736) );
  AND_GATE U1151 ( .I1(n736), .I2(n737), .O(n7705) );
  OR_GATE U1152 ( .I1(n7717), .I2(n7710), .O(n737) );
  AND_GATE U1153 ( .I1(n7708), .I2(n7459), .O(n738) );
  NAND_GATE U1154 ( .I1(n7112), .I2(n741), .O(n739) );
  AND_GATE U1155 ( .I1(n739), .I2(n740), .O(n7117) );
  OR_GATE U1156 ( .I1(n7115), .I2(n7106), .O(n740) );
  AND_GATE U1157 ( .I1(n7105), .I2(n6547), .O(n741) );
  AND3_GATE U1158 ( .I1(n9354), .I2(n9353), .I3(n9352), .O(n742) );
  AND_GATE U1159 ( .I1(n4728), .I2(n4724), .O(n743) );
  OR_GATE U1160 ( .I1(n3741), .I2(n3819), .O(n744) );
  AND_GATE U1161 ( .I1(n3588), .I2(n3587), .O(n745) );
  AND_GATE U1162 ( .I1(n4348), .I2(n3813), .O(n746) );
  INV_GATE U1163 ( .I1(n746), .O(n4351) );
  OR_GATE U1164 ( .I1(n3810), .I2(n929), .O(n3812) );
  AND_GATE U1165 ( .I1(n6239), .I2(n6238), .O(n747) );
  INV_GATE U1166 ( .I1(n747), .O(n6542) );
  AND3_GATE U1167 ( .I1(n12216), .I2(n12215), .I3(n12609), .O(n748) );
  OR_GATE U1168 ( .I1(B[18]), .I2(n1444), .O(n6988) );
  AND_GATE U1169 ( .I1(n9983), .I2(n9982), .O(n749) );
  INV_GATE U1170 ( .I1(n749), .O(n10317) );
  INV_GATE U1171 ( .I1(n750), .O(n6626) );
  AND3_GATE U1172 ( .I1(n11268), .I2(n11489), .I3(n11488), .O(n751) );
  INV_GATE U1173 ( .I1(n751), .O(n11479) );
  NAND_GATE U1174 ( .I1(n359), .I2(n620), .O(n752) );
  AND_GATE U1175 ( .I1(n752), .I2(n753), .O(n10115) );
  AND3_GATE U1176 ( .I1(n10955), .I2(n10954), .I3(n10953), .O(n754) );
  OR_GATE U1177 ( .I1(n1390), .I2(n755), .O(n11796) );
  AND_GATE U1178 ( .I1(n11414), .I2(n775), .O(n755) );
  AND_GATE U1179 ( .I1(n11743), .I2(n11742), .O(n756) );
  AND_GATE U1180 ( .I1(n6937), .I2(n6936), .O(n757) );
  NAND_GATE U1181 ( .I1(n5286), .I2(n4686), .O(n758) );
  AND_GATE U1182 ( .I1(n5512), .I2(n5511), .O(n759) );
  AND_GATE U1183 ( .I1(n4403), .I2(n4408), .O(n760) );
  INV_GATE U1184 ( .I1(n760), .O(n4618) );
  AND3_GATE U1185 ( .I1(n7937), .I2(n7408), .I3(n7936), .O(n761) );
  INV_GATE U1186 ( .I1(n761), .O(n7956) );
  AND3_GATE U1187 ( .I1(n9139), .I2(n8795), .I3(n9145), .O(n762) );
  INV_GATE U1188 ( .I1(n762), .O(n8961) );
  OR_GATE U1189 ( .I1(n10320), .I2(n749), .O(n10322) );
  OR_GATE U1190 ( .I1(n11093), .I2(n11095), .O(n10838) );
  OR_GATE U1191 ( .I1(n10595), .I2(n569), .O(n10594) );
  AND_GATE U1192 ( .I1(n5286), .I2(n4686), .O(n764) );
  OR_GATE U1193 ( .I1(n6203), .I2(n729), .O(n6209) );
  AND_GATE U1194 ( .I1(n6192), .I2(n5590), .O(n765) );
  INV_GATE U1195 ( .I1(n765), .O(n6211) );
  AND_GATE U1196 ( .I1(n766), .I2(n767), .O(n14330) );
  NAND_GATE U1197 ( .I1(n6998), .I2(n770), .O(n768) );
  AND_GATE U1198 ( .I1(n768), .I2(n769), .O(n7004) );
  AND_GATE U1199 ( .I1(n6997), .I2(n7003), .O(n770) );
  AND3_GATE U1200 ( .I1(n11669), .I2(n11964), .I3(n11963), .O(n771) );
  NAND_GATE U1201 ( .I1(n11484), .I2(n774), .O(n772) );
  AND_GATE U1202 ( .I1(n772), .I2(n773), .O(n11964) );
  OR_GATE U1203 ( .I1(n11969), .I2(n11487), .O(n773) );
  AND_GATE U1204 ( .I1(n11485), .I2(n11668), .O(n774) );
  NOR3_GATE U1205 ( .I1(n928), .I2(n776), .I3(n777), .O(n775) );
  AND_GATE U1206 ( .I1(n357), .I2(n11410), .O(n776) );
  AND_GATE U1207 ( .I1(n1414), .I2(A[31]), .O(n777) );
  OR_GATE U1208 ( .I1(n6325), .I2(n666), .O(n6326) );
  AND3_GATE U1209 ( .I1(n10483), .I2(n9987), .I3(n10482), .O(n778) );
  INV_GATE U1210 ( .I1(n778), .O(n10306) );
  OR_GATE U1211 ( .I1(n10655), .I2(n779), .O(n10657) );
  NOR_GATE U1212 ( .I1(n9204), .I2(n9205), .O(n780) );
  INV_GATE U1213 ( .I1(n780), .O(n9406) );
  AND3_GATE U1214 ( .I1(n11018), .I2(n11017), .I3(n11016), .O(n781) );
  AND_GATE U1215 ( .I1(n5354), .I2(n5353), .O(n782) );
  OR_GATE U1216 ( .I1(n10201), .I2(n10114), .O(n10111) );
  AND_GATE U1217 ( .I1(n6535), .I2(n6534), .O(n783) );
  AND_GATE U1218 ( .I1(n7453), .I2(n7124), .O(n784) );
  INV_GATE U1219 ( .I1(n784), .O(n7199) );
  AND_GATE U1220 ( .I1(n785), .I2(n786), .O(n13457) );
  NAND_GATE U1221 ( .I1(n11098), .I2(n790), .O(n787) );
  AND_GATE U1222 ( .I1(n787), .I2(n788), .O(n11674) );
  OR_GATE U1223 ( .I1(n789), .I2(n11100), .O(n788) );
  INV_GATE U1224 ( .I1(n11101), .O(n789) );
  AND_GATE U1225 ( .I1(n11099), .I2(n11101), .O(n790) );
  OR_GATE U1226 ( .I1(n6448), .I2(n6447), .O(n6450) );
  AND_GATE U1227 ( .I1(n14282), .I2(n14531), .O(n791) );
  INV_GATE U1228 ( .I1(n791), .O(n14509) );
  OR_GATE U1229 ( .I1(n778), .I2(n10307), .O(n10309) );
  AND3_GATE U1230 ( .I1(n6977), .I2(n6458), .I3(n6976), .O(n792) );
  INV_GATE U1231 ( .I1(n792), .O(n7016) );
  AND3_GATE U1232 ( .I1(n7258), .I2(n7257), .I3(n7256), .O(n793) );
  OR_GATE U1233 ( .I1(n7014), .I2(n792), .O(n7018) );
  AND3_GATE U1234 ( .I1(n13959), .I2(n13958), .I3(n13957), .O(n794) );
  INV_GATE U1235 ( .I1(n794), .O(n14419) );
  AND_GATE U1236 ( .I1(n8632), .I2(n8628), .O(n795) );
  INV_GATE U1237 ( .I1(n795), .O(n8759) );
  AND3_GATE U1238 ( .I1(n6204), .I2(n5600), .I3(n5599), .O(n796) );
  AND_GATE U1239 ( .I1(n5939), .I2(n5938), .O(n797) );
  INV_GATE U1240 ( .I1(n797), .O(n6611) );
  AND_GATE U1241 ( .I1(n5110), .I2(n5109), .O(n798) );
  INV_GATE U1242 ( .I1(n798), .O(n5437) );
  INV_GATE U1243 ( .I1(n799), .O(n8886) );
  AND_GATE U1244 ( .I1(n5099), .I2(n5098), .O(n800) );
  AND_GATE U1245 ( .I1(n4274), .I2(n4273), .O(n801) );
  INV_GATE U1246 ( .I1(n801), .O(n4822) );
  AND3_GATE U1247 ( .I1(n8753), .I2(n8752), .I3(n8751), .O(n802) );
  INV_GATE U1248 ( .I1(n802), .O(n8993) );
  NAND_GATE U1249 ( .I1(n5172), .I2(n805), .O(n803) );
  AND_GATE U1250 ( .I1(n803), .I2(n804), .O(n5355) );
  OR_GATE U1251 ( .I1(n782), .I2(n5998), .O(n804) );
  AND_GATE U1252 ( .I1(n5171), .I2(n5622), .O(n805) );
  AND_GATE U1253 ( .I1(n9344), .I2(n9343), .O(n806) );
  AND_GATE U1254 ( .I1(n8508), .I2(n8507), .O(n807) );
  NAND_GATE U1255 ( .I1(n6847), .I2(n6846), .O(n808) );
  AND_GATE U1256 ( .I1(n7463), .I2(n7130), .O(n809) );
  AND3_GATE U1257 ( .I1(n4337), .I2(n4336), .I3(n4335), .O(n810) );
  NAND_GATE U1258 ( .I1(n3853), .I2(n3852), .O(n811) );
  AND3_GATE U1259 ( .I1(n2683), .I2(n2682), .I3(n2681), .O(n812) );
  AND_GATE U1260 ( .I1(n1996), .I2(n1874), .O(n813) );
  AND_GATE U1261 ( .I1(n9258), .I2(n9257), .O(n814) );
  NAND_GATE U1262 ( .I1(n8370), .I2(n817), .O(n815) );
  AND_GATE U1263 ( .I1(n815), .I2(n816), .O(n8498) );
  OR_GATE U1264 ( .I1(n8504), .I2(n8373), .O(n816) );
  NAND_GATE U1265 ( .I1(n4751), .I2(n820), .O(n818) );
  AND_GATE U1266 ( .I1(n818), .I2(n819), .O(n5161) );
  OR_GATE U1267 ( .I1(n5170), .I2(n4756), .O(n819) );
  AND_GATE U1268 ( .I1(n4752), .I2(n4758), .O(n820) );
  AND_GATE U1269 ( .I1(n3623), .I2(n3622), .O(n821) );
  INV_GATE U1270 ( .I1(n822), .O(n3943) );
  AND_GATE U1271 ( .I1(n2609), .I2(n2608), .O(n823) );
  INV_GATE U1272 ( .I1(n823), .O(n3041) );
  INV_GATE U1273 ( .I1(n824), .O(n8422) );
  AND_GATE U1274 ( .I1(n6847), .I2(n6846), .O(n825) );
  OR_GATE U1275 ( .I1(n8650), .I2(n8649), .O(n8654) );
  AND3_GATE U1276 ( .I1(n9603), .I2(n9104), .I3(n9602), .O(n826) );
  INV_GATE U1277 ( .I1(n826), .O(n9484) );
  OR_GATE U1278 ( .I1(n825), .I2(n7467), .O(n7465) );
  AND_GATE U1279 ( .I1(n6553), .I2(n6247), .O(n827) );
  NAND_GATE U1280 ( .I1(n1858), .I2(n1857), .O(n828) );
  OR_GATE U1281 ( .I1(n11789), .I2(n911), .O(n11792) );
  OR_GATE U1282 ( .I1(n829), .I2(n5450), .O(n5453) );
  AND_GATE U1283 ( .I1(n10151), .I2(n10147), .O(n830) );
  AND_GATE U1284 ( .I1(n8486), .I2(n8485), .O(n831) );
  AND_GATE U1285 ( .I1(n7669), .I2(n7668), .O(n832) );
  AND_GATE U1286 ( .I1(n6825), .I2(n6824), .O(n833) );
  AND_GATE U1287 ( .I1(n5961), .I2(n5960), .O(n834) );
  AND_GATE U1288 ( .I1(n5121), .I2(n5120), .O(n836) );
  AND_GATE U1289 ( .I1(n3471), .I2(n3470), .O(n837) );
  AND_GATE U1290 ( .I1(n2992), .I2(n2755), .O(n838) );
  AND_GATE U1291 ( .I1(n1990), .I2(n1876), .O(n839) );
  AND_GATE U1292 ( .I1(n2056), .I2(n2055), .O(n840) );
  NAND_GATE U1293 ( .I1(n8400), .I2(n843), .O(n841) );
  AND_GATE U1294 ( .I1(n841), .I2(n842), .O(n8476) );
  OR_GATE U1295 ( .I1(n8482), .I2(n8403), .O(n842) );
  AND_GATE U1296 ( .I1(n8401), .I2(n8404), .O(n843) );
  NAND_GATE U1297 ( .I1(n7498), .I2(n846), .O(n844) );
  AND_GATE U1298 ( .I1(n844), .I2(n845), .O(n7659) );
  OR_GATE U1299 ( .I1(n7665), .I2(n7501), .O(n845) );
  AND_GATE U1300 ( .I1(n7499), .I2(n7502), .O(n846) );
  OR_GATE U1301 ( .I1(n6821), .I2(n6591), .O(n847) );
  NAND_GATE U1302 ( .I1(n5693), .I2(n850), .O(n848) );
  AND_GATE U1303 ( .I1(n848), .I2(n849), .O(n5951) );
  OR_GATE U1304 ( .I1(n5957), .I2(n5696), .O(n849) );
  AND_GATE U1305 ( .I1(n5694), .I2(n5697), .O(n850) );
  NAND_GATE U1306 ( .I1(n4814), .I2(n853), .O(n851) );
  AND_GATE U1307 ( .I1(n851), .I2(n852), .O(n5111) );
  OR_GATE U1308 ( .I1(n5117), .I2(n4817), .O(n852) );
  AND_GATE U1309 ( .I1(n4815), .I2(n4818), .O(n853) );
  NAND_GATE U1310 ( .I1(n3017), .I2(n856), .O(n854) );
  AND_GATE U1311 ( .I1(n854), .I2(n855), .O(n3461) );
  OR_GATE U1312 ( .I1(n3467), .I2(n3020), .O(n855) );
  AND_GATE U1313 ( .I1(n3018), .I2(n3021), .O(n856) );
  INV_GATE U1314 ( .I1(n857), .O(n8393) );
  AND_GATE U1315 ( .I1(n9262), .I2(n8868), .O(n858) );
  INV_GATE U1316 ( .I1(n858), .O(n9280) );
  OR_GATE U1317 ( .I1(n8492), .I2(n1336), .O(n8495) );
  AND_GATE U1318 ( .I1(n859), .I2(n860), .O(n10900) );
  NAND_GATE U1319 ( .I1(n640), .I2(n863), .O(n861) );
  AND_GATE U1320 ( .I1(n861), .I2(n862), .O(n9665) );
  OR_GATE U1321 ( .I1(n9664), .I2(n9663), .O(n862) );
  AND_GATE U1322 ( .I1(n9659), .I2(n9797), .O(n863) );
  NAND_GATE U1323 ( .I1(n7372), .I2(n866), .O(n864) );
  AND_GATE U1324 ( .I1(n864), .I2(n865), .O(n7375) );
  OR_GATE U1325 ( .I1(n7368), .I2(n7374), .O(n865) );
  AND_GATE U1326 ( .I1(n7371), .I2(n7900), .O(n866) );
  AND_GATE U1327 ( .I1(n6136), .I2(n5575), .O(n867) );
  AND_GATE U1328 ( .I1(n13094), .I2(n13098), .O(n868) );
  AND3_GATE U1329 ( .I1(n12649), .I2(n12651), .I3(n12650), .O(n869) );
  NAND_GATE U1330 ( .I1(n8060), .I2(n872), .O(n870) );
  AND_GATE U1331 ( .I1(n870), .I2(n871), .O(n8068) );
  OR_GATE U1332 ( .I1(n8063), .I2(n8057), .O(n871) );
  AND_GATE U1333 ( .I1(n8056), .I2(n7973), .O(n872) );
  NOR_GATE U1334 ( .I1(n869), .I2(n12648), .O(n873) );
  AND3_GATE U1335 ( .I1(n9773), .I2(n9772), .I3(n9771), .O(n874) );
  AND_GATE U1336 ( .I1(n8937), .I2(n8936), .O(n875) );
  AND3_GATE U1337 ( .I1(n8072), .I2(n8071), .I3(n8070), .O(n876) );
  AND3_GATE U1338 ( .I1(n7220), .I2(n7219), .I3(n277), .O(n877) );
  AND3_GATE U1339 ( .I1(n6078), .I2(n6077), .I3(n6076), .O(n878) );
  AND_GATE U1340 ( .I1(n6231), .I2(n6230), .O(n879) );
  AND3_GATE U1341 ( .I1(n5213), .I2(n5212), .I3(n5211), .O(n880) );
  AND3_GATE U1342 ( .I1(n5327), .I2(n5326), .I3(n5329), .O(n881) );
  AND_GATE U1343 ( .I1(n3798), .I2(n3799), .O(n882) );
  AND_GATE U1344 ( .I1(n3572), .I2(n3571), .O(n883) );
  AND3_GATE U1345 ( .I1(n10548), .I2(n10547), .I3(n10616), .O(n884) );
  AND3_GATE U1346 ( .I1(n11054), .I2(n11053), .I3(n11052), .O(n885) );
  AND3_GATE U1347 ( .I1(n9805), .I2(n9668), .I3(n9793), .O(n886) );
  INV_GATE U1348 ( .I1(n886), .O(n10050) );
  OR_GATE U1349 ( .I1(n887), .I2(n12673), .O(n12675) );
  OR_GATE U1350 ( .I1(n11848), .I2(n11859), .O(n11865) );
  OR3_GATE U1351 ( .I1(n12677), .I2(n887), .I3(n12673), .O(n12672) );
  OR_GATE U1352 ( .I1(n888), .I2(n8267), .O(n8270) );
  INV_GATE U1353 ( .I1(n8269), .O(n888) );
  NAND_GATE U1354 ( .I1(n7480), .I2(n891), .O(n889) );
  AND_GATE U1355 ( .I1(n889), .I2(n890), .O(n7483) );
  OR_GATE U1356 ( .I1(n7478), .I2(n7477), .O(n890) );
  AND_GATE U1357 ( .I1(n7479), .I2(n7482), .O(n891) );
  NAND_GATE U1358 ( .I1(n892), .I2(n6830), .O(n6829) );
  NOR_GATE U1359 ( .I1(n6832), .I2(n6831), .O(n892) );
  NAND3_GATE U1360 ( .I1(n5146), .I2(n5145), .I3(n4776), .O(n893) );
  NAND_GATE U1361 ( .I1(n3849), .I2(n3628), .O(n894) );
  NOR_GATE U1362 ( .I1(n1255), .I2(n1224), .O(n895) );
  AND_GATE U1363 ( .I1(n2740), .I2(n2038), .O(n896) );
  OR_GATE U1364 ( .I1(n897), .I2(n2680), .O(n2675) );
  NAND_GATE U1365 ( .I1(n903), .I2(n900), .O(n898) );
  AND_GATE U1366 ( .I1(n898), .I2(n899), .O(n4574) );
  OR_GATE U1367 ( .I1(n4572), .I2(n4571), .O(n899) );
  AND_GATE U1368 ( .I1(n8497), .I2(n8496), .O(n901) );
  AND_GATE U1369 ( .I1(n3492), .I2(n3491), .O(n902) );
  OR_GATE U1370 ( .I1(n826), .I2(n9481), .O(n9485) );
  OR_GATE U1371 ( .I1(n903), .I2(n4576), .O(n4571) );
  NAND_GATE U1372 ( .I1(n904), .I2(n6841), .O(n6840) );
  NOR_GATE U1373 ( .I1(n6843), .I2(n6842), .O(n904) );
  AND_GATE U1374 ( .I1(n4328), .I2(n4327), .O(n905) );
  AND_GATE U1375 ( .I1(n2879), .I2(n2878), .O(n906) );
  AND_GATE U1376 ( .I1(n2018), .I2(n2017), .O(n907) );
  OR_GATE U1377 ( .I1(n4331), .I2(n1266), .O(n4333) );
  AND_GATE U1378 ( .I1(n5668), .I2(n5364), .O(n908) );
  INV_GATE U1379 ( .I1(n908), .O(n5688) );
  AND3_GATE U1380 ( .I1(n5156), .I2(n5155), .I3(n4774), .O(n909) );
  INV_GATE U1381 ( .I1(n909), .O(n5147) );
  OR_GATE U1382 ( .I1(n798), .I2(n5439), .O(n5441) );
  AND_GATE U1383 ( .I1(n6814), .I2(n6813), .O(n910) );
  INV_GATE U1384 ( .I1(n910), .O(n7506) );
  OR_GATE U1385 ( .I1(n810), .I2(n4754), .O(n4748) );
  OR_GATE U1386 ( .I1(n613), .I2(n13093), .O(n13095) );
  AND_GATE U1387 ( .I1(n11409), .I2(n11408), .O(n911) );
  NOR_GATE U1388 ( .I1(n12258), .I2(n12256), .O(n912) );
  OR_GATE U1389 ( .I1(n12608), .I2(n913), .O(n12613) );
  INV_GATE U1390 ( .I1(n12610), .O(n913) );
  INV_GATE U1391 ( .I1(n11866), .O(n914) );
  AND_GATE U1392 ( .I1(n2907), .I2(n2908), .O(n915) );
  NAND_GATE U1393 ( .I1(n916), .I2(n9359), .O(n9357) );
  NOR_GATE U1394 ( .I1(n9363), .I2(n9360), .O(n916) );
  NAND_GATE U1395 ( .I1(n917), .I2(n8523), .O(n8522) );
  NOR_GATE U1396 ( .I1(n8527), .I2(n8524), .O(n917) );
  NAND_GATE U1397 ( .I1(n7696), .I2(n918), .O(n7694) );
  NOR_GATE U1398 ( .I1(n7700), .I2(n7697), .O(n918) );
  AND_GATE U1399 ( .I1(n2720), .I2(n2717), .O(n919) );
  NAND_GATE U1400 ( .I1(n806), .I2(n922), .O(n920) );
  AND_GATE U1401 ( .I1(n920), .I2(n921), .O(n10139) );
  OR_GATE U1402 ( .I1(n10135), .I2(n10134), .O(n921) );
  AND_GATE U1403 ( .I1(n10136), .I2(n10138), .O(n922) );
  NAND_GATE U1404 ( .I1(n702), .I2(n925), .O(n923) );
  AND_GATE U1405 ( .I1(n923), .I2(n924), .O(n3839) );
  OR_GATE U1406 ( .I1(n3831), .I2(n3838), .O(n924) );
  AND_GATE U1407 ( .I1(n3836), .I2(n4454), .O(n925) );
  OR_GATE U1408 ( .I1(n857), .I2(n8395), .O(n8397) );
  AND_GATE U1409 ( .I1(n10956), .I2(n10567), .O(n926) );
  INV_GATE U1410 ( .I1(n926), .O(n10578) );
  AND3_GATE U1411 ( .I1(n10575), .I2(n10570), .I3(n10569), .O(n927) );
  NOR_GATE U1412 ( .I1(n11790), .I2(n11789), .O(n928) );
  AND3_GATE U1413 ( .I1(n3750), .I2(n3585), .I3(n3584), .O(n929) );
  INV_GATE U1414 ( .I1(n929), .O(n3811) );
  OR_GATE U1415 ( .I1(n3914), .I2(n3913), .O(n3916) );
  OR3_GATE U1416 ( .I1(n930), .I2(n931), .I3(n10151), .O(n10154) );
  INV_GATE U1417 ( .I1(n10153), .O(n930) );
  INV_GATE U1418 ( .I1(n10152), .O(n931) );
  AND_GATE U1419 ( .I1(n1444), .I2(A[1]), .O(n932) );
  NAND_GATE U1420 ( .I1(n933), .I2(n4290), .O(n4289) );
  NOR_GATE U1421 ( .I1(n4292), .I2(n4291), .O(n933) );
  AND3_GATE U1422 ( .I1(n5140), .I2(n5139), .I3(n5138), .O(n935) );
  AND3_GATE U1423 ( .I1(n5146), .I2(n5145), .I3(n4776), .O(n937) );
  INV_GATE U1424 ( .I1(n938), .O(n7521) );
  AND_GATE U1425 ( .I1(n5950), .I2(n5949), .O(n939) );
  INV_GATE U1426 ( .I1(n939), .O(n6596) );
  OR_GATE U1427 ( .I1(n5686), .I2(n908), .O(n5689) );
  NAND_GATE U1428 ( .I1(n7601), .I2(n941), .O(n7603) );
  INV_GATE U1429 ( .I1(n7600), .O(n941) );
  NAND_GATE U1430 ( .I1(n4269), .I2(n942), .O(n4271) );
  INV_GATE U1431 ( .I1(n4268), .O(n942) );
  AND_GATE U1432 ( .I1(n868), .I2(n614), .O(\A2[33] ) );
  NAND_GATE U1433 ( .I1(n5934), .I2(n943), .O(n5936) );
  INV_GATE U1434 ( .I1(n5933), .O(n943) );
  NAND_GATE U1435 ( .I1(n5686), .I2(n908), .O(n5690) );
  NAND_GATE U1436 ( .I1(n5188), .I2(n743), .O(n5190) );
  NAND_GATE U1437 ( .I1(n3513), .I2(n944), .O(n3515) );
  INV_GATE U1438 ( .I1(n3520), .O(n944) );
  NAND_GATE U1439 ( .I1(n945), .I2(n13353), .O(n13358) );
  INV_GATE U1440 ( .I1(n13356), .O(n945) );
  NAND_GATE U1441 ( .I1(n946), .I2(n13787), .O(n13792) );
  INV_GATE U1442 ( .I1(n13790), .O(n946) );
  NAND_GATE U1443 ( .I1(n947), .I2(n14228), .O(n14233) );
  INV_GATE U1444 ( .I1(n14231), .O(n947) );
  OR_GATE U1445 ( .I1(n948), .I2(n6703), .O(n6727) );
  INV_GATE U1446 ( .I1(n6702), .O(n948) );
  OR_GATE U1447 ( .I1(n949), .I2(n6830), .O(n6833) );
  INV_GATE U1448 ( .I1(n6831), .O(n949) );
  OR_GATE U1449 ( .I1(n594), .I2(n8502), .O(n8505) );
  OR_GATE U1450 ( .I1(n950), .I2(n10162), .O(n10157) );
  INV_GATE U1451 ( .I1(n10159), .O(n950) );
  OR_GATE U1452 ( .I1(n199), .I2(n7674), .O(n7677) );
  OR_GATE U1453 ( .I1(n9402), .I2(n780), .O(n9413) );
  AND_GATE U1454 ( .I1(n10978), .I2(n10977), .O(n951) );
  OR_GATE U1455 ( .I1(n754), .I2(n10980), .O(n10972) );
  OR_GATE U1456 ( .I1(n8554), .I2(n8564), .O(n8852) );
  OR_GATE U1457 ( .I1(n10234), .I2(n10233), .O(n10552) );
  OR_GATE U1458 ( .I1(n10283), .I2(n1393), .O(n10640) );
  OR_GATE U1459 ( .I1(n952), .I2(n11019), .O(n11023) );
  INV_GATE U1460 ( .I1(n11020), .O(n952) );
  OR_GATE U1461 ( .I1(n953), .I2(n6841), .O(n6844) );
  INV_GATE U1462 ( .I1(n6842), .O(n953) );
  OR_GATE U1463 ( .I1(n954), .I2(n8513), .O(n8516) );
  INV_GATE U1464 ( .I1(n8514), .O(n954) );
  OR_GATE U1465 ( .I1(n955), .I2(n7685), .O(n7688) );
  INV_GATE U1466 ( .I1(n7686), .O(n955) );
  OR_GATE U1467 ( .I1(n7696), .I2(n956), .O(n7698) );
  INV_GATE U1468 ( .I1(n7697), .O(n956) );
  OR_GATE U1469 ( .I1(n957), .I2(n8523), .O(n8525) );
  INV_GATE U1470 ( .I1(n8524), .O(n957) );
  OR_GATE U1471 ( .I1(n958), .I2(n9359), .O(n9361) );
  INV_GATE U1472 ( .I1(n9360), .O(n958) );
  OR_GATE U1473 ( .I1(n6849), .I2(n505), .O(n6850) );
  OR_GATE U1474 ( .I1(n603), .I2(n9351), .O(n9346) );
  OR_GATE U1475 ( .I1(n6861), .I2(n665), .O(n6858) );
  OR_GATE U1476 ( .I1(n13048), .I2(n489), .O(n13050) );
  OR_GATE U1477 ( .I1(n13078), .I2(n959), .O(n13088) );
  INV_GATE U1478 ( .I1(n13079), .O(n959) );
  OR_GATE U1479 ( .I1(n960), .I2(n6808), .O(n6811) );
  INV_GATE U1480 ( .I1(n6809), .O(n960) );
  OR_GATE U1481 ( .I1(n13549), .I2(n961), .O(n13552) );
  INV_GATE U1482 ( .I1(n13553), .O(n961) );
  OR_GATE U1483 ( .I1(n962), .I2(n6819), .O(n6822) );
  INV_GATE U1484 ( .I1(n6820), .O(n962) );
  OR_GATE U1485 ( .I1(n963), .I2(n7653), .O(n7656) );
  INV_GATE U1486 ( .I1(n7654), .O(n963) );
  OR_GATE U1487 ( .I1(n964), .I2(n7663), .O(n7666) );
  INV_GATE U1488 ( .I1(n7664), .O(n964) );
  OR_GATE U1489 ( .I1(n965), .I2(n8480), .O(n8483) );
  INV_GATE U1490 ( .I1(n8481), .O(n965) );
  OR_GATE U1491 ( .I1(n9991), .I2(n966), .O(n9995) );
  INV_GATE U1492 ( .I1(n9993), .O(n966) );
  OR_GATE U1493 ( .I1(n11431), .I2(n11439), .O(n11739) );
  OR_GATE U1494 ( .I1(n13104), .I2(n967), .O(n13067) );
  INV_GATE U1495 ( .I1(n13107), .O(n967) );
  OR_GATE U1496 ( .I1(n12284), .I2(n78), .O(n12719) );
  OR_GATE U1497 ( .I1(n10883), .I2(n10886), .O(n11326) );
  OR_GATE U1498 ( .I1(n10920), .I2(n884), .O(n11040) );
  AND_GATE U1499 ( .I1(n10923), .I2(n10925), .O(n968) );
  OR_GATE U1500 ( .I1(n9385), .I2(n969), .O(n9390) );
  INV_GATE U1501 ( .I1(n9386), .O(n969) );
  AND_GATE U1502 ( .I1(n13924), .I2(n13923), .O(n970) );
  OR_GATE U1503 ( .I1(n20), .I2(n9794), .O(n9801) );
  OR_GATE U1504 ( .I1(n13895), .I2(n13893), .O(n13965) );
  OR_GATE U1505 ( .I1(n971), .I2(n6941), .O(n6954) );
  INV_GATE U1506 ( .I1(n6942), .O(n971) );
  OR_GATE U1507 ( .I1(n7367), .I2(n7369), .O(n7903) );
  OR_GATE U1508 ( .I1(n972), .I2(n6711), .O(n6715) );
  INV_GATE U1509 ( .I1(n6712), .O(n972) );
  OR_GATE U1510 ( .I1(n11858), .I2(n11857), .O(n11864) );
  OR_GATE U1511 ( .I1(n12256), .I2(n12257), .O(n12260) );
  OR_GATE U1512 ( .I1(n973), .I2(n6798), .O(n6801) );
  INV_GATE U1513 ( .I1(n6799), .O(n973) );
  OR_GATE U1514 ( .I1(n974), .I2(n7643), .O(n7646) );
  INV_GATE U1515 ( .I1(n7644), .O(n974) );
  OR_GATE U1516 ( .I1(n975), .I2(n8470), .O(n8473) );
  INV_GATE U1517 ( .I1(n8471), .O(n975) );
  OR_GATE U1518 ( .I1(n976), .I2(n9305), .O(n9308) );
  INV_GATE U1519 ( .I1(n9306), .O(n976) );
  OR_GATE U1520 ( .I1(n11726), .I2(n977), .O(n11894) );
  INV_GATE U1521 ( .I1(n11730), .O(n977) );
  OR_GATE U1522 ( .I1(n14356), .I2(n978), .O(n13917) );
  INV_GATE U1523 ( .I1(n14357), .O(n978) );
  OR_GATE U1524 ( .I1(n10076), .I2(n979), .O(n10243) );
  INV_GATE U1525 ( .I1(n10078), .O(n979) );
  OR_GATE U1526 ( .I1(n11744), .I2(n980), .O(n11755) );
  INV_GATE U1527 ( .I1(n11747), .O(n980) );
  OR_GATE U1528 ( .I1(n11372), .I2(n1389), .O(n11380) );
  OR_GATE U1529 ( .I1(n7952), .I2(n761), .O(n8289) );
  OR_GATE U1530 ( .I1(n8834), .I2(n8832), .O(n8943) );
  OR_GATE U1531 ( .I1(n10605), .I2(n981), .O(n10608) );
  INV_GATE U1532 ( .I1(n10606), .O(n981) );
  OR_GATE U1533 ( .I1(n9479), .I2(n9476), .O(n9993) );
  OR_GATE U1534 ( .I1(n12297), .I2(n12302), .O(n12725) );
  OR_GATE U1535 ( .I1(n9683), .I2(n9686), .O(n9759) );
  OR_GATE U1536 ( .I1(n982), .I2(n6787), .O(n6790) );
  INV_GATE U1537 ( .I1(n6788), .O(n982) );
  OR_GATE U1538 ( .I1(n983), .I2(n7633), .O(n7636) );
  INV_GATE U1539 ( .I1(n7634), .O(n983) );
  OR_GATE U1540 ( .I1(n984), .I2(n8460), .O(n8463) );
  INV_GATE U1541 ( .I1(n8461), .O(n984) );
  OR_GATE U1542 ( .I1(n8249), .I2(n985), .O(n8797) );
  INV_GATE U1543 ( .I1(n8251), .O(n985) );
  OR_GATE U1544 ( .I1(n6735), .I2(n6744), .O(n6746) );
  OR_GATE U1545 ( .I1(n986), .I2(n6765), .O(n6768) );
  INV_GATE U1546 ( .I1(n6766), .O(n986) );
  OR_GATE U1547 ( .I1(n987), .I2(n6776), .O(n6779) );
  INV_GATE U1548 ( .I1(n6777), .O(n987) );
  OR_GATE U1549 ( .I1(n988), .I2(n7622), .O(n7625) );
  INV_GATE U1550 ( .I1(n7623), .O(n988) );
  OR_GATE U1551 ( .I1(n989), .I2(n8449), .O(n8452) );
  INV_GATE U1552 ( .I1(n8450), .O(n989) );
  OR_GATE U1553 ( .I1(n990), .I2(n7611), .O(n7614) );
  INV_GATE U1554 ( .I1(n7612), .O(n990) );
  NOR_GATE U1555 ( .I1(n14382), .I2(n14376), .O(\A2[31] ) );
  OR_GATE U1556 ( .I1(n10111), .I2(n991), .O(n10200) );
  INV_GATE U1557 ( .I1(n10113), .O(n991) );
  AND_GATE U1558 ( .I1(n11769), .I2(n11847), .O(n992) );
  OR_GATE U1559 ( .I1(n939), .I2(n6598), .O(n6600) );
  AND_GATE U1560 ( .I1(n12656), .I2(n12658), .O(n993) );
  OR_GATE U1561 ( .I1(n910), .I2(n7508), .O(n7510) );
  OR_GATE U1562 ( .I1(n347), .I2(n6557), .O(n6555) );
  OR_GATE U1563 ( .I1(n641), .I2(n13495), .O(n13490) );
  OR_GATE U1564 ( .I1(n77), .I2(n11448), .O(n11444) );
  OR_GATE U1565 ( .I1(n469), .I2(n11075), .O(n11077) );
  OR_GATE U1566 ( .I1(n10121), .I2(n10120), .O(n10124) );
  OR_GATE U1567 ( .I1(n994), .I2(n8535), .O(n8537) );
  INV_GATE U1568 ( .I1(n8534), .O(n994) );
  OR_GATE U1569 ( .I1(n8322), .I2(n8321), .O(n8324) );
  OR_GATE U1570 ( .I1(n11907), .I2(n11906), .O(n11909) );
  OR_GATE U1571 ( .I1(n695), .I2(n10645), .O(n10648) );
  OR_GATE U1572 ( .I1(n7430), .I2(n7434), .O(n7431) );
  OR_GATE U1573 ( .I1(n995), .I2(n12663), .O(n12665) );
  INV_GATE U1574 ( .I1(n12664), .O(n995) );
  OR_GATE U1575 ( .I1(n996), .I2(n11935), .O(n11938) );
  INV_GATE U1576 ( .I1(n11936), .O(n996) );
  OR_GATE U1577 ( .I1(n997), .I2(n14361), .O(n14364) );
  INV_GATE U1578 ( .I1(n14362), .O(n997) );
  OR_GATE U1579 ( .I1(n110), .I2(n11469), .O(n11472) );
  OR_GATE U1580 ( .I1(n998), .I2(n10847), .O(n10850) );
  INV_GATE U1581 ( .I1(n10846), .O(n998) );
  OR_GATE U1582 ( .I1(n124), .I2(n13136), .O(n13139) );
  OR_GATE U1583 ( .I1(n999), .I2(n11945), .O(n11948) );
  INV_GATE U1584 ( .I1(n11946), .O(n999) );
  OR_GATE U1585 ( .I1(n10486), .I2(n1000), .O(n10489) );
  INV_GATE U1586 ( .I1(n10487), .O(n1000) );
  OR_GATE U1587 ( .I1(n11287), .I2(n1001), .O(n11290) );
  INV_GATE U1588 ( .I1(n11288), .O(n1001) );
  OR_GATE U1589 ( .I1(n8255), .I2(n1002), .O(n8257) );
  INV_GATE U1590 ( .I1(n8260), .O(n1002) );
  OR_GATE U1591 ( .I1(n10831), .I2(n1003), .O(n10834) );
  INV_GATE U1592 ( .I1(n10832), .O(n1003) );
  OR_GATE U1593 ( .I1(n1004), .I2(n13969), .O(n13972) );
  INV_GATE U1594 ( .I1(n13970), .O(n1004) );
  OR_GATE U1595 ( .I1(n13016), .I2(n1005), .O(n13019) );
  INV_GATE U1596 ( .I1(n13017), .O(n1005) );
  OR_GATE U1597 ( .I1(n11674), .I2(n1006), .O(n11677) );
  INV_GATE U1598 ( .I1(n11675), .O(n1006) );
  OR_GATE U1599 ( .I1(n12566), .I2(n1007), .O(n12569) );
  INV_GATE U1600 ( .I1(n12567), .O(n1007) );
  OR_GATE U1601 ( .I1(n10471), .I2(n1008), .O(n10474) );
  INV_GATE U1602 ( .I1(n10472), .O(n1008) );
  OR_GATE U1603 ( .I1(n13871), .I2(n1009), .O(n13874) );
  INV_GATE U1604 ( .I1(n13872), .O(n1009) );
  OR_GATE U1605 ( .I1(n9109), .I2(n1010), .O(n9112) );
  INV_GATE U1606 ( .I1(n9110), .O(n1010) );
  OR_GATE U1607 ( .I1(n13422), .I2(n1011), .O(n13425) );
  INV_GATE U1608 ( .I1(n13423), .O(n1011) );
  OR_GATE U1609 ( .I1(n8733), .I2(n1012), .O(n8736) );
  INV_GATE U1610 ( .I1(n8734), .O(n1012) );
  OR3_GATE U1611 ( .I1(n1013), .I2(n1014), .I3(n1396), .O(n6903) );
  INV_GATE U1612 ( .I1(n6909), .O(n1013) );
  AND3_GATE U1613 ( .I1(n6914), .I2(n6520), .I3(n6916), .O(n1014) );
  OR_GATE U1614 ( .I1(n1298), .I2(n1015), .O(n7053) );
  NAND_GATE U1615 ( .I1(n1343), .I2(n1344), .O(n1015) );
  OR_GATE U1616 ( .I1(n10252), .I2(n10253), .O(n10923) );
  OR_GATE U1617 ( .I1(n5873), .I2(n402), .O(n6688) );
  AND_GATE U1618 ( .I1(n13108), .I2(n13067), .O(n1016) );
  OR_GATE U1619 ( .I1(n8923), .I2(n1017), .O(n8925) );
  INV_GATE U1620 ( .I1(n8924), .O(n1017) );
  OR_GATE U1621 ( .I1(n8906), .I2(n1018), .O(n9373) );
  INV_GATE U1622 ( .I1(n8908), .O(n1018) );
  OR_GATE U1623 ( .I1(n7196), .I2(n784), .O(n7710) );
  OR_GATE U1624 ( .I1(n797), .I2(n6613), .O(n6615) );
  OR_GATE U1625 ( .I1(n84), .I2(n12199), .O(n12200) );
  OR_GATE U1626 ( .I1(n938), .I2(n7523), .O(n7525) );
  OR_GATE U1627 ( .I1(n13146), .I2(n13148), .O(n13142) );
  OR_GATE U1628 ( .I1(n6052), .I2(n1285), .O(n6344) );
  OR_GATE U1629 ( .I1(n763), .I2(n8409), .O(n8411) );
  OR_GATE U1630 ( .I1(n1019), .I2(n7105), .O(n7110) );
  INV_GATE U1631 ( .I1(n7106), .O(n1019) );
  OR_GATE U1632 ( .I1(n726), .I2(n8899), .O(n8900) );
  OR_GATE U1633 ( .I1(n7802), .I2(n7803), .O(n8202) );
  OR_GATE U1634 ( .I1(n6938), .I2(n6940), .O(n7057) );
  OR_GATE U1635 ( .I1(n642), .I2(n13535), .O(n13531) );
  OR_GATE U1636 ( .I1(n12701), .I2(n1020), .O(n13488) );
  INV_GATE U1637 ( .I1(n12705), .O(n1020) );
  OR_GATE U1638 ( .I1(n8552), .I2(n8553), .O(n8851) );
  OR_GATE U1639 ( .I1(n1021), .I2(n11332), .O(n11328) );
  INV_GATE U1640 ( .I1(n11327), .O(n1021) );
  OR_GATE U1641 ( .I1(n11440), .I2(n11436), .O(n11433) );
  OR_GATE U1642 ( .I1(n7724), .I2(n306), .O(n7721) );
  OR_GATE U1643 ( .I1(n1022), .I2(n10297), .O(n10299) );
  INV_GATE U1644 ( .I1(n10296), .O(n1022) );
  OR_GATE U1645 ( .I1(n1024), .I2(n8931), .O(n8933) );
  INV_GATE U1646 ( .I1(n8932), .O(n1024) );
  OR_GATE U1647 ( .I1(n129), .I2(n11084), .O(n11087) );
  OR_GATE U1648 ( .I1(n134), .I2(n12313), .O(n12308) );
  OR_GATE U1649 ( .I1(n1025), .I2(n9454), .O(n9456) );
  INV_GATE U1650 ( .I1(n9453), .O(n1025) );
  OR_GATE U1651 ( .I1(n10497), .I2(n1026), .O(n10499) );
  INV_GATE U1652 ( .I1(n10502), .O(n1026) );
  OR_GATE U1653 ( .I1(n9646), .I2(n1027), .O(n9648) );
  INV_GATE U1654 ( .I1(n9651), .O(n1027) );
  OR_GATE U1655 ( .I1(n479), .I2(n12741), .O(n12744) );
  OR_GATE U1656 ( .I1(n1028), .I2(n12321), .O(n12324) );
  INV_GATE U1657 ( .I1(n12322), .O(n1028) );
  OR_GATE U1658 ( .I1(n9636), .I2(n1029), .O(n9632) );
  INV_GATE U1659 ( .I1(n9635), .O(n1029) );
  OR_GATE U1660 ( .I1(n13558), .I2(n13565), .O(n13560) );
  OR_GATE U1661 ( .I1(n1030), .I2(n9140), .O(n9142) );
  INV_GATE U1662 ( .I1(n9144), .O(n1030) );
  OR_GATE U1663 ( .I1(n13436), .I2(n1031), .O(n13439) );
  INV_GATE U1664 ( .I1(n13437), .O(n1031) );
  OR_GATE U1665 ( .I1(n1032), .I2(n7927), .O(n7929) );
  INV_GATE U1666 ( .I1(n7926), .O(n1032) );
  OR_GATE U1667 ( .I1(n14295), .I2(n1033), .O(n14298) );
  INV_GATE U1668 ( .I1(n14296), .O(n1033) );
  OR_GATE U1669 ( .I1(n7382), .I2(n1346), .O(n7384) );
  OR_GATE U1670 ( .I1(n11273), .I2(n1034), .O(n11276) );
  INV_GATE U1671 ( .I1(n11274), .O(n1034) );
  OR_GATE U1672 ( .I1(n10817), .I2(n1035), .O(n10820) );
  INV_GATE U1673 ( .I1(n10818), .O(n1035) );
  OR_GATE U1674 ( .I1(n11967), .I2(n1036), .O(n11970) );
  INV_GATE U1675 ( .I1(n11968), .O(n1036) );
  OR_GATE U1676 ( .I1(n13002), .I2(n1037), .O(n13005) );
  INV_GATE U1677 ( .I1(n13003), .O(n1037) );
  OR_GATE U1678 ( .I1(n9963), .I2(n1038), .O(n9966) );
  INV_GATE U1679 ( .I1(n9964), .O(n1038) );
  OR_GATE U1680 ( .I1(n11492), .I2(n1039), .O(n11495) );
  INV_GATE U1681 ( .I1(n11493), .O(n1039) );
  OR_GATE U1682 ( .I1(n9095), .I2(n1040), .O(n9098) );
  INV_GATE U1683 ( .I1(n9096), .O(n1040) );
  OR_GATE U1684 ( .I1(n13407), .I2(n1041), .O(n13410) );
  INV_GATE U1685 ( .I1(n13408), .O(n1041) );
  OR_GATE U1686 ( .I1(n12354), .I2(n1042), .O(n12357) );
  INV_GATE U1687 ( .I1(n12355), .O(n1042) );
  OR_GATE U1688 ( .I1(n1043), .I2(n7280), .O(n7274) );
  INV_GATE U1689 ( .I1(n7277), .O(n1043) );
  OR_GATE U1690 ( .I1(n7030), .I2(n1044), .O(n7038) );
  INV_GATE U1691 ( .I1(n7039), .O(n1044) );
  OR_GATE U1692 ( .I1(n14018), .I2(n1045), .O(n14021) );
  INV_GATE U1693 ( .I1(n14019), .O(n1045) );
  OR_GATE U1694 ( .I1(n7775), .I2(n7779), .O(n7787) );
  OR_GATE U1695 ( .I1(n6745), .I2(n6747), .O(n7158) );
  OR_GATE U1696 ( .I1(n6674), .I2(n6673), .O(n6676) );
  OR_GATE U1697 ( .I1(n6303), .I2(n6302), .O(n6305) );
  OR_GATE U1698 ( .I1(n750), .I2(n6628), .O(n6630) );
  OR_GATE U1699 ( .I1(n318), .I2(n7538), .O(n7540) );
  OR_GATE U1700 ( .I1(n11314), .I2(n11313), .O(n11315) );
  OR_GATE U1701 ( .I1(n824), .I2(n8424), .O(n8426) );
  AND_GATE U1702 ( .I1(n13539), .I2(n13540), .O(n1046) );
  OR_GATE U1703 ( .I1(n799), .I2(n8888), .O(n8889) );
  OR_GATE U1704 ( .I1(n6658), .I2(n6657), .O(n6660) );
  OR_GATE U1705 ( .I1(n6686), .I2(n6687), .O(n6699) );
  OR_GATE U1706 ( .I1(n1047), .I2(n10631), .O(n10634) );
  INV_GATE U1707 ( .I1(n10632), .O(n1047) );
  OR_GATE U1708 ( .I1(n58), .I2(n10873), .O(n10875) );
  OR_GATE U1709 ( .I1(n657), .I2(n9445), .O(n9439) );
  OR_GATE U1710 ( .I1(n10016), .I2(n1048), .O(n10018) );
  INV_GATE U1711 ( .I1(n10015), .O(n1048) );
  OR_GATE U1712 ( .I1(n9277), .I2(n858), .O(n9287) );
  OR_GATE U1713 ( .I1(n13885), .I2(n491), .O(n13888) );
  OR_GATE U1714 ( .I1(n13856), .I2(n1049), .O(n13859) );
  INV_GATE U1715 ( .I1(n13857), .O(n1049) );
  OR_GATE U1716 ( .I1(n13992), .I2(n1050), .O(n13995) );
  INV_GATE U1717 ( .I1(n13993), .O(n1050) );
  OR_GATE U1718 ( .I1(n10457), .I2(n1051), .O(n10460) );
  INV_GATE U1719 ( .I1(n10458), .O(n1051) );
  OR_GATE U1720 ( .I1(n11120), .I2(n1052), .O(n11123) );
  INV_GATE U1721 ( .I1(n11121), .O(n1052) );
  OR_GATE U1722 ( .I1(n9592), .I2(n1053), .O(n9595) );
  INV_GATE U1723 ( .I1(n9593), .O(n1053) );
  OR_GATE U1724 ( .I1(n11992), .I2(n1054), .O(n11995) );
  INV_GATE U1725 ( .I1(n11993), .O(n1054) );
  OR_GATE U1726 ( .I1(n13841), .I2(n1055), .O(n13844) );
  INV_GATE U1727 ( .I1(n13842), .O(n1055) );
  OR_GATE U1728 ( .I1(n12789), .I2(n1056), .O(n12792) );
  INV_GATE U1729 ( .I1(n12790), .O(n1056) );
  OR_GATE U1730 ( .I1(n8376), .I2(n8377), .O(n8388) );
  OR_GATE U1731 ( .I1(n1057), .I2(n6926), .O(n6930) );
  INV_GATE U1732 ( .I1(n6927), .O(n1057) );
  OR_GATE U1733 ( .I1(n10692), .I2(n1058), .O(n10695) );
  INV_GATE U1734 ( .I1(n10693), .O(n1058) );
  OR_GATE U1735 ( .I1(n9949), .I2(n1059), .O(n9952) );
  INV_GATE U1736 ( .I1(n9950), .O(n1059) );
  OR_GATE U1737 ( .I1(n11516), .I2(n1060), .O(n11519) );
  INV_GATE U1738 ( .I1(n11517), .O(n1060) );
  OR_GATE U1739 ( .I1(n12378), .I2(n1061), .O(n12381) );
  INV_GATE U1740 ( .I1(n12379), .O(n1061) );
  OR_GATE U1741 ( .I1(n13194), .I2(n1062), .O(n13197) );
  INV_GATE U1742 ( .I1(n13195), .O(n1062) );
  OR_GATE U1743 ( .I1(n14044), .I2(n1063), .O(n14047) );
  INV_GATE U1744 ( .I1(n14045), .O(n1063) );
  OR_GATE U1745 ( .I1(n10361), .I2(n1064), .O(n10364) );
  INV_GATE U1746 ( .I1(n10362), .O(n1064) );
  OR_GATE U1747 ( .I1(n11144), .I2(n1065), .O(n11147) );
  INV_GATE U1748 ( .I1(n11145), .O(n1065) );
  OR_GATE U1749 ( .I1(n12016), .I2(n1066), .O(n12019) );
  INV_GATE U1750 ( .I1(n12017), .O(n1066) );
  OR_GATE U1751 ( .I1(n12814), .I2(n1067), .O(n12817) );
  INV_GATE U1752 ( .I1(n12815), .O(n1067) );
  OR_GATE U1753 ( .I1(n13628), .I2(n1068), .O(n13631) );
  INV_GATE U1754 ( .I1(n13629), .O(n1068) );
  OR_GATE U1755 ( .I1(n10716), .I2(n1069), .O(n10719) );
  INV_GATE U1756 ( .I1(n10717), .O(n1069) );
  OR_GATE U1757 ( .I1(n11540), .I2(n1070), .O(n11543) );
  INV_GATE U1758 ( .I1(n11541), .O(n1070) );
  OR_GATE U1759 ( .I1(n12403), .I2(n1071), .O(n12406) );
  INV_GATE U1760 ( .I1(n12404), .O(n1071) );
  OR_GATE U1761 ( .I1(n13219), .I2(n1072), .O(n13222) );
  INV_GATE U1762 ( .I1(n13220), .O(n1072) );
  OR_GATE U1763 ( .I1(n14069), .I2(n1073), .O(n14072) );
  INV_GATE U1764 ( .I1(n14070), .O(n1073) );
  OR_GATE U1765 ( .I1(n11168), .I2(n1074), .O(n11171) );
  INV_GATE U1766 ( .I1(n11169), .O(n1074) );
  OR_GATE U1767 ( .I1(n12041), .I2(n1075), .O(n12044) );
  INV_GATE U1768 ( .I1(n12042), .O(n1075) );
  OR_GATE U1769 ( .I1(n12839), .I2(n1076), .O(n12842) );
  INV_GATE U1770 ( .I1(n12840), .O(n1076) );
  OR_GATE U1771 ( .I1(n13653), .I2(n1077), .O(n13656) );
  INV_GATE U1772 ( .I1(n13654), .O(n1077) );
  OR_GATE U1773 ( .I1(n13244), .I2(n1078), .O(n13247) );
  INV_GATE U1774 ( .I1(n13245), .O(n1078) );
  OR_GATE U1775 ( .I1(n12428), .I2(n1079), .O(n12431) );
  INV_GATE U1776 ( .I1(n12429), .O(n1079) );
  OR_GATE U1777 ( .I1(n11565), .I2(n1080), .O(n11568) );
  INV_GATE U1778 ( .I1(n11566), .O(n1080) );
  OR_GATE U1779 ( .I1(n14094), .I2(n1081), .O(n14097) );
  INV_GATE U1780 ( .I1(n14095), .O(n1081) );
  OR_GATE U1781 ( .I1(n12864), .I2(n1082), .O(n12867) );
  INV_GATE U1782 ( .I1(n12865), .O(n1082) );
  OR_GATE U1783 ( .I1(n12066), .I2(n1083), .O(n12069) );
  INV_GATE U1784 ( .I1(n12067), .O(n1083) );
  OR_GATE U1785 ( .I1(n13678), .I2(n1084), .O(n13681) );
  INV_GATE U1786 ( .I1(n13679), .O(n1084) );
  OR_GATE U1787 ( .I1(n13269), .I2(n1085), .O(n13272) );
  INV_GATE U1788 ( .I1(n13270), .O(n1085) );
  OR_GATE U1789 ( .I1(n12453), .I2(n1086), .O(n12456) );
  INV_GATE U1790 ( .I1(n12454), .O(n1086) );
  OR_GATE U1791 ( .I1(n14119), .I2(n1087), .O(n14122) );
  INV_GATE U1792 ( .I1(n14120), .O(n1087) );
  OR_GATE U1793 ( .I1(n12889), .I2(n1088), .O(n12892) );
  INV_GATE U1794 ( .I1(n12890), .O(n1088) );
  OR_GATE U1795 ( .I1(n13703), .I2(n1089), .O(n13706) );
  INV_GATE U1796 ( .I1(n13704), .O(n1089) );
  OR_GATE U1797 ( .I1(n7175), .I2(n7174), .O(n7177) );
  OR_GATE U1798 ( .I1(n13294), .I2(n1090), .O(n13297) );
  INV_GATE U1799 ( .I1(n13295), .O(n1090) );
  OR_GATE U1800 ( .I1(n14144), .I2(n1091), .O(n14147) );
  INV_GATE U1801 ( .I1(n14145), .O(n1091) );
  OR_GATE U1802 ( .I1(n13728), .I2(n1092), .O(n13731) );
  INV_GATE U1803 ( .I1(n13729), .O(n1092) );
  OR_GATE U1804 ( .I1(n14169), .I2(n1093), .O(n14172) );
  INV_GATE U1805 ( .I1(n14170), .O(n1093) );
  OR_GATE U1806 ( .I1(n14412), .I2(n794), .O(n14414) );
  OR_GATE U1807 ( .I1(n1094), .I2(n4301), .O(n4304) );
  INV_GATE U1808 ( .I1(n4302), .O(n1094) );
  OR_GATE U1809 ( .I1(n1095), .I2(n5128), .O(n5123) );
  INV_GATE U1810 ( .I1(n5125), .O(n1095) );
  OR_GATE U1811 ( .I1(n180), .I2(n6252), .O(n6255) );
  OR_GATE U1812 ( .I1(n10193), .I2(n10194), .O(n10197) );
  NOR_GATE U1813 ( .I1(n13092), .I2(n12645), .O(\A2[35] ) );
  OR_GATE U1814 ( .I1(n1096), .I2(n12597), .O(n12598) );
  INV_GATE U1815 ( .I1(n13046), .O(n1096) );
  NOR_GATE U1816 ( .I1(n11796), .I2(n12238), .O(\A2[37] ) );
  OR_GATE U1817 ( .I1(n1271), .I2(n1097), .O(n11010) );
  AND_GATE U1818 ( .I1(n11009), .I2(n11008), .O(n1097) );
  OR_GATE U1819 ( .I1(n3730), .I2(n731), .O(n3830) );
  OR_GATE U1820 ( .I1(n3589), .I2(n3591), .O(n3608) );
  OR_GATE U1821 ( .I1(n1289), .I2(n1098), .O(n8340) );
  AND_GATE U1822 ( .I1(n8326), .I2(n7983), .O(n1098) );
  OR_GATE U1823 ( .I1(n1383), .I2(n1099), .O(n11892) );
  AND_GATE U1824 ( .I1(n11911), .I2(n11723), .O(n1099) );
  OR_GATE U1825 ( .I1(n937), .I2(n5137), .O(n5133) );
  OR_GATE U1826 ( .I1(n370), .I2(n3476), .O(n3479) );
  OR_GATE U1827 ( .I1(n1100), .I2(n5966), .O(n5969) );
  INV_GATE U1828 ( .I1(n5967), .O(n1100) );
  OR_GATE U1829 ( .I1(n10119), .I2(n1101), .O(n10122) );
  AND_GATE U1830 ( .I1(n10121), .I2(n10120), .O(n1101) );
  OR_GATE U1831 ( .I1(n8320), .I2(n1102), .O(n8325) );
  AND_GATE U1832 ( .I1(n8322), .I2(n8321), .O(n1102) );
  OR_GATE U1833 ( .I1(n5144), .I2(n909), .O(n5141) );
  OR_GATE U1834 ( .I1(n13046), .I2(n1103), .O(n13049) );
  AND_GATE U1835 ( .I1(n13048), .I2(n489), .O(n1103) );
  OR_GATE U1836 ( .I1(n3498), .I2(n1104), .O(n3494) );
  INV_GATE U1837 ( .I1(n3497), .O(n1104) );
  OR_GATE U1838 ( .I1(n704), .I2(n5157), .O(n5151) );
  OR_GATE U1839 ( .I1(n319), .I2(n2657), .O(n2660) );
  OR_GATE U1840 ( .I1(n700), .I2(n5955), .O(n5958) );
  OR_GATE U1841 ( .I1(n1105), .I2(n2648), .O(n2644) );
  INV_GATE U1842 ( .I1(n2645), .O(n1105) );
  OR_GATE U1843 ( .I1(n4332), .I2(n1266), .O(n4329) );
  OR_GATE U1844 ( .I1(n2637), .I2(n1106), .O(n2640) );
  INV_GATE U1845 ( .I1(n2636), .O(n1106) );
  OR_GATE U1846 ( .I1(n6183), .I2(n6185), .O(n6181) );
  OR_GATE U1847 ( .I1(n1356), .I2(n1107), .O(n11836) );
  AND_GATE U1848 ( .I1(n11849), .I2(n11383), .O(n1107) );
  OR_GATE U1849 ( .I1(n1108), .I2(n1362), .O(n8082) );
  AND_GATE U1850 ( .I1(n8594), .I2(n8593), .O(n1108) );
  OR_GATE U1851 ( .I1(n8636), .I2(n1109), .O(n8209) );
  AND_GATE U1852 ( .I1(n8643), .I2(n8637), .O(n1109) );
  OR_GATE U1853 ( .I1(n6153), .I2(n6157), .O(n6396) );
  OR_GATE U1854 ( .I1(n11850), .I2(n1110), .O(n11854) );
  AND_GATE U1855 ( .I1(n11851), .I2(n372), .O(n1110) );
  OR_GATE U1856 ( .I1(n1111), .I2(n6021), .O(n6026) );
  INV_GATE U1857 ( .I1(n6022), .O(n1111) );
  OR_GATE U1858 ( .I1(n1392), .I2(n1112), .O(n8228) );
  AND_GATE U1859 ( .I1(n8227), .I2(n8226), .O(n1112) );
  OR_GATE U1860 ( .I1(n6420), .I2(n6419), .O(n6423) );
  OR_GATE U1861 ( .I1(n1284), .I2(n1113), .O(n9749) );
  AND_GATE U1862 ( .I1(n10125), .I2(n9702), .O(n1113) );
  OR_GATE U1863 ( .I1(n13516), .I2(n1114), .O(n13519) );
  AND_GATE U1864 ( .I1(n13518), .I2(n1387), .O(n1114) );
  OR_GATE U1865 ( .I1(n11355), .I2(n1115), .O(n11361) );
  AND_GATE U1866 ( .I1(n11357), .I2(n11356), .O(n1115) );
  OR_GATE U1867 ( .I1(n1116), .I2(n4290), .O(n4293) );
  INV_GATE U1868 ( .I1(n4291), .O(n1116) );
  OR_GATE U1869 ( .I1(n1117), .I2(n5093), .O(n5096) );
  INV_GATE U1870 ( .I1(n5094), .O(n1117) );
  OR_GATE U1871 ( .I1(n5872), .I2(n5868), .O(n5865) );
  OR_GATE U1872 ( .I1(n5944), .I2(n1118), .O(n5947) );
  INV_GATE U1873 ( .I1(n5945), .O(n1118) );
  OR_GATE U1874 ( .I1(n1119), .I2(n5104), .O(n5107) );
  INV_GATE U1875 ( .I1(n5105), .O(n1119) );
  OR_GATE U1876 ( .I1(n1120), .I2(n5115), .O(n5118) );
  INV_GATE U1877 ( .I1(n5116), .O(n1120) );
  OR_GATE U1878 ( .I1(n1121), .I2(n4222), .O(n4225) );
  INV_GATE U1879 ( .I1(n4223), .O(n1121) );
  OR_GATE U1880 ( .I1(n1122), .I2(n5040), .O(n5043) );
  INV_GATE U1881 ( .I1(n5041), .O(n1122) );
  OR_GATE U1882 ( .I1(n1123), .I2(n4211), .O(n4214) );
  INV_GATE U1883 ( .I1(n4212), .O(n1123) );
  OR_GATE U1884 ( .I1(n1124), .I2(n4279), .O(n4282) );
  INV_GATE U1885 ( .I1(n4280), .O(n1124) );
  OR_GATE U1886 ( .I1(n1125), .I2(n3465), .O(n3468) );
  INV_GATE U1887 ( .I1(n3466), .O(n1125) );
  NAND_GATE U1888 ( .I1(n7957), .I2(n1126), .O(n1358) );
  AND_GATE U1889 ( .I1(n7955), .I2(n761), .O(n1126) );
  OR_GATE U1890 ( .I1(n1127), .I2(n3407), .O(n3410) );
  INV_GATE U1891 ( .I1(n3408), .O(n1127) );
  OR_GATE U1892 ( .I1(n321), .I2(n3454), .O(n3457) );
  OR_GATE U1893 ( .I1(n7381), .I2(n1128), .O(n7385) );
  AND_GATE U1894 ( .I1(n7382), .I2(n1346), .O(n1128) );
  OR_GATE U1895 ( .I1(n1129), .I2(n3383), .O(n3386) );
  INV_GATE U1896 ( .I1(n3384), .O(n1129) );
  OR_GATE U1897 ( .I1(n1130), .I2(n2625), .O(n2628) );
  INV_GATE U1898 ( .I1(n2626), .O(n1130) );
  OR_GATE U1899 ( .I1(n1131), .I2(n2581), .O(n2584) );
  INV_GATE U1900 ( .I1(n2582), .O(n1131) );
  OR_GATE U1901 ( .I1(n2571), .I2(n1132), .O(n2574) );
  INV_GATE U1902 ( .I1(n2570), .O(n1132) );
  OR_GATE U1903 ( .I1(n1133), .I2(n2559), .O(n2562) );
  INV_GATE U1904 ( .I1(n2560), .O(n1133) );
  OR_GATE U1905 ( .I1(n8185), .I2(n1134), .O(n8188) );
  INV_GATE U1906 ( .I1(n8186), .O(n1134) );
  NOR_GATE U1907 ( .I1(n9428), .I2(n1135), .O(n1276) );
  AND_GATE U1908 ( .I1(n8923), .I2(n1017), .O(n1135) );
  OR_GATE U1909 ( .I1(n1136), .I2(n6366), .O(n6370) );
  INV_GATE U1910 ( .I1(n6367), .O(n1136) );
  OR_GATE U1911 ( .I1(n6063), .I2(n1137), .O(n6067) );
  INV_GATE U1912 ( .I1(n6064), .O(n1137) );
  OR_GATE U1913 ( .I1(n10858), .I2(n1138), .O(n10506) );
  AND_GATE U1914 ( .I1(n10861), .I2(n10859), .O(n1138) );
  OR_GATE U1915 ( .I1(n5890), .I2(n1139), .O(n5893) );
  INV_GATE U1916 ( .I1(n5889), .O(n1139) );
  OR_GATE U1917 ( .I1(n5901), .I2(n1140), .O(n5904) );
  INV_GATE U1918 ( .I1(n5900), .O(n1140) );
  OR_GATE U1919 ( .I1(n1141), .I2(n5911), .O(n5914) );
  INV_GATE U1920 ( .I1(n5912), .O(n1141) );
  OR_GATE U1921 ( .I1(n1142), .I2(n5922), .O(n5925) );
  INV_GATE U1922 ( .I1(n5923), .O(n1142) );
  OR3_GATE U1923 ( .I1(n12258), .I2(n1143), .I3(n1144), .O(n12261) );
  NOR_GATE U1924 ( .I1(n12263), .I2(n12255), .O(n1143) );
  AND_GATE U1925 ( .I1(n11866), .I2(n12257), .O(n1144) );
  OR_GATE U1926 ( .I1(n1145), .I2(n5060), .O(n5063) );
  INV_GATE U1927 ( .I1(n5061), .O(n1145) );
  OR_GATE U1928 ( .I1(n1146), .I2(n5050), .O(n5053) );
  INV_GATE U1929 ( .I1(n5051), .O(n1146) );
  OR_GATE U1930 ( .I1(n1385), .I2(n1147), .O(n11039) );
  AND_GATE U1931 ( .I1(n11044), .I2(n11043), .O(n1147) );
  OR_GATE U1932 ( .I1(n1148), .I2(n4246), .O(n4249) );
  INV_GATE U1933 ( .I1(n4247), .O(n1148) );
  OR_GATE U1934 ( .I1(n1149), .I2(n4257), .O(n4260) );
  INV_GATE U1935 ( .I1(n4258), .O(n1149) );
  OR_GATE U1936 ( .I1(n1150), .I2(n4498), .O(n4501) );
  INV_GATE U1937 ( .I1(n4499), .O(n1150) );
  OR_GATE U1938 ( .I1(n1151), .I2(n3431), .O(n3434) );
  INV_GATE U1939 ( .I1(n3432), .O(n1151) );
  OR_GATE U1940 ( .I1(n2593), .I2(n1152), .O(n2596) );
  INV_GATE U1941 ( .I1(n2592), .O(n1152) );
  OR_GATE U1942 ( .I1(n1153), .I2(n2603), .O(n2606) );
  INV_GATE U1943 ( .I1(n2604), .O(n1153) );
  OR_GATE U1944 ( .I1(n2615), .I2(n1154), .O(n2618) );
  INV_GATE U1945 ( .I1(n2614), .O(n1154) );
  OR_GATE U1946 ( .I1(n8719), .I2(n1155), .O(n8722) );
  INV_GATE U1947 ( .I1(n8720), .O(n1155) );
  OR_GATE U1948 ( .I1(n2550), .I2(n1156), .O(n2553) );
  INV_GATE U1949 ( .I1(n2549), .O(n1156) );
  OR3_GATE U1950 ( .I1(n411), .I2(n1157), .I3(n11840), .O(n12246) );
  AND3_GATE U1951 ( .I1(n11839), .I2(n11838), .I3(n11837), .O(n1157) );
  OR_GATE U1952 ( .I1(n1275), .I2(n1158), .O(n11066) );
  AND_GATE U1953 ( .I1(n11362), .I2(n10908), .O(n1158) );
  OR_GATE U1954 ( .I1(n5879), .I2(n1159), .O(n5882) );
  INV_GATE U1955 ( .I1(n5878), .O(n1159) );
  OR_GATE U1956 ( .I1(n1160), .I2(n5082), .O(n5085) );
  INV_GATE U1957 ( .I1(n5083), .O(n1160) );
  OR_GATE U1958 ( .I1(n5071), .I2(n1161), .O(n5074) );
  INV_GATE U1959 ( .I1(n5072), .O(n1161) );
  OR_GATE U1960 ( .I1(n1162), .I2(n5375), .O(n5378) );
  INV_GATE U1961 ( .I1(n5376), .O(n1162) );
  OR_GATE U1962 ( .I1(n1163), .I2(n5856), .O(n5859) );
  INV_GATE U1963 ( .I1(n5857), .O(n1163) );
  OR_GATE U1964 ( .I1(n1164), .I2(n4200), .O(n4203) );
  INV_GATE U1965 ( .I1(n4201), .O(n1164) );
  OR_GATE U1966 ( .I1(n1165), .I2(n3372), .O(n3375) );
  INV_GATE U1967 ( .I1(n3373), .O(n1165) );
  OR_GATE U1968 ( .I1(n9081), .I2(n1166), .O(n9084) );
  INV_GATE U1969 ( .I1(n9082), .O(n1166) );
  OR_GATE U1970 ( .I1(n1167), .I2(n3361), .O(n3364) );
  INV_GATE U1971 ( .I1(n3362), .O(n1167) );
  OR_GATE U1972 ( .I1(n1168), .I2(n2538), .O(n2541) );
  INV_GATE U1973 ( .I1(n2539), .O(n1168) );
  OR_GATE U1974 ( .I1(n5031), .I2(n1169), .O(n5034) );
  INV_GATE U1975 ( .I1(n5030), .O(n1169) );
  OR_GATE U1976 ( .I1(n9578), .I2(n1170), .O(n9581) );
  INV_GATE U1977 ( .I1(n9579), .O(n1170) );
  OR_GATE U1978 ( .I1(n2528), .I2(n1171), .O(n2531) );
  INV_GATE U1979 ( .I1(n2527), .O(n1171) );
  OR_GATE U1980 ( .I1(n1172), .I2(n4190), .O(n4193) );
  INV_GATE U1981 ( .I1(n4189), .O(n1172) );
  OR_GATE U1982 ( .I1(n9881), .I2(n1173), .O(n9884) );
  INV_GATE U1983 ( .I1(n9882), .O(n1173) );
  OR_GATE U1984 ( .I1(n5020), .I2(n1174), .O(n5023) );
  INV_GATE U1985 ( .I1(n5019), .O(n1174) );
  OR_GATE U1986 ( .I1(n1175), .I2(n3350), .O(n3353) );
  INV_GATE U1987 ( .I1(n3351), .O(n1175) );
  OR_GATE U1988 ( .I1(n10385), .I2(n1176), .O(n10388) );
  INV_GATE U1989 ( .I1(n10386), .O(n1176) );
  OR_GATE U1990 ( .I1(n1177), .I2(n3339), .O(n3342) );
  INV_GATE U1991 ( .I1(n3340), .O(n1177) );
  OR_GATE U1992 ( .I1(n1178), .I2(n4178), .O(n4181) );
  INV_GATE U1993 ( .I1(n4179), .O(n1178) );
  OR_GATE U1994 ( .I1(n10741), .I2(n1179), .O(n10744) );
  INV_GATE U1995 ( .I1(n10742), .O(n1179) );
  OR_GATE U1996 ( .I1(n1180), .I2(n2516), .O(n2519) );
  INV_GATE U1997 ( .I1(n2517), .O(n1180) );
  OR_GATE U1998 ( .I1(n5009), .I2(n1181), .O(n5012) );
  INV_GATE U1999 ( .I1(n5008), .O(n1181) );
  OR_GATE U2000 ( .I1(n1182), .I2(n4167), .O(n4170) );
  INV_GATE U2001 ( .I1(n4168), .O(n1182) );
  OR_GATE U2002 ( .I1(n2506), .I2(n1183), .O(n2509) );
  INV_GATE U2003 ( .I1(n2505), .O(n1183) );
  OR_GATE U2004 ( .I1(n11193), .I2(n1184), .O(n11196) );
  INV_GATE U2005 ( .I1(n11194), .O(n1184) );
  OR_GATE U2006 ( .I1(n1185), .I2(n2494), .O(n2497) );
  INV_GATE U2007 ( .I1(n2495), .O(n1185) );
  OR_GATE U2008 ( .I1(n11590), .I2(n1186), .O(n11593) );
  INV_GATE U2009 ( .I1(n11591), .O(n1186) );
  OR_GATE U2010 ( .I1(n12091), .I2(n1187), .O(n12094) );
  INV_GATE U2011 ( .I1(n12092), .O(n1187) );
  OR_GATE U2012 ( .I1(n1188), .I2(n4156), .O(n4159) );
  INV_GATE U2013 ( .I1(n4157), .O(n1188) );
  OR_GATE U2014 ( .I1(n12478), .I2(n1189), .O(n12481) );
  INV_GATE U2015 ( .I1(n12479), .O(n1189) );
  OR_GATE U2016 ( .I1(n1190), .I2(n4997), .O(n5000) );
  INV_GATE U2017 ( .I1(n4998), .O(n1190) );
  OR_GATE U2018 ( .I1(n12914), .I2(n1191), .O(n12917) );
  INV_GATE U2019 ( .I1(n12915), .O(n1191) );
  OR_GATE U2020 ( .I1(n1192), .I2(n3328), .O(n3331) );
  INV_GATE U2021 ( .I1(n3329), .O(n1192) );
  OR_GATE U2022 ( .I1(n13319), .I2(n1193), .O(n13322) );
  INV_GATE U2023 ( .I1(n13320), .O(n1193) );
  OR_GATE U2024 ( .I1(n2484), .I2(n1194), .O(n2487) );
  INV_GATE U2025 ( .I1(n2483), .O(n1194) );
  OR_GATE U2026 ( .I1(n13753), .I2(n1195), .O(n13756) );
  INV_GATE U2027 ( .I1(n13754), .O(n1195) );
  OR_GATE U2028 ( .I1(n14194), .I2(n1196), .O(n14197) );
  INV_GATE U2029 ( .I1(n14195), .O(n1196) );
  OR_GATE U2030 ( .I1(n4146), .I2(n1197), .O(n4149) );
  INV_GATE U2031 ( .I1(n4145), .O(n1197) );
  OR_GATE U2032 ( .I1(n14804), .I2(n7154), .O(n7151) );
  OR_GATE U2033 ( .I1(n1198), .I2(n2472), .O(n2475) );
  INV_GATE U2034 ( .I1(n2473), .O(n1198) );
  OR_GATE U2035 ( .I1(n4135), .I2(n1199), .O(n4138) );
  INV_GATE U2036 ( .I1(n4134), .O(n1199) );
  OR_GATE U2037 ( .I1(n1200), .I2(n3304), .O(n3307) );
  INV_GATE U2038 ( .I1(n3305), .O(n1200) );
  OR_GATE U2039 ( .I1(n2462), .I2(n1201), .O(n2465) );
  INV_GATE U2040 ( .I1(n2461), .O(n1201) );
  OR_GATE U2041 ( .I1(n1202), .I2(n2792), .O(n2795) );
  INV_GATE U2042 ( .I1(n2793), .O(n1202) );
  OR_GATE U2043 ( .I1(n1203), .I2(n3280), .O(n3283) );
  INV_GATE U2044 ( .I1(n3281), .O(n1203) );
  OR_GATE U2045 ( .I1(n2451), .I2(n1204), .O(n2454) );
  INV_GATE U2046 ( .I1(n2450), .O(n1204) );
  OR_GATE U2047 ( .I1(n1205), .I2(n2439), .O(n2442) );
  INV_GATE U2048 ( .I1(n2440), .O(n1205) );
  OR_GATE U2049 ( .I1(n2429), .I2(n1206), .O(n2432) );
  INV_GATE U2050 ( .I1(n2428), .O(n1206) );
  OR_GATE U2051 ( .I1(n934), .I2(n3884), .O(n3882) );
  OR_GATE U2052 ( .I1(n6193), .I2(n759), .O(n6197) );
  OR_GATE U2053 ( .I1(n4781), .I2(n4785), .O(n4777) );
  OR_GATE U2054 ( .I1(n330), .I2(n5650), .O(n5641) );
  OR_GATE U2055 ( .I1(n326), .I2(n2884), .O(n2934) );
  OR_GATE U2056 ( .I1(n745), .I2(n3735), .O(n3816) );
  OR_GATE U2057 ( .I1(n3775), .I2(n3788), .O(n3794) );
  OR_GATE U2058 ( .I1(n333), .I2(n4322), .O(n4324) );
  OR3_GATE U2059 ( .I1(n1256), .I2(n1207), .I3(n1208), .O(n4425) );
  AND3_GATE U2060 ( .I1(n4372), .I2(n4370), .I3(n4363), .O(n1207) );
  AND_GATE U2061 ( .I1(n4363), .I2(n1216), .O(n1208) );
  AND_GATE U2062 ( .I1(n6173), .I2(n6174), .O(n1209) );
  AND_GATE U2063 ( .I1(n2957), .I2(n2956), .O(n1210) );
  AND_GATE U2064 ( .I1(n2742), .I2(n2739), .O(n1211) );
  OR_GATE U2065 ( .I1(n800), .I2(n5704), .O(n5706) );
  OR_GATE U2066 ( .I1(n619), .I2(n9715), .O(n9716) );
  OR_GATE U2067 ( .I1(n4840), .I2(n4839), .O(n4842) );
  OR_GATE U2068 ( .I1(n801), .I2(n4824), .O(n4826) );
  OR_GATE U2069 ( .I1(n3930), .I2(n3929), .O(n3932) );
  OR_GATE U2070 ( .I1(n3993), .I2(n3992), .O(n3995) );
  OR_GATE U2071 ( .I1(n4922), .I2(n4921), .O(n4924) );
  AND_GATE U2072 ( .I1(n3828), .I2(n3827), .O(n1212) );
  AND_GATE U2073 ( .I1(n2932), .I2(n2931), .O(n1213) );
  OR_GATE U2074 ( .I1(n3028), .I2(n3027), .O(n3030) );
  OR_GATE U2075 ( .I1(n3091), .I2(n3090), .O(n3093) );
  AND_GATE U2076 ( .I1(n4413), .I2(n4412), .O(n1214) );
  OR_GATE U2077 ( .I1(n3107), .I2(n3106), .O(n3109) );
  OR_GATE U2078 ( .I1(n5283), .I2(n5284), .O(n6170) );
  AND_GATE U2079 ( .I1(n3583), .I2(n3581), .O(n1215) );
  AND_GATE U2080 ( .I1(n3806), .I2(n4370), .O(n1216) );
  OR_GATE U2081 ( .I1(n2100), .I2(n2099), .O(n2102) );
  AND_GATE U2082 ( .I1(n4409), .I2(n4626), .O(n1217) );
  OR_GATE U2083 ( .I1(n6142), .I2(n6141), .O(n6136) );
  OR_GATE U2084 ( .I1(n2166), .I2(n2165), .O(n2168) );
  OR_GATE U2085 ( .I1(n6136), .I2(n1304), .O(n6148) );
  OR_GATE U2086 ( .I1(n2199), .I2(n2198), .O(n2201) );
  OR_GATE U2087 ( .I1(n5576), .I2(n6082), .O(n6081) );
  OR_GATE U2088 ( .I1(n5735), .I2(n5734), .O(n5737) );
  OR_GATE U2089 ( .I1(n935), .I2(n5660), .O(n5658) );
  AND_GATE U2090 ( .I1(n5544), .I2(n5540), .O(n1218) );
  OR_GATE U2091 ( .I1(n5751), .I2(n5750), .O(n5753) );
  OR_GATE U2092 ( .I1(n5767), .I2(n5766), .O(n5769) );
  OR_GATE U2093 ( .I1(n5783), .I2(n5782), .O(n5785) );
  OR_GATE U2094 ( .I1(n9471), .I2(n1219), .O(n9467) );
  INV_GATE U2095 ( .I1(n9472), .O(n1219) );
  OR_GATE U2096 ( .I1(n4890), .I2(n4889), .O(n4892) );
  OR_GATE U2097 ( .I1(n3961), .I2(n3960), .O(n3963) );
  OR_GATE U2098 ( .I1(n822), .I2(n3945), .O(n3947) );
  OR_GATE U2099 ( .I1(n3977), .I2(n3976), .O(n3979) );
  AND_GATE U2100 ( .I1(n5333), .I2(n5331), .O(n1220) );
  OR_GATE U2101 ( .I1(n3059), .I2(n3058), .O(n3061) );
  OR_GATE U2102 ( .I1(n4025), .I2(n4024), .O(n4027) );
  OR_GATE U2103 ( .I1(n823), .I2(n3043), .O(n3045) );
  OR_GATE U2104 ( .I1(n3075), .I2(n3074), .O(n3077) );
  AND_GATE U2105 ( .I1(n4709), .I2(n4705), .O(n1221) );
  OR_GATE U2106 ( .I1(n7331), .I2(n7332), .O(n7344) );
  OR_GATE U2107 ( .I1(n2133), .I2(n2132), .O(n2135) );
  OR_GATE U2108 ( .I1(n4872), .I2(n4871), .O(n4874) );
  OR_GATE U2109 ( .I1(n4560), .I2(n4559), .O(n4562) );
  OR_GATE U2110 ( .I1(n4856), .I2(n4855), .O(n4858) );
  AND_GATE U2111 ( .I1(n4726), .I2(n4725), .O(n1222) );
  AND_GATE U2112 ( .I1(n4708), .I2(n4707), .O(n1223) );
  OR_GATE U2113 ( .I1(n4041), .I2(n4040), .O(n4043) );
  OR_GATE U2114 ( .I1(n3139), .I2(n3138), .O(n3141) );
  OR_GATE U2115 ( .I1(n3155), .I2(n3154), .O(n3157) );
  OR_GATE U2116 ( .I1(n403), .I2(n6286), .O(n6287) );
  OR_GATE U2117 ( .I1(n2232), .I2(n2231), .O(n2234) );
  OR_GATE U2118 ( .I1(n5426), .I2(n5425), .O(n5428) );
  OR_GATE U2119 ( .I1(n4954), .I2(n4953), .O(n4956) );
  OR_GATE U2120 ( .I1(n3171), .I2(n3170), .O(n3173) );
  OR_GATE U2121 ( .I1(n5412), .I2(n5411), .O(n5414) );
  OR_GATE U2122 ( .I1(n4970), .I2(n4969), .O(n4972) );
  OR_GATE U2123 ( .I1(n4059), .I2(n4058), .O(n4061) );
  OR_GATE U2124 ( .I1(n3187), .I2(n3186), .O(n3189) );
  OR_GATE U2125 ( .I1(n2265), .I2(n2264), .O(n2267) );
  OR_GATE U2126 ( .I1(n3203), .I2(n3202), .O(n3205) );
  OR_GATE U2127 ( .I1(n2298), .I2(n2297), .O(n2300) );
  OR_GATE U2128 ( .I1(n404), .I2(n8006), .O(n8007) );
  OR_GATE U2129 ( .I1(n4091), .I2(n4090), .O(n4093) );
  OR_GATE U2130 ( .I1(n3219), .I2(n3218), .O(n3221) );
  OR_GATE U2131 ( .I1(n4531), .I2(n4530), .O(n4533) );
  OR_GATE U2132 ( .I1(n415), .I2(n14806), .O(n7153) );
  OR_GATE U2133 ( .I1(n4107), .I2(n4106), .O(n4109) );
  OR_GATE U2134 ( .I1(n2845), .I2(n2844), .O(n2847) );
  OR_GATE U2135 ( .I1(n2331), .I2(n2330), .O(n2333) );
  OR_GATE U2136 ( .I1(n3707), .I2(n3706), .O(n3709) );
  OR_GATE U2137 ( .I1(n3237), .I2(n3236), .O(n3239) );
  OR_GATE U2138 ( .I1(n3693), .I2(n3692), .O(n3695) );
  OR_GATE U2139 ( .I1(n2364), .I2(n2363), .O(n2366) );
  OR_GATE U2140 ( .I1(n2831), .I2(n2830), .O(n2833) );
  OR_GATE U2141 ( .I1(n2817), .I2(n2816), .O(n2819) );
  OR_GATE U2142 ( .I1(n2397), .I2(n2396), .O(n2399) );
  OR_GATE U2143 ( .I1(n1944), .I2(n1943), .O(n1946) );
  OR_GATE U2144 ( .I1(n1255), .I2(n1224), .O(n3874) );
  AND_GATE U2145 ( .I1(n894), .I2(n3629), .O(n1224) );
  OR_GATE U2146 ( .I1(n1225), .I2(n2705), .O(n2706) );
  OR_GATE U2147 ( .I1(n3778), .I2(n3770), .O(n4384) );
  OR_GATE U2148 ( .I1(n3857), .I2(n1226), .O(n3861) );
  AND_GATE U2149 ( .I1(n3858), .I2(n1324), .O(n1226) );
  OR_GATE U2150 ( .I1(n1227), .I2(n6428), .O(n6431) );
  INV_GATE U2151 ( .I1(n6429), .O(n1227) );
  OR3_GATE U2152 ( .I1(n1228), .I2(n1229), .I3(n4603), .O(n5327) );
  INV_GATE U2153 ( .I1(n4607), .O(n1228) );
  AND_GATE U2154 ( .I1(n4602), .I2(n4601), .O(n1229) );
  OR_GATE U2155 ( .I1(n1397), .I2(n2922), .O(n2929) );
  OR_GATE U2156 ( .I1(n4641), .I2(n4646), .O(n5231) );
  OR_GATE U2157 ( .I1(n5537), .I2(n1230), .O(n5253) );
  INV_GATE U2158 ( .I1(n5539), .O(n1230) );
  OR_GATE U2159 ( .I1(n1231), .I2(n7298), .O(n7301) );
  INV_GATE U2160 ( .I1(n7299), .O(n1231) );
  OR_GATE U2161 ( .I1(n1232), .I2(n6108), .O(n6103) );
  INV_GATE U2162 ( .I1(n6105), .O(n1232) );
  OR3_GATE U2163 ( .I1(n4347), .I2(n1233), .I3(n1234), .O(n4702) );
  INV_GATE U2164 ( .I1(n4352), .O(n1233) );
  AND_GATE U2165 ( .I1(n4351), .I2(n4356), .O(n1234) );
  OR3_GATE U2166 ( .I1(n729), .I2(n1235), .I3(n6204), .O(n6217) );
  AND_GATE U2167 ( .I1(n6203), .I2(n6205), .O(n1235) );
  OR_GATE U2168 ( .I1(n5243), .I2(n5240), .O(n5539) );
  OR_GATE U2169 ( .I1(n5294), .I2(n5503), .O(n5505) );
  OR_GATE U2170 ( .I1(n1236), .I2(n7856), .O(n7859) );
  INV_GATE U2171 ( .I1(n7857), .O(n1236) );
  OR_GATE U2172 ( .I1(n8171), .I2(n1237), .O(n8174) );
  INV_GATE U2173 ( .I1(n8172), .O(n1237) );
  OR_GATE U2174 ( .I1(n8704), .I2(n1238), .O(n8707) );
  INV_GATE U2175 ( .I1(n8705), .O(n1238) );
  OR_GATE U2176 ( .I1(n9066), .I2(n1239), .O(n9069) );
  INV_GATE U2177 ( .I1(n9067), .O(n1239) );
  OR_GATE U2178 ( .I1(n9539), .I2(n1240), .O(n9542) );
  INV_GATE U2179 ( .I1(n9540), .O(n1240) );
  OR_GATE U2180 ( .I1(n9906), .I2(n1241), .O(n9909) );
  INV_GATE U2181 ( .I1(n9907), .O(n1241) );
  OR_GATE U2182 ( .I1(n10410), .I2(n1242), .O(n10413) );
  INV_GATE U2183 ( .I1(n10411), .O(n1242) );
  OR_GATE U2184 ( .I1(n10766), .I2(n1243), .O(n10769) );
  INV_GATE U2185 ( .I1(n10767), .O(n1243) );
  OR_GATE U2186 ( .I1(n11218), .I2(n1244), .O(n11221) );
  INV_GATE U2187 ( .I1(n11219), .O(n1244) );
  OR_GATE U2188 ( .I1(n11615), .I2(n1245), .O(n11618) );
  INV_GATE U2189 ( .I1(n11616), .O(n1245) );
  OR_GATE U2190 ( .I1(n12116), .I2(n1246), .O(n12119) );
  INV_GATE U2191 ( .I1(n12117), .O(n1246) );
  OR_GATE U2192 ( .I1(n12503), .I2(n1247), .O(n12506) );
  INV_GATE U2193 ( .I1(n12504), .O(n1247) );
  OR_GATE U2194 ( .I1(n12939), .I2(n1248), .O(n12942) );
  INV_GATE U2195 ( .I1(n12940), .O(n1248) );
  OR_GATE U2196 ( .I1(n13344), .I2(n1249), .O(n13347) );
  INV_GATE U2197 ( .I1(n13345), .O(n1249) );
  OR_GATE U2198 ( .I1(n13778), .I2(n1250), .O(n13781) );
  INV_GATE U2199 ( .I1(n13779), .O(n1250) );
  OR_GATE U2200 ( .I1(n14219), .I2(n1251), .O(n14222) );
  INV_GATE U2201 ( .I1(n14220), .O(n1251) );
  OR_GATE U2202 ( .I1(n2423), .I2(n409), .O(n14783) );
  OR_GATE U2203 ( .I1(n1937), .I2(n410), .O(n14782) );
  OR_GATE U2204 ( .I1(n8681), .I2(n8680), .O(n8683) );
  OR_GATE U2205 ( .I1(n9043), .I2(n9042), .O(n9045) );
  OR_GATE U2206 ( .I1(n9551), .I2(n9550), .O(n9553) );
  OR_GATE U2207 ( .I1(n9918), .I2(n9917), .O(n9920) );
  OR_GATE U2208 ( .I1(n10422), .I2(n10421), .O(n10424) );
  OR_GATE U2209 ( .I1(n10778), .I2(n10777), .O(n10780) );
  OR_GATE U2210 ( .I1(n5404), .I2(n405), .O(n5406) );
  OR_GATE U2211 ( .I1(n11230), .I2(n11229), .O(n11232) );
  OR_GATE U2212 ( .I1(n11627), .I2(n11626), .O(n11629) );
  OR_GATE U2213 ( .I1(n12128), .I2(n12127), .O(n12130) );
  OR_GATE U2214 ( .I1(n12515), .I2(n12514), .O(n12517) );
  OR_GATE U2215 ( .I1(n12951), .I2(n12950), .O(n12953) );
  OR_GATE U2216 ( .I1(n406), .I2(n4523), .O(n4524) );
  OR_GATE U2217 ( .I1(n3685), .I2(n407), .O(n3687) );
  OR_GATE U2218 ( .I1(n408), .I2(n2809), .O(n2810) );
  AND_GATE U2219 ( .I1(A[1]), .I2(n1401), .O(n1252) );
  OR_GATE U2220 ( .I1(n2028), .I2(n2025), .O(n2700) );
  OR_GATE U2221 ( .I1(A[0]), .I2(n1253), .O(n2025) );
  AND_GATE U2222 ( .I1(n1400), .I2(n1864), .O(n1253) );
  AND_GATE U2223 ( .I1(A[0]), .I2(A[1]), .O(n1254) );
  NOR_GATE U2224 ( .I1(n3858), .I2(n3857), .O(n1255) );
  AND_GATE U2225 ( .I1(n3806), .I2(n4372), .O(n1256) );
  OR_GATE U2226 ( .I1(n9428), .I2(n8923), .O(n8922) );
  OR_GATE U2227 ( .I1(n932), .I2(n1257), .O(n2712) );
  AND_GATE U2228 ( .I1(n1441), .I2(A[1]), .O(n1257) );
  OR_GATE U2229 ( .I1(n10922), .I2(n1147), .O(n10931) );
  OR_GATE U2230 ( .I1(n7735), .I2(n7734), .O(n7736) );
  OR_GATE U2231 ( .I1(n6221), .I2(n796), .O(n6223) );
  AND_GATE U2232 ( .I1(n5586), .I2(n5585), .O(n1258) );
  OR_GATE U2233 ( .I1(n11905), .I2(n1259), .O(n11910) );
  AND_GATE U2234 ( .I1(n11907), .I2(n11906), .O(n1259) );
  OR_GATE U2235 ( .I1(n483), .I2(n12611), .O(n1261) );
  AND_GATE U2236 ( .I1(n12615), .I2(n12614), .O(n1262) );
  AND_GATE U2237 ( .I1(n10976), .I2(n10975), .O(n1263) );
  AND_GATE U2238 ( .I1(n3512), .I2(n3511), .O(n1264) );
  NAND_GATE U2239 ( .I1(n2870), .I2(n2747), .O(n1265) );
  AND_GATE U2240 ( .I1(n3853), .I2(n3852), .O(n1266) );
  AND_GATE U2241 ( .I1(n2972), .I2(n2971), .O(n1267) );
  NOR_GATE U2242 ( .I1(n3741), .I2(n3819), .O(n1268) );
  OR_GATE U2243 ( .I1(n303), .I2(n4339), .O(n4441) );
  NOR_GATE U2244 ( .I1(n2735), .I2(n2736), .O(n1269) );
  INV_GATE U2245 ( .I1(n1269), .O(n2740) );
  OR_GATE U2246 ( .I1(n2946), .I2(n2941), .O(n2954) );
  OR_GATE U2247 ( .I1(n1270), .I2(n14487), .O(n14491) );
  AND_GATE U2248 ( .I1(n14286), .I2(n14503), .O(n1270) );
  OR_GATE U2249 ( .I1(n280), .I2(n12645), .O(n12646) );
  OR_GATE U2250 ( .I1(n5621), .I2(n782), .O(n5623) );
  AND_GATE U2251 ( .I1(n10597), .I2(n10596), .O(n1271) );
  NOR_GATE U2252 ( .I1(n1365), .I2(n1273), .O(n1272) );
  OR_GATE U2253 ( .I1(n1365), .I2(n1273), .O(n6956) );
  AND_GATE U2254 ( .I1(n7039), .I2(n6478), .O(n1273) );
  OR_GATE U2255 ( .I1(n4797), .I2(n4796), .O(n4798) );
  OR_GATE U2256 ( .I1(n11796), .I2(n350), .O(n11798) );
  OR_GATE U2257 ( .I1(n9618), .I2(n664), .O(n9620) );
  OR_GATE U2258 ( .I1(n13922), .I2(n1274), .O(n13929) );
  INV_GATE U2259 ( .I1(n13930), .O(n1274) );
  NOR_GATE U2260 ( .I1(n11355), .I2(n11357), .O(n1275) );
  OR_GATE U2261 ( .I1(n13518), .I2(n13516), .O(n13522) );
  INV_GATE U2262 ( .I1(n1276), .O(n9421) );
  OR_GATE U2263 ( .I1(n7206), .I2(n1277), .O(n7210) );
  INV_GATE U2264 ( .I1(n7207), .O(n1277) );
  AND3_GATE U2265 ( .I1(n11758), .I2(n11757), .I3(n11756), .O(n1278) );
  INV_GATE U2266 ( .I1(n1278), .O(n11869) );
  OR_GATE U2267 ( .I1(n362), .I2(n9462), .O(n9461) );
  OR_GATE U2268 ( .I1(n932), .I2(n1279), .O(n2021) );
  AND_GATE U2269 ( .I1(n1442), .I2(A[1]), .O(n1279) );
  AND_GATE U2270 ( .I1(n3831), .I2(n3837), .O(n1280) );
  NAND_GATE U2271 ( .I1(n2716), .I2(n2717), .O(n1281) );
  OR_GATE U2272 ( .I1(n2982), .I2(n1391), .O(n2987) );
  OR_GATE U2273 ( .I1(n2970), .I2(n1371), .O(n2971) );
  OR_GATE U2274 ( .I1(n8637), .I2(n8636), .O(n8640) );
  AND3_GATE U2275 ( .I1(n13025), .I2(n13433), .I3(n13432), .O(n1282) );
  INV_GATE U2276 ( .I1(n1282), .O(n13147) );
  OR3_GATE U2277 ( .I1(n4709), .I2(n4705), .I3(n1301), .O(n4707) );
  OR3_GATE U2278 ( .I1(n2930), .I2(n2922), .I3(n1397), .O(n2931) );
  AND3_GATE U2279 ( .I1(n8068), .I2(n7974), .I3(n8067), .O(n1283) );
  NOR_GATE U2280 ( .I1(n10119), .I2(n10121), .O(n1284) );
  AND3_GATE U2281 ( .I1(n6074), .I2(n5605), .I3(n6073), .O(n1285) );
  INV_GATE U2282 ( .I1(n1285), .O(n6055) );
  NAND_GATE U2283 ( .I1(n8633), .I2(n1288), .O(n1286) );
  AND_GATE U2284 ( .I1(n1286), .I2(n1287), .O(n8758) );
  OR_GATE U2285 ( .I1(n8632), .I2(n8628), .O(n1287) );
  AND_GATE U2286 ( .I1(n8627), .I2(n8757), .O(n1288) );
  OR_GATE U2287 ( .I1(n7791), .I2(n7790), .O(n7789) );
  NOR_GATE U2288 ( .I1(n8320), .I2(n8322), .O(n1289) );
  AND3_GATE U2289 ( .I1(n7100), .I2(n7216), .I3(n7217), .O(n1290) );
  AND3_GATE U2290 ( .I1(n6101), .I2(n6100), .I3(n6099), .O(n1291) );
  INV_GATE U2291 ( .I1(n1291), .O(n6484) );
  OR_GATE U2292 ( .I1(n1291), .I2(n6482), .O(n6485) );
  NAND_GATE U2293 ( .I1(n7260), .I2(n1295), .O(n1292) );
  AND_GATE U2294 ( .I1(n1292), .I2(n1293), .O(n7266) );
  OR_GATE U2295 ( .I1(n1294), .I2(n7263), .O(n1293) );
  INV_GATE U2296 ( .I1(n7264), .O(n1294) );
  AND_GATE U2297 ( .I1(n7261), .I2(n7264), .O(n1295) );
  AND_GATE U2298 ( .I1(n4674), .I2(n4675), .O(n1296) );
  AND_GATE U2299 ( .I1(n8244), .I2(n8243), .O(n1297) );
  AND_GATE U2300 ( .I1(n7047), .I2(n7046), .O(n1298) );
  OR_GATE U2301 ( .I1(n1973), .I2(n1972), .O(n1975) );
  OR_GATE U2302 ( .I1(n1299), .I2(n10279), .O(n10276) );
  INV_GATE U2303 ( .I1(n10274), .O(n1299) );
  OR_GATE U2304 ( .I1(n6192), .I2(n7), .O(n6382) );
  OR_GATE U2305 ( .I1(n6168), .I2(n1322), .O(n5515) );
  OR_GATE U2306 ( .I1(n9977), .I2(n1300), .O(n9980) );
  INV_GATE U2307 ( .I1(n9978), .O(n1300) );
  OR_GATE U2308 ( .I1(n647), .I2(n11424), .O(n11426) );
  AND3_GATE U2309 ( .I1(n4701), .I2(n4702), .I3(n4700), .O(n1301) );
  NOR_GATE U2310 ( .I1(n10571), .I2(n1302), .O(\A2[40] ) );
  INV_GATE U2311 ( .I1(n1323), .O(n1302) );
  AND_GATE U2312 ( .I1(n4446), .I2(n4445), .O(n1303) );
  OR_GATE U2313 ( .I1(n764), .I2(n5312), .O(n5307) );
  OR_GATE U2314 ( .I1(n6142), .I2(n1304), .O(n6139) );
  INV_GATE U2315 ( .I1(n6138), .O(n1304) );
  NAND_GATE U2316 ( .I1(n13034), .I2(n1307), .O(n1305) );
  AND_GATE U2317 ( .I1(n1305), .I2(n1306), .O(n13036) );
  OR_GATE U2318 ( .I1(n13031), .I2(n13030), .O(n1306) );
  AND_GATE U2319 ( .I1(n13033), .I2(n13035), .O(n1307) );
  NAND_GATE U2320 ( .I1(n1308), .I2(n7872), .O(n7870) );
  NOR_GATE U2321 ( .I1(n7874), .I2(n7873), .O(n1308) );
  NAND_GATE U2322 ( .I1(n1309), .I2(n6981), .O(n6979) );
  NOR_GATE U2323 ( .I1(n6983), .I2(n6982), .O(n1309) );
  AND3_GATE U2324 ( .I1(n9974), .I2(n9616), .I3(n9973), .O(n1310) );
  AND_GATE U2325 ( .I1(n9009), .I2(n9008), .O(n1311) );
  NAND_GATE U2326 ( .I1(n8125), .I2(n1314), .O(n1312) );
  AND_GATE U2327 ( .I1(n1312), .I2(n1313), .O(n8730) );
  OR_GATE U2328 ( .I1(n8735), .I2(n8128), .O(n1313) );
  AND_GATE U2329 ( .I1(n8126), .I2(n8193), .O(n1314) );
  AND_GATE U2330 ( .I1(n7344), .I2(n7343), .O(n1315) );
  AND_GATE U2331 ( .I1(n6456), .I2(n6455), .O(n1316) );
  AND_GATE U2332 ( .I1(n8635), .I2(n8209), .O(n1317) );
  INV_GATE U2333 ( .I1(n1317), .O(n8750) );
  OR_GATE U2334 ( .I1(n9158), .I2(n1318), .O(n9160) );
  INV_GATE U2335 ( .I1(n9157), .O(n1318) );
  OR_GATE U2336 ( .I1(n1319), .I2(n7290), .O(n7285) );
  INV_GATE U2337 ( .I1(n7287), .O(n1319) );
  NOR_GATE U2338 ( .I1(n1323), .I2(n1321), .O(n1320) );
  AND_GATE U2339 ( .I1(n10574), .I2(n927), .O(n1321) );
  OR_GATE U2340 ( .I1(n322), .I2(n3486), .O(n3489) );
  OR3_GATE U2341 ( .I1(n6168), .I2(n6172), .I3(n1322), .O(n6174) );
  INV_GATE U2342 ( .I1(n5514), .O(n1322) );
  OR_GATE U2343 ( .I1(n8982), .I2(n802), .O(n8983) );
  NOR_GATE U2344 ( .I1(n10574), .I2(n927), .O(n1323) );
  AND_GATE U2345 ( .I1(n3849), .I2(n3628), .O(n1324) );
  OR_GATE U2346 ( .I1(n2870), .I2(n1375), .O(n2879) );
  NAND_GATE U2347 ( .I1(n2998), .I2(n1327), .O(n1325) );
  AND_GATE U2348 ( .I1(n1325), .I2(n1326), .O(n3002) );
  OR_GATE U2349 ( .I1(n2995), .I2(n3000), .O(n1326) );
  AND_GATE U2350 ( .I1(n2999), .I2(n3001), .O(n1327) );
  NAND_GATE U2351 ( .I1(n1328), .I2(n8491), .O(n8490) );
  NOR_GATE U2352 ( .I1(n8493), .I2(n8492), .O(n1328) );
  NAND_GATE U2353 ( .I1(n1329), .I2(n7674), .O(n7673) );
  NOR_GATE U2354 ( .I1(n7676), .I2(n7675), .O(n1329) );
  NAND_GATE U2355 ( .I1(n1330), .I2(n6252), .O(n6251) );
  NOR_GATE U2356 ( .I1(n6254), .I2(n6253), .O(n1330) );
  AND_GATE U2357 ( .I1(n9323), .I2(n9322), .O(n1331) );
  AND_GATE U2358 ( .I1(n3880), .I2(n3633), .O(n1332) );
  NAND_GATE U2359 ( .I1(n9285), .I2(n1335), .O(n1333) );
  AND_GATE U2360 ( .I1(n1333), .I2(n1334), .O(n9312) );
  OR_GATE U2361 ( .I1(n9319), .I2(n9287), .O(n1334) );
  AND_GATE U2362 ( .I1(n9286), .I2(n9288), .O(n1335) );
  OR_GATE U2363 ( .I1(n1337), .I2(n9330), .O(n9325) );
  INV_GATE U2364 ( .I1(n9327), .O(n1337) );
  AND_GATE U2365 ( .I1(n3626), .I2(n3625), .O(n1338) );
  OR_GATE U2366 ( .I1(n10956), .I2(n10960), .O(n10957) );
  AND_GATE U2367 ( .I1(n2716), .I2(n2717), .O(n1339) );
  OR_GATE U2368 ( .I1(n8922), .I2(n1017), .O(n9423) );
  NAND_GATE U2369 ( .I1(n11706), .I2(n1342), .O(n1340) );
  AND_GATE U2370 ( .I1(n1340), .I2(n1341), .O(n11708) );
  AND_GATE U2371 ( .I1(n11705), .I2(n11707), .O(n1342) );
  NAND_GATE U2372 ( .I1(n5545), .I2(n1218), .O(n5543) );
  NAND_GATE U2373 ( .I1(n7051), .I2(n1345), .O(n1343) );
  OR_GATE U2374 ( .I1(n7047), .I2(n7046), .O(n1344) );
  AND_GATE U2375 ( .I1(n7050), .I2(n7261), .O(n1345) );
  AND3_GATE U2376 ( .I1(n7269), .I2(n7055), .I3(n7054), .O(n1346) );
  OR_GATE U2377 ( .I1(n793), .I2(n7771), .O(n7764) );
  OR_GATE U2378 ( .I1(n7381), .I2(n7382), .O(n7386) );
  OR_GATE U2379 ( .I1(n5287), .I2(n5290), .O(n5286) );
  AND_GATE U2380 ( .I1(n7066), .I2(n7065), .O(n1347) );
  INV_GATE U2381 ( .I1(n1347), .O(n7073) );
  OR_GATE U2382 ( .I1(n2914), .I2(n1348), .O(n3564) );
  INV_GATE U2383 ( .I1(n3556), .O(n1348) );
  OR_GATE U2384 ( .I1(n5165), .I2(n5166), .O(n5168) );
  AND_GATE U2385 ( .I1(n4575), .I2(n4475), .O(n1349) );
  INV_GATE U2386 ( .I1(n1349), .O(n4780) );
  NAND_GATE U2387 ( .I1(n7350), .I2(n1352), .O(n1350) );
  AND_GATE U2388 ( .I1(n1350), .I2(n1351), .O(n7355) );
  OR_GATE U2389 ( .I1(n7349), .I2(n7353), .O(n1351) );
  AND_GATE U2390 ( .I1(n7358), .I2(n7354), .O(n1352) );
  AND_GATE U2391 ( .I1(n5250), .I2(n5249), .O(n1354) );
  AND_GATE U2392 ( .I1(n2883), .I2(n2882), .O(n1355) );
  INV_GATE U2393 ( .I1(n1355), .O(n3602) );
  OR_GATE U2394 ( .I1(n11411), .I2(n1390), .O(n11413) );
  OR_GATE U2395 ( .I1(n10170), .I2(n10171), .O(n10173) );
  NOR_GATE U2396 ( .I1(n11850), .I2(n11851), .O(n1356) );
  NAND_GATE U2397 ( .I1(n293), .I2(n1359), .O(n1357) );
  AND_GATE U2398 ( .I1(n7956), .I2(n7957), .O(n1359) );
  AND_GATE U2399 ( .I1(n1360), .I2(n1361), .O(n6929) );
  AND_GATE U2400 ( .I1(n8078), .I2(n8074), .O(n1362) );
  OR_GATE U2401 ( .I1(n9672), .I2(n9674), .O(n9780) );
  OR_GATE U2402 ( .I1(n5544), .I2(n5545), .O(n5547) );
  OR_GATE U2403 ( .I1(n8588), .I2(n1363), .O(n8846) );
  INV_GATE U2404 ( .I1(n8589), .O(n1363) );
  OR_GATE U2405 ( .I1(n13527), .I2(n614), .O(n13529) );
  OR_GATE U2406 ( .I1(n2856), .I2(n1398), .O(n2858) );
  INV_GATE U2407 ( .I1(n6969), .O(n1364) );
  OR_GATE U2408 ( .I1(n12702), .I2(n12704), .O(n12701) );
  NOR_GATE U2409 ( .I1(n7030), .I2(n7031), .O(n1365) );
  OR_GATE U2410 ( .I1(n1366), .I2(n10637), .O(n10639) );
  INV_GATE U2411 ( .I1(n10638), .O(n1366) );
  OR_GATE U2412 ( .I1(n10058), .I2(n10059), .O(n10061) );
  OR_GATE U2413 ( .I1(n264), .I2(n12599), .O(n12706) );
  OR_GATE U2414 ( .I1(n169), .I2(n10182), .O(n10184) );
  NAND_GATE U2415 ( .I1(n1367), .I2(n13992), .O(n13991) );
  NOR_GATE U2416 ( .I1(n13993), .I2(n13994), .O(n1367) );
  NAND_GATE U2417 ( .I1(n14450), .I2(n14319), .O(n1368) );
  AND_GATE U2418 ( .I1(n14474), .I2(n14491), .O(n1369) );
  AND_GATE U2419 ( .I1(n5557), .I2(n5556), .O(n1370) );
  OR_GATE U2420 ( .I1(n4781), .I2(n1349), .O(n4783) );
  AND_GATE U2421 ( .I1(n2870), .I2(n2747), .O(n1371) );
  AND3_GATE U2422 ( .I1(n2706), .I2(n2707), .I3(n2708), .O(n1372) );
  INV_GATE U2423 ( .I1(n1372), .O(n2924) );
  OR_GATE U2424 ( .I1(n10981), .I2(n10980), .O(n10983) );
  OR_GATE U2425 ( .I1(n1373), .I2(n1855), .O(n1857) );
  INV_GATE U2426 ( .I1(n1856), .O(n1373) );
  NOR_GATE U2427 ( .I1(n11900), .I2(n11901), .O(n1374) );
  AND_GATE U2428 ( .I1(n2946), .I2(n2746), .O(n1375) );
  INV_GATE U2429 ( .I1(n1375), .O(n2871) );
  NAND_GATE U2430 ( .I1(n1382), .I2(n1378), .O(n1376) );
  AND_GATE U2431 ( .I1(n1376), .I2(n1377), .O(n6316) );
  NAND_GATE U2432 ( .I1(n895), .I2(n1381), .O(n1379) );
  AND_GATE U2433 ( .I1(n1379), .I2(n1380), .O(n3872) );
  OR_GATE U2434 ( .I1(n3870), .I2(n3866), .O(n1380) );
  AND_GATE U2435 ( .I1(n3868), .I2(n3867), .O(n1381) );
  AND_GATE U2436 ( .I1(n5984), .I2(n5983), .O(n1382) );
  NOR_GATE U2437 ( .I1(n11905), .I2(n11907), .O(n1383) );
  AND_GATE U2438 ( .I1(n5598), .I2(n6209), .O(n1384) );
  AND_GATE U2439 ( .I1(n10919), .I2(n10918), .O(n1385) );
  OR_GATE U2440 ( .I1(n388), .I2(n5290), .O(n5503) );
  OR_GATE U2441 ( .I1(n7395), .I2(n7396), .O(n7944) );
  AND3_GATE U2442 ( .I1(n8280), .I2(n8279), .I3(n8814), .O(n1386) );
  OR_GATE U2443 ( .I1(n294), .I2(n7239), .O(n7234) );
  AND3_GATE U2444 ( .I1(n13070), .I2(n13069), .I3(n13068), .O(n1387) );
  INV_GATE U2445 ( .I1(n1387), .O(n13523) );
  AND_GATE U2446 ( .I1(n14450), .I2(n14319), .O(n1388) );
  AND_GATE U2447 ( .I1(n10914), .I2(n10913), .O(n1389) );
  OR_GATE U2448 ( .I1(n5989), .I2(n5990), .O(n5992) );
  OR_GATE U2449 ( .I1(n869), .I2(n12648), .O(n12633) );
  OR_GATE U2450 ( .I1(n14382), .I2(n14826), .O(n14378) );
  NOR_GATE U2451 ( .I1(n2984), .I2(n2983), .O(n1391) );
  AND_GATE U2452 ( .I1(n8093), .I2(n8092), .O(n1392) );
  AND3_GATE U2453 ( .I1(n10293), .I2(n10038), .I3(n10292), .O(n1393) );
  INV_GATE U2454 ( .I1(n1393), .O(n10286) );
  OR_GATE U2455 ( .I1(n8745), .I2(n1317), .O(n8747) );
  OR_GATE U2456 ( .I1(n1394), .I2(n4314), .O(n4308) );
  INV_GATE U2457 ( .I1(n4311), .O(n1394) );
  INV_GATE U2458 ( .I1(n1395), .O(n11888) );
  AND_GATE U2459 ( .I1(n6521), .I2(n6916), .O(n1396) );
  OR_GATE U2460 ( .I1(n11868), .I2(n1278), .O(n12274) );
  NOR_GATE U2461 ( .I1(n2709), .I2(n1372), .O(n1397) );
  OR_GATE U2462 ( .I1(n7889), .I2(n7888), .O(n7891) );
  NOR_GATE U2463 ( .I1(n2854), .I2(n2862), .O(n1398) );
  NOR_GATE U2464 ( .I1(n13921), .I2(n13922), .O(n1399) );
  OR_GATE U2465 ( .I1(n13925), .I2(n727), .O(n13922) );
  INV_GATE U2466 ( .I1(n1402), .O(n1401) );
  INV_GATE U2467 ( .I1(B[0]), .O(n1402) );
  INV_GATE U2468 ( .I1(B[1]), .O(n1403) );
  INV_GATE U2469 ( .I1(n1406), .O(n1404) );
  INV_GATE U2470 ( .I1(n1406), .O(n1405) );
  INV_GATE U2471 ( .I1(B[2]), .O(n1406) );
  INV_GATE U2472 ( .I1(B[3]), .O(n1407) );
  INV_GATE U2473 ( .I1(B[4]), .O(n1408) );
  INV_GATE U2474 ( .I1(n1411), .O(n1409) );
  INV_GATE U2475 ( .I1(n1411), .O(n1410) );
  INV_GATE U2476 ( .I1(B[5]), .O(n1411) );
  INV_GATE U2477 ( .I1(B[6]), .O(n1412) );
  INV_GATE U2478 ( .I1(n1414), .O(n1413) );
  INV_GATE U2479 ( .I1(B[7]), .O(n1414) );
  INV_GATE U2480 ( .I1(n1417), .O(n1415) );
  INV_GATE U2481 ( .I1(n1417), .O(n1416) );
  INV_GATE U2482 ( .I1(B[8]), .O(n1417) );
  INV_GATE U2483 ( .I1(n1419), .O(n1418) );
  INV_GATE U2484 ( .I1(B[9]), .O(n1419) );
  INV_GATE U2485 ( .I1(B[10]), .O(n1420) );
  INV_GATE U2486 ( .I1(B[11]), .O(n1421) );
  INV_GATE U2487 ( .I1(n1423), .O(n1422) );
  INV_GATE U2488 ( .I1(B[12]), .O(n1423) );
  INV_GATE U2489 ( .I1(B[13]), .O(n1424) );
  INV_GATE U2490 ( .I1(n1426), .O(n1425) );
  INV_GATE U2491 ( .I1(B[14]), .O(n1426) );
  INV_GATE U2492 ( .I1(B[15]), .O(n1427) );
  INV_GATE U2493 ( .I1(B[16]), .O(n1428) );
  INV_GATE U2494 ( .I1(B[17]), .O(n1429) );
  INV_GATE U2495 ( .I1(B[18]), .O(n1430) );
  INV_GATE U2496 ( .I1(B[19]), .O(n1431) );
  INV_GATE U2497 ( .I1(B[20]), .O(n1432) );
  INV_GATE U2498 ( .I1(B[21]), .O(n1433) );
  INV_GATE U2499 ( .I1(B[22]), .O(n1434) );
  INV_GATE U2500 ( .I1(B[23]), .O(n1435) );
  INV_GATE U2501 ( .I1(B[24]), .O(n1436) );
  INV_GATE U2502 ( .I1(B[25]), .O(n1437) );
  INV_GATE U2503 ( .I1(B[26]), .O(n1438) );
  INV_GATE U2504 ( .I1(B[27]), .O(n1439) );
  INV_GATE U2505 ( .I1(B[28]), .O(n1440) );
  INV_GATE U2506 ( .I1(B[29]), .O(n1441) );
  INV_GATE U2507 ( .I1(B[30]), .O(n1442) );
  INV_GATE U2508 ( .I1(B[31]), .O(n1443) );
  INV_GATE U2509 ( .I1(A[0]), .O(n1444) );
  INV_GATE U2510 ( .I1(A[1]), .O(n1445) );
  INV_GATE U2511 ( .I1(A[2]), .O(n1446) );
  INV_GATE U2512 ( .I1(A[3]), .O(n1447) );
  INV_GATE U2513 ( .I1(A[4]), .O(n1448) );
  INV_GATE U2514 ( .I1(A[5]), .O(n1449) );
  INV_GATE U2515 ( .I1(A[6]), .O(n1450) );
  INV_GATE U2516 ( .I1(A[7]), .O(n1451) );
  INV_GATE U2517 ( .I1(A[8]), .O(n1452) );
  INV_GATE U2518 ( .I1(A[9]), .O(n1453) );
  INV_GATE U2519 ( .I1(A[10]), .O(n1454) );
  INV_GATE U2520 ( .I1(A[11]), .O(n1455) );
  INV_GATE U2521 ( .I1(A[12]), .O(n1456) );
  INV_GATE U2522 ( .I1(A[13]), .O(n1457) );
  INV_GATE U2523 ( .I1(A[14]), .O(n1458) );
  INV_GATE U2524 ( .I1(A[15]), .O(n1459) );
  INV_GATE U2525 ( .I1(A[16]), .O(n1460) );
  INV_GATE U2526 ( .I1(A[17]), .O(n1461) );
  INV_GATE U2527 ( .I1(A[18]), .O(n1462) );
  INV_GATE U2528 ( .I1(A[19]), .O(n1463) );
  INV_GATE U2529 ( .I1(A[20]), .O(n1464) );
  INV_GATE U2530 ( .I1(A[21]), .O(n1465) );
  INV_GATE U2531 ( .I1(A[22]), .O(n1466) );
  INV_GATE U2532 ( .I1(A[23]), .O(n1467) );
  INV_GATE U2533 ( .I1(A[24]), .O(n1468) );
  INV_GATE U2534 ( .I1(A[25]), .O(n1469) );
  INV_GATE U2535 ( .I1(A[26]), .O(n1470) );
  INV_GATE U2536 ( .I1(A[27]), .O(n1471) );
  INV_GATE U2537 ( .I1(A[28]), .O(n1472) );
  INV_GATE U2538 ( .I1(A[29]), .O(n1473) );
  INV_GATE U2539 ( .I1(A[30]), .O(n1474) );
  INV_GATE U2540 ( .I1(A[31]), .O(n1475) );
  NAND_GATE U2541 ( .I1(n14839), .I2(n1252), .O(n1477) );
  OR_GATE U2542 ( .I1(n1252), .I2(n14839), .O(n1476) );
  NAND_GATE U2543 ( .I1(n1477), .I2(n1476), .O(PRODUCT[1]) );
  OR_GATE U2544 ( .I1(A[31]), .I2(B[31]), .O(\A1[61] ) );
  NAND_GATE U2545 ( .I1(B[31]), .I2(A[31]), .O(n14829) );
  OR_GATE U2546 ( .I1(n14829), .I2(A[30]), .O(n1481) );
  NAND_GATE U2547 ( .I1(B[31]), .I2(n1475), .O(n1479) );
  NAND_GATE U2548 ( .I1(n1443), .I2(A[31]), .O(n1478) );
  NAND_GATE U2549 ( .I1(n1479), .I2(n1478), .O(n14384) );
  INV_GATE U2550 ( .I1(n14384), .O(n14386) );
  NAND_GATE U2551 ( .I1(n14829), .I2(n14386), .O(n1480) );
  NAND_GATE U2552 ( .I1(n1481), .I2(n1480), .O(n1482) );
  NAND_GATE U2553 ( .I1(B[30]), .I2(B[31]), .O(n1483) );
  NAND_GATE U2554 ( .I1(n1482), .I2(n1483), .O(\A1[60] ) );
  INV_GATE U2555 ( .I1(n1483), .O(n1929) );
  NAND3_GATE U2556 ( .I1(n1929), .I2(n1472), .I3(A[29]), .O(n1539) );
  NAND_GATE U2557 ( .I1(A[29]), .I2(B[30]), .O(n1550) );
  NAND3_GATE U2558 ( .I1(n1929), .I2(n1470), .I3(A[27]), .O(n1535) );
  NAND_GATE U2559 ( .I1(A[27]), .I2(B[30]), .O(n1573) );
  NAND3_GATE U2560 ( .I1(n1929), .I2(n1468), .I3(A[25]), .O(n1531) );
  NAND_GATE U2561 ( .I1(A[25]), .I2(B[30]), .O(n1596) );
  NAND3_GATE U2562 ( .I1(n1929), .I2(n1466), .I3(A[23]), .O(n1527) );
  NAND_GATE U2563 ( .I1(A[23]), .I2(B[30]), .O(n1619) );
  NAND3_GATE U2564 ( .I1(n1929), .I2(n1464), .I3(A[21]), .O(n1523) );
  NAND_GATE U2565 ( .I1(A[21]), .I2(B[30]), .O(n1642) );
  NAND3_GATE U2566 ( .I1(n1929), .I2(n1462), .I3(A[19]), .O(n1519) );
  NAND_GATE U2567 ( .I1(A[19]), .I2(B[30]), .O(n1665) );
  NAND3_GATE U2568 ( .I1(n1929), .I2(n1460), .I3(A[17]), .O(n1515) );
  NAND_GATE U2569 ( .I1(A[17]), .I2(B[30]), .O(n1688) );
  NAND3_GATE U2570 ( .I1(n1929), .I2(n1458), .I3(A[15]), .O(n1511) );
  NAND_GATE U2571 ( .I1(A[15]), .I2(B[30]), .O(n1711) );
  NAND3_GATE U2572 ( .I1(n1929), .I2(n1456), .I3(A[13]), .O(n1507) );
  NAND_GATE U2573 ( .I1(A[13]), .I2(B[30]), .O(n1734) );
  NAND3_GATE U2574 ( .I1(n1929), .I2(n1454), .I3(A[11]), .O(n1503) );
  NAND_GATE U2575 ( .I1(A[11]), .I2(B[30]), .O(n1757) );
  NAND3_GATE U2576 ( .I1(n1929), .I2(n1452), .I3(A[9]), .O(n1499) );
  NAND_GATE U2577 ( .I1(A[9]), .I2(B[30]), .O(n1780) );
  NAND3_GATE U2578 ( .I1(n1929), .I2(n1450), .I3(A[7]), .O(n1495) );
  NAND_GATE U2579 ( .I1(A[7]), .I2(B[30]), .O(n1803) );
  NAND3_GATE U2580 ( .I1(n1929), .I2(n1448), .I3(A[5]), .O(n1491) );
  NAND_GATE U2581 ( .I1(A[5]), .I2(B[30]), .O(n1826) );
  NAND3_GATE U2582 ( .I1(A[3]), .I2(n1929), .I3(n1446), .O(n1487) );
  INV_GATE U2583 ( .I1(n1850), .O(n1485) );
  NAND3_GATE U2584 ( .I1(n932), .I2(n1929), .I3(A[2]), .O(n1863) );
  NAND3_GATE U2585 ( .I1(A[2]), .I2(n1445), .I3(n1929), .O(n1484) );
  NAND_GATE U2586 ( .I1(n1863), .I2(n1484), .O(n1856) );
  NAND_GATE U2587 ( .I1(n1485), .I2(n1856), .O(n1486) );
  NAND_GATE U2588 ( .I1(n1447), .I2(n1929), .O(n1488) );
  NAND_GATE U2589 ( .I1(n301), .I2(n1488), .O(n1489) );
  NAND_GATE U2590 ( .I1(A[4]), .I2(n1489), .O(n1834) );
  OR_GATE U2591 ( .I1(n1826), .I2(n1834), .O(n1490) );
  NAND_GATE U2592 ( .I1(n1491), .I2(n1490), .O(n1822) );
  NAND_GATE U2593 ( .I1(n1449), .I2(n1929), .O(n1492) );
  NAND_GATE U2594 ( .I1(n1819), .I2(n1492), .O(n1493) );
  NAND_GATE U2595 ( .I1(A[6]), .I2(n1493), .O(n1811) );
  OR_GATE U2596 ( .I1(n1803), .I2(n1811), .O(n1494) );
  NAND_GATE U2597 ( .I1(n1495), .I2(n1494), .O(n1799) );
  NAND_GATE U2598 ( .I1(n1451), .I2(n1929), .O(n1496) );
  NAND_GATE U2599 ( .I1(n1796), .I2(n1496), .O(n1497) );
  NAND_GATE U2600 ( .I1(A[8]), .I2(n1497), .O(n1788) );
  OR_GATE U2601 ( .I1(n1780), .I2(n1788), .O(n1498) );
  NAND_GATE U2602 ( .I1(n1499), .I2(n1498), .O(n1776) );
  INV_GATE U2603 ( .I1(n1776), .O(n1773) );
  NAND_GATE U2604 ( .I1(n1453), .I2(n1929), .O(n1500) );
  NAND_GATE U2605 ( .I1(n1773), .I2(n1500), .O(n1501) );
  NAND_GATE U2606 ( .I1(A[10]), .I2(n1501), .O(n1765) );
  OR_GATE U2607 ( .I1(n1757), .I2(n1765), .O(n1502) );
  NAND_GATE U2608 ( .I1(n1503), .I2(n1502), .O(n1753) );
  INV_GATE U2609 ( .I1(n1753), .O(n1750) );
  NAND_GATE U2610 ( .I1(n1455), .I2(n1929), .O(n1504) );
  NAND_GATE U2611 ( .I1(n1750), .I2(n1504), .O(n1505) );
  NAND_GATE U2612 ( .I1(A[12]), .I2(n1505), .O(n1742) );
  OR_GATE U2613 ( .I1(n1734), .I2(n1742), .O(n1506) );
  NAND_GATE U2614 ( .I1(n1507), .I2(n1506), .O(n1730) );
  INV_GATE U2615 ( .I1(n1730), .O(n1727) );
  NAND_GATE U2616 ( .I1(n1457), .I2(n1929), .O(n1508) );
  NAND_GATE U2617 ( .I1(n1727), .I2(n1508), .O(n1509) );
  NAND_GATE U2618 ( .I1(A[14]), .I2(n1509), .O(n1719) );
  OR_GATE U2619 ( .I1(n1711), .I2(n1719), .O(n1510) );
  NAND_GATE U2620 ( .I1(n1511), .I2(n1510), .O(n1707) );
  INV_GATE U2621 ( .I1(n1707), .O(n1704) );
  NAND_GATE U2622 ( .I1(n1459), .I2(n1929), .O(n1512) );
  NAND_GATE U2623 ( .I1(n1704), .I2(n1512), .O(n1513) );
  NAND_GATE U2624 ( .I1(A[16]), .I2(n1513), .O(n1696) );
  OR_GATE U2625 ( .I1(n1688), .I2(n1696), .O(n1514) );
  NAND_GATE U2626 ( .I1(n1515), .I2(n1514), .O(n1684) );
  INV_GATE U2627 ( .I1(n1684), .O(n1681) );
  NAND_GATE U2628 ( .I1(n1461), .I2(n1929), .O(n1516) );
  NAND_GATE U2629 ( .I1(n1681), .I2(n1516), .O(n1517) );
  NAND_GATE U2630 ( .I1(A[18]), .I2(n1517), .O(n1673) );
  OR_GATE U2631 ( .I1(n1665), .I2(n1673), .O(n1518) );
  NAND_GATE U2632 ( .I1(n1519), .I2(n1518), .O(n1661) );
  INV_GATE U2633 ( .I1(n1661), .O(n1658) );
  NAND_GATE U2634 ( .I1(n1463), .I2(n1929), .O(n1520) );
  NAND_GATE U2635 ( .I1(n1658), .I2(n1520), .O(n1521) );
  NAND_GATE U2636 ( .I1(A[20]), .I2(n1521), .O(n1650) );
  OR_GATE U2637 ( .I1(n1642), .I2(n1650), .O(n1522) );
  NAND_GATE U2638 ( .I1(n1523), .I2(n1522), .O(n1638) );
  INV_GATE U2639 ( .I1(n1638), .O(n1635) );
  NAND_GATE U2640 ( .I1(n1465), .I2(n1929), .O(n1524) );
  NAND_GATE U2641 ( .I1(n1635), .I2(n1524), .O(n1525) );
  NAND_GATE U2642 ( .I1(A[22]), .I2(n1525), .O(n1627) );
  OR_GATE U2643 ( .I1(n1619), .I2(n1627), .O(n1526) );
  NAND_GATE U2644 ( .I1(n1527), .I2(n1526), .O(n1615) );
  INV_GATE U2645 ( .I1(n1615), .O(n1612) );
  NAND_GATE U2646 ( .I1(n1467), .I2(n1929), .O(n1528) );
  NAND_GATE U2647 ( .I1(n1612), .I2(n1528), .O(n1529) );
  NAND_GATE U2648 ( .I1(A[24]), .I2(n1529), .O(n1604) );
  OR_GATE U2649 ( .I1(n1596), .I2(n1604), .O(n1530) );
  NAND_GATE U2650 ( .I1(n1531), .I2(n1530), .O(n1592) );
  INV_GATE U2651 ( .I1(n1592), .O(n1589) );
  NAND_GATE U2652 ( .I1(n1469), .I2(n1929), .O(n1532) );
  NAND_GATE U2653 ( .I1(n1589), .I2(n1532), .O(n1533) );
  NAND_GATE U2654 ( .I1(A[26]), .I2(n1533), .O(n1581) );
  OR_GATE U2655 ( .I1(n1573), .I2(n1581), .O(n1534) );
  NAND_GATE U2656 ( .I1(n1535), .I2(n1534), .O(n1569) );
  INV_GATE U2657 ( .I1(n1569), .O(n1566) );
  NAND_GATE U2658 ( .I1(n1471), .I2(n1929), .O(n1536) );
  NAND_GATE U2659 ( .I1(n1566), .I2(n1536), .O(n1537) );
  NAND_GATE U2660 ( .I1(A[28]), .I2(n1537), .O(n1558) );
  OR_GATE U2661 ( .I1(n1550), .I2(n1558), .O(n1538) );
  NAND_GATE U2662 ( .I1(n1539), .I2(n1538), .O(n1546) );
  INV_GATE U2663 ( .I1(n1546), .O(n1936) );
  NAND_GATE U2664 ( .I1(B[30]), .I2(n1443), .O(n1837) );
  NAND_GATE U2665 ( .I1(n1550), .I2(n1837), .O(n1540) );
  NAND_GATE U2666 ( .I1(A[30]), .I2(n1540), .O(n1543) );
  NAND_GATE U2667 ( .I1(n1474), .I2(B[31]), .O(n1930) );
  NAND_GATE U2668 ( .I1(n1400), .I2(n1930), .O(n1541) );
  NAND_GATE U2669 ( .I1(n1473), .I2(n1541), .O(n1542) );
  NAND_GATE U2670 ( .I1(n1543), .I2(n1542), .O(n1544) );
  NAND_GATE U2671 ( .I1(n1936), .I2(n1544), .O(n1548) );
  INV_GATE U2672 ( .I1(n1544), .O(n1545) );
  NAND_GATE U2673 ( .I1(n1546), .I2(n1545), .O(n1547) );
  NAND_GATE U2674 ( .I1(n1548), .I2(n1547), .O(n2412) );
  NAND_GATE U2675 ( .I1(B[29]), .I2(A[30]), .O(n1948) );
  INV_GATE U2676 ( .I1(n1948), .O(n1942) );
  INV_GATE U2677 ( .I1(n1558), .O(n1555) );
  INV_GATE U2678 ( .I1(n1837), .O(n1848) );
  NAND_GATE U2679 ( .I1(A[29]), .I2(n1848), .O(n1554) );
  NAND_GATE U2680 ( .I1(n1473), .I2(B[31]), .O(n1549) );
  NAND3_GATE U2681 ( .I1(n1472), .I2(n1400), .I3(n1549), .O(n1552) );
  NAND_GATE U2682 ( .I1(A[28]), .I2(n1550), .O(n1551) );
  NAND_GATE U2683 ( .I1(n1552), .I2(n1551), .O(n1553) );
  NAND_GATE U2684 ( .I1(n1554), .I2(n1553), .O(n1556) );
  NAND_GATE U2685 ( .I1(n1555), .I2(n1556), .O(n1560) );
  INV_GATE U2686 ( .I1(n1556), .O(n1557) );
  NAND_GATE U2687 ( .I1(n1558), .I2(n1557), .O(n1559) );
  NAND_GATE U2688 ( .I1(n1560), .I2(n1559), .O(n1941) );
  INV_GATE U2689 ( .I1(n1941), .O(n1944) );
  NAND_GATE U2690 ( .I1(n1942), .I2(n1944), .O(n1939) );
  NAND_GATE U2691 ( .I1(B[29]), .I2(A[29]), .O(n1963) );
  INV_GATE U2692 ( .I1(n1963), .O(n1956) );
  NAND_GATE U2693 ( .I1(n1573), .I2(n1837), .O(n1561) );
  NAND_GATE U2694 ( .I1(A[28]), .I2(n1561), .O(n1565) );
  NAND_GATE U2695 ( .I1(n1472), .I2(B[31]), .O(n1562) );
  NAND_GATE U2696 ( .I1(n1400), .I2(n1562), .O(n1563) );
  NAND_GATE U2697 ( .I1(n1471), .I2(n1563), .O(n1564) );
  NAND_GATE U2698 ( .I1(n1565), .I2(n1564), .O(n1567) );
  NAND_GATE U2699 ( .I1(n1566), .I2(n1567), .O(n1571) );
  INV_GATE U2700 ( .I1(n1567), .O(n1568) );
  NAND_GATE U2701 ( .I1(n1569), .I2(n1568), .O(n1570) );
  NAND_GATE U2702 ( .I1(n1571), .I2(n1570), .O(n1958) );
  NAND_GATE U2703 ( .I1(n1956), .I2(n1958), .O(n1953) );
  NAND_GATE U2704 ( .I1(B[29]), .I2(A[28]), .O(n2401) );
  INV_GATE U2705 ( .I1(n2401), .O(n2395) );
  INV_GATE U2706 ( .I1(n1581), .O(n1578) );
  NAND_GATE U2707 ( .I1(A[27]), .I2(n1848), .O(n1577) );
  NAND_GATE U2708 ( .I1(n1471), .I2(B[31]), .O(n1572) );
  NAND3_GATE U2709 ( .I1(n1470), .I2(n1400), .I3(n1572), .O(n1575) );
  NAND_GATE U2710 ( .I1(A[26]), .I2(n1573), .O(n1574) );
  NAND_GATE U2711 ( .I1(n1575), .I2(n1574), .O(n1576) );
  NAND_GATE U2712 ( .I1(n1577), .I2(n1576), .O(n1579) );
  NAND_GATE U2713 ( .I1(n1578), .I2(n1579), .O(n1583) );
  INV_GATE U2714 ( .I1(n1579), .O(n1580) );
  NAND_GATE U2715 ( .I1(n1581), .I2(n1580), .O(n1582) );
  NAND_GATE U2716 ( .I1(n1583), .I2(n1582), .O(n2394) );
  INV_GATE U2717 ( .I1(n2394), .O(n2397) );
  NAND_GATE U2718 ( .I1(n2395), .I2(n2397), .O(n2392) );
  NAND_GATE U2719 ( .I1(B[29]), .I2(A[27]), .O(n2385) );
  INV_GATE U2720 ( .I1(n2385), .O(n2378) );
  NAND_GATE U2721 ( .I1(n1596), .I2(n1837), .O(n1584) );
  NAND_GATE U2722 ( .I1(A[26]), .I2(n1584), .O(n1588) );
  NAND_GATE U2723 ( .I1(n1470), .I2(B[31]), .O(n1585) );
  NAND_GATE U2724 ( .I1(n1400), .I2(n1585), .O(n1586) );
  NAND_GATE U2725 ( .I1(n1469), .I2(n1586), .O(n1587) );
  NAND_GATE U2726 ( .I1(n1588), .I2(n1587), .O(n1590) );
  NAND_GATE U2727 ( .I1(n1589), .I2(n1590), .O(n1594) );
  INV_GATE U2728 ( .I1(n1590), .O(n1591) );
  NAND_GATE U2729 ( .I1(n1592), .I2(n1591), .O(n1593) );
  NAND_GATE U2730 ( .I1(n1594), .I2(n1593), .O(n2380) );
  NAND_GATE U2731 ( .I1(n2378), .I2(n2380), .O(n2375) );
  NAND_GATE U2732 ( .I1(B[29]), .I2(A[26]), .O(n2368) );
  INV_GATE U2733 ( .I1(n2368), .O(n2362) );
  INV_GATE U2734 ( .I1(n1604), .O(n1601) );
  NAND_GATE U2735 ( .I1(A[25]), .I2(n1848), .O(n1600) );
  NAND_GATE U2736 ( .I1(n1469), .I2(B[31]), .O(n1595) );
  NAND3_GATE U2737 ( .I1(n1468), .I2(n1400), .I3(n1595), .O(n1598) );
  NAND_GATE U2738 ( .I1(A[24]), .I2(n1596), .O(n1597) );
  NAND_GATE U2739 ( .I1(n1598), .I2(n1597), .O(n1599) );
  NAND_GATE U2740 ( .I1(n1600), .I2(n1599), .O(n1602) );
  NAND_GATE U2741 ( .I1(n1601), .I2(n1602), .O(n1606) );
  INV_GATE U2742 ( .I1(n1602), .O(n1603) );
  NAND_GATE U2743 ( .I1(n1604), .I2(n1603), .O(n1605) );
  NAND_GATE U2744 ( .I1(n1606), .I2(n1605), .O(n2361) );
  INV_GATE U2745 ( .I1(n2361), .O(n2364) );
  NAND_GATE U2746 ( .I1(n2362), .I2(n2364), .O(n2359) );
  NAND_GATE U2747 ( .I1(B[29]), .I2(A[25]), .O(n2352) );
  INV_GATE U2748 ( .I1(n2352), .O(n2345) );
  NAND_GATE U2749 ( .I1(n1619), .I2(n1837), .O(n1607) );
  NAND_GATE U2750 ( .I1(A[24]), .I2(n1607), .O(n1611) );
  NAND_GATE U2751 ( .I1(n1468), .I2(B[31]), .O(n1608) );
  NAND_GATE U2752 ( .I1(n1400), .I2(n1608), .O(n1609) );
  NAND_GATE U2753 ( .I1(n1467), .I2(n1609), .O(n1610) );
  NAND_GATE U2754 ( .I1(n1611), .I2(n1610), .O(n1613) );
  NAND_GATE U2755 ( .I1(n1612), .I2(n1613), .O(n1617) );
  INV_GATE U2756 ( .I1(n1613), .O(n1614) );
  NAND_GATE U2757 ( .I1(n1615), .I2(n1614), .O(n1616) );
  NAND_GATE U2758 ( .I1(n1617), .I2(n1616), .O(n2347) );
  NAND_GATE U2759 ( .I1(n2345), .I2(n2347), .O(n2342) );
  NAND_GATE U2760 ( .I1(B[29]), .I2(A[24]), .O(n2335) );
  INV_GATE U2761 ( .I1(n2335), .O(n2329) );
  INV_GATE U2762 ( .I1(n1627), .O(n1624) );
  NAND_GATE U2763 ( .I1(A[23]), .I2(n1848), .O(n1623) );
  NAND_GATE U2764 ( .I1(n1467), .I2(B[31]), .O(n1618) );
  NAND3_GATE U2765 ( .I1(n1466), .I2(n1400), .I3(n1618), .O(n1621) );
  NAND_GATE U2766 ( .I1(A[22]), .I2(n1619), .O(n1620) );
  NAND_GATE U2767 ( .I1(n1621), .I2(n1620), .O(n1622) );
  NAND_GATE U2768 ( .I1(n1623), .I2(n1622), .O(n1625) );
  NAND_GATE U2769 ( .I1(n1624), .I2(n1625), .O(n1629) );
  INV_GATE U2770 ( .I1(n1625), .O(n1626) );
  NAND_GATE U2771 ( .I1(n1627), .I2(n1626), .O(n1628) );
  NAND_GATE U2772 ( .I1(n1629), .I2(n1628), .O(n2328) );
  INV_GATE U2773 ( .I1(n2328), .O(n2331) );
  NAND_GATE U2774 ( .I1(n2329), .I2(n2331), .O(n2326) );
  NAND_GATE U2775 ( .I1(B[29]), .I2(A[23]), .O(n2319) );
  INV_GATE U2776 ( .I1(n2319), .O(n2312) );
  NAND_GATE U2777 ( .I1(n1642), .I2(n1837), .O(n1630) );
  NAND_GATE U2778 ( .I1(A[22]), .I2(n1630), .O(n1634) );
  NAND_GATE U2779 ( .I1(n1466), .I2(B[31]), .O(n1631) );
  NAND_GATE U2780 ( .I1(n1400), .I2(n1631), .O(n1632) );
  NAND_GATE U2781 ( .I1(n1465), .I2(n1632), .O(n1633) );
  NAND_GATE U2782 ( .I1(n1634), .I2(n1633), .O(n1636) );
  NAND_GATE U2783 ( .I1(n1635), .I2(n1636), .O(n1640) );
  INV_GATE U2784 ( .I1(n1636), .O(n1637) );
  NAND_GATE U2785 ( .I1(n1638), .I2(n1637), .O(n1639) );
  NAND_GATE U2786 ( .I1(n1640), .I2(n1639), .O(n2314) );
  NAND_GATE U2787 ( .I1(n2312), .I2(n2314), .O(n2309) );
  NAND_GATE U2788 ( .I1(B[29]), .I2(A[22]), .O(n2302) );
  INV_GATE U2789 ( .I1(n2302), .O(n2296) );
  INV_GATE U2790 ( .I1(n1650), .O(n1647) );
  NAND_GATE U2791 ( .I1(A[21]), .I2(n1848), .O(n1646) );
  NAND_GATE U2792 ( .I1(n1465), .I2(B[31]), .O(n1641) );
  NAND3_GATE U2793 ( .I1(n1464), .I2(n1400), .I3(n1641), .O(n1644) );
  NAND_GATE U2794 ( .I1(A[20]), .I2(n1642), .O(n1643) );
  NAND_GATE U2795 ( .I1(n1644), .I2(n1643), .O(n1645) );
  NAND_GATE U2796 ( .I1(n1646), .I2(n1645), .O(n1648) );
  NAND_GATE U2797 ( .I1(n1647), .I2(n1648), .O(n1652) );
  INV_GATE U2798 ( .I1(n1648), .O(n1649) );
  NAND_GATE U2799 ( .I1(n1650), .I2(n1649), .O(n1651) );
  NAND_GATE U2800 ( .I1(n1652), .I2(n1651), .O(n2295) );
  INV_GATE U2801 ( .I1(n2295), .O(n2298) );
  NAND_GATE U2802 ( .I1(n2296), .I2(n2298), .O(n2293) );
  NAND_GATE U2803 ( .I1(B[29]), .I2(A[21]), .O(n2286) );
  INV_GATE U2804 ( .I1(n2286), .O(n2279) );
  NAND_GATE U2805 ( .I1(n1665), .I2(n1837), .O(n1653) );
  NAND_GATE U2806 ( .I1(A[20]), .I2(n1653), .O(n1657) );
  NAND_GATE U2807 ( .I1(n1464), .I2(B[31]), .O(n1654) );
  NAND_GATE U2808 ( .I1(n1400), .I2(n1654), .O(n1655) );
  NAND_GATE U2809 ( .I1(n1463), .I2(n1655), .O(n1656) );
  NAND_GATE U2810 ( .I1(n1657), .I2(n1656), .O(n1659) );
  NAND_GATE U2811 ( .I1(n1658), .I2(n1659), .O(n1663) );
  INV_GATE U2812 ( .I1(n1659), .O(n1660) );
  NAND_GATE U2813 ( .I1(n1661), .I2(n1660), .O(n1662) );
  NAND_GATE U2814 ( .I1(n1663), .I2(n1662), .O(n2281) );
  NAND_GATE U2815 ( .I1(n2279), .I2(n2281), .O(n2276) );
  NAND_GATE U2816 ( .I1(B[29]), .I2(A[20]), .O(n2269) );
  INV_GATE U2817 ( .I1(n2269), .O(n2263) );
  INV_GATE U2818 ( .I1(n1673), .O(n1670) );
  NAND_GATE U2819 ( .I1(A[19]), .I2(n1848), .O(n1669) );
  NAND_GATE U2820 ( .I1(n1463), .I2(B[31]), .O(n1664) );
  NAND3_GATE U2821 ( .I1(n1462), .I2(n1400), .I3(n1664), .O(n1667) );
  NAND_GATE U2822 ( .I1(A[18]), .I2(n1665), .O(n1666) );
  NAND_GATE U2823 ( .I1(n1667), .I2(n1666), .O(n1668) );
  NAND_GATE U2824 ( .I1(n1669), .I2(n1668), .O(n1671) );
  NAND_GATE U2825 ( .I1(n1670), .I2(n1671), .O(n1675) );
  INV_GATE U2826 ( .I1(n1671), .O(n1672) );
  NAND_GATE U2827 ( .I1(n1673), .I2(n1672), .O(n1674) );
  NAND_GATE U2828 ( .I1(n1675), .I2(n1674), .O(n2262) );
  INV_GATE U2829 ( .I1(n2262), .O(n2265) );
  NAND_GATE U2830 ( .I1(n2263), .I2(n2265), .O(n2260) );
  NAND_GATE U2831 ( .I1(B[29]), .I2(A[19]), .O(n2253) );
  INV_GATE U2832 ( .I1(n2253), .O(n2246) );
  NAND_GATE U2833 ( .I1(n1688), .I2(n1837), .O(n1676) );
  NAND_GATE U2834 ( .I1(A[18]), .I2(n1676), .O(n1680) );
  NAND_GATE U2835 ( .I1(n1462), .I2(B[31]), .O(n1677) );
  NAND_GATE U2836 ( .I1(n1400), .I2(n1677), .O(n1678) );
  NAND_GATE U2837 ( .I1(n1461), .I2(n1678), .O(n1679) );
  NAND_GATE U2838 ( .I1(n1680), .I2(n1679), .O(n1682) );
  NAND_GATE U2839 ( .I1(n1681), .I2(n1682), .O(n1686) );
  INV_GATE U2840 ( .I1(n1682), .O(n1683) );
  NAND_GATE U2841 ( .I1(n1684), .I2(n1683), .O(n1685) );
  NAND_GATE U2842 ( .I1(n1686), .I2(n1685), .O(n2248) );
  NAND_GATE U2843 ( .I1(n2246), .I2(n2248), .O(n2243) );
  NAND_GATE U2844 ( .I1(B[29]), .I2(A[18]), .O(n2236) );
  INV_GATE U2845 ( .I1(n2236), .O(n2230) );
  INV_GATE U2846 ( .I1(n1696), .O(n1693) );
  NAND_GATE U2847 ( .I1(A[17]), .I2(n1848), .O(n1692) );
  NAND_GATE U2848 ( .I1(n1461), .I2(B[31]), .O(n1687) );
  NAND3_GATE U2849 ( .I1(n1460), .I2(n1400), .I3(n1687), .O(n1690) );
  NAND_GATE U2850 ( .I1(A[16]), .I2(n1688), .O(n1689) );
  NAND_GATE U2851 ( .I1(n1690), .I2(n1689), .O(n1691) );
  NAND_GATE U2852 ( .I1(n1692), .I2(n1691), .O(n1694) );
  NAND_GATE U2853 ( .I1(n1693), .I2(n1694), .O(n1698) );
  INV_GATE U2854 ( .I1(n1694), .O(n1695) );
  NAND_GATE U2855 ( .I1(n1696), .I2(n1695), .O(n1697) );
  NAND_GATE U2856 ( .I1(n1698), .I2(n1697), .O(n2229) );
  INV_GATE U2857 ( .I1(n2229), .O(n2232) );
  NAND_GATE U2858 ( .I1(n2230), .I2(n2232), .O(n2227) );
  NAND_GATE U2859 ( .I1(B[29]), .I2(A[17]), .O(n2220) );
  INV_GATE U2860 ( .I1(n2220), .O(n2213) );
  NAND_GATE U2861 ( .I1(n1711), .I2(n1837), .O(n1699) );
  NAND_GATE U2862 ( .I1(A[16]), .I2(n1699), .O(n1703) );
  NAND_GATE U2863 ( .I1(n1460), .I2(B[31]), .O(n1700) );
  NAND_GATE U2864 ( .I1(n1400), .I2(n1700), .O(n1701) );
  NAND_GATE U2865 ( .I1(n1459), .I2(n1701), .O(n1702) );
  NAND_GATE U2866 ( .I1(n1703), .I2(n1702), .O(n1705) );
  NAND_GATE U2867 ( .I1(n1704), .I2(n1705), .O(n1709) );
  INV_GATE U2868 ( .I1(n1705), .O(n1706) );
  NAND_GATE U2869 ( .I1(n1707), .I2(n1706), .O(n1708) );
  NAND_GATE U2870 ( .I1(n1709), .I2(n1708), .O(n2215) );
  NAND_GATE U2871 ( .I1(n2213), .I2(n2215), .O(n2210) );
  NAND_GATE U2872 ( .I1(B[29]), .I2(A[16]), .O(n2203) );
  INV_GATE U2873 ( .I1(n2203), .O(n2197) );
  INV_GATE U2874 ( .I1(n1719), .O(n1716) );
  NAND_GATE U2875 ( .I1(A[15]), .I2(n1848), .O(n1715) );
  NAND_GATE U2876 ( .I1(n1459), .I2(B[31]), .O(n1710) );
  NAND3_GATE U2877 ( .I1(n1458), .I2(n1400), .I3(n1710), .O(n1713) );
  NAND_GATE U2878 ( .I1(A[14]), .I2(n1711), .O(n1712) );
  NAND_GATE U2879 ( .I1(n1713), .I2(n1712), .O(n1714) );
  NAND_GATE U2880 ( .I1(n1715), .I2(n1714), .O(n1717) );
  NAND_GATE U2881 ( .I1(n1716), .I2(n1717), .O(n1721) );
  INV_GATE U2882 ( .I1(n1717), .O(n1718) );
  NAND_GATE U2883 ( .I1(n1719), .I2(n1718), .O(n1720) );
  NAND_GATE U2884 ( .I1(n1721), .I2(n1720), .O(n2196) );
  INV_GATE U2885 ( .I1(n2196), .O(n2199) );
  NAND_GATE U2886 ( .I1(n2197), .I2(n2199), .O(n2194) );
  NAND_GATE U2887 ( .I1(B[29]), .I2(A[15]), .O(n2187) );
  INV_GATE U2888 ( .I1(n2187), .O(n2180) );
  NAND_GATE U2889 ( .I1(n1734), .I2(n1837), .O(n1722) );
  NAND_GATE U2890 ( .I1(A[14]), .I2(n1722), .O(n1726) );
  NAND_GATE U2891 ( .I1(n1458), .I2(B[31]), .O(n1723) );
  NAND_GATE U2892 ( .I1(n1400), .I2(n1723), .O(n1724) );
  NAND_GATE U2893 ( .I1(n1457), .I2(n1724), .O(n1725) );
  NAND_GATE U2894 ( .I1(n1726), .I2(n1725), .O(n1728) );
  NAND_GATE U2895 ( .I1(n1727), .I2(n1728), .O(n1732) );
  INV_GATE U2896 ( .I1(n1728), .O(n1729) );
  NAND_GATE U2897 ( .I1(n1730), .I2(n1729), .O(n1731) );
  NAND_GATE U2898 ( .I1(n1732), .I2(n1731), .O(n2182) );
  NAND_GATE U2899 ( .I1(n2180), .I2(n2182), .O(n2177) );
  NAND_GATE U2900 ( .I1(B[29]), .I2(A[14]), .O(n2170) );
  INV_GATE U2901 ( .I1(n2170), .O(n2164) );
  INV_GATE U2902 ( .I1(n1742), .O(n1739) );
  NAND_GATE U2903 ( .I1(A[13]), .I2(n1848), .O(n1738) );
  NAND_GATE U2904 ( .I1(n1457), .I2(B[31]), .O(n1733) );
  NAND3_GATE U2905 ( .I1(n1456), .I2(n1400), .I3(n1733), .O(n1736) );
  NAND_GATE U2906 ( .I1(A[12]), .I2(n1734), .O(n1735) );
  NAND_GATE U2907 ( .I1(n1736), .I2(n1735), .O(n1737) );
  NAND_GATE U2908 ( .I1(n1738), .I2(n1737), .O(n1740) );
  NAND_GATE U2909 ( .I1(n1739), .I2(n1740), .O(n1744) );
  INV_GATE U2910 ( .I1(n1740), .O(n1741) );
  NAND_GATE U2911 ( .I1(n1742), .I2(n1741), .O(n1743) );
  NAND_GATE U2912 ( .I1(n1744), .I2(n1743), .O(n2163) );
  INV_GATE U2913 ( .I1(n2163), .O(n2166) );
  NAND_GATE U2914 ( .I1(n2164), .I2(n2166), .O(n2161) );
  NAND_GATE U2915 ( .I1(B[29]), .I2(A[13]), .O(n2154) );
  INV_GATE U2916 ( .I1(n2154), .O(n2147) );
  NAND_GATE U2917 ( .I1(n1757), .I2(n1837), .O(n1745) );
  NAND_GATE U2918 ( .I1(A[12]), .I2(n1745), .O(n1749) );
  NAND_GATE U2919 ( .I1(n1456), .I2(B[31]), .O(n1746) );
  NAND_GATE U2920 ( .I1(n1400), .I2(n1746), .O(n1747) );
  NAND_GATE U2921 ( .I1(n1455), .I2(n1747), .O(n1748) );
  NAND_GATE U2922 ( .I1(n1749), .I2(n1748), .O(n1751) );
  NAND_GATE U2923 ( .I1(n1750), .I2(n1751), .O(n1755) );
  INV_GATE U2924 ( .I1(n1751), .O(n1752) );
  NAND_GATE U2925 ( .I1(n1753), .I2(n1752), .O(n1754) );
  NAND_GATE U2926 ( .I1(n1755), .I2(n1754), .O(n2149) );
  NAND_GATE U2927 ( .I1(n2147), .I2(n2149), .O(n2144) );
  NAND_GATE U2928 ( .I1(B[29]), .I2(A[12]), .O(n2137) );
  INV_GATE U2929 ( .I1(n2137), .O(n2131) );
  INV_GATE U2930 ( .I1(n1765), .O(n1762) );
  NAND_GATE U2931 ( .I1(A[11]), .I2(n1848), .O(n1761) );
  NAND_GATE U2932 ( .I1(n1455), .I2(B[31]), .O(n1756) );
  NAND3_GATE U2933 ( .I1(n1454), .I2(n1400), .I3(n1756), .O(n1759) );
  NAND_GATE U2934 ( .I1(A[10]), .I2(n1757), .O(n1758) );
  NAND_GATE U2935 ( .I1(n1759), .I2(n1758), .O(n1760) );
  NAND_GATE U2936 ( .I1(n1761), .I2(n1760), .O(n1763) );
  NAND_GATE U2937 ( .I1(n1762), .I2(n1763), .O(n1767) );
  INV_GATE U2938 ( .I1(n1763), .O(n1764) );
  NAND_GATE U2939 ( .I1(n1765), .I2(n1764), .O(n1766) );
  NAND_GATE U2940 ( .I1(n1767), .I2(n1766), .O(n2130) );
  INV_GATE U2941 ( .I1(n2130), .O(n2133) );
  NAND_GATE U2942 ( .I1(n2131), .I2(n2133), .O(n2128) );
  NAND_GATE U2943 ( .I1(B[29]), .I2(A[11]), .O(n2121) );
  INV_GATE U2944 ( .I1(n2121), .O(n2114) );
  NAND_GATE U2945 ( .I1(n1780), .I2(n1837), .O(n1768) );
  NAND_GATE U2946 ( .I1(A[10]), .I2(n1768), .O(n1772) );
  NAND_GATE U2947 ( .I1(n1454), .I2(B[31]), .O(n1769) );
  NAND_GATE U2948 ( .I1(n1400), .I2(n1769), .O(n1770) );
  NAND_GATE U2949 ( .I1(n1453), .I2(n1770), .O(n1771) );
  NAND_GATE U2950 ( .I1(n1772), .I2(n1771), .O(n1774) );
  NAND_GATE U2951 ( .I1(n1773), .I2(n1774), .O(n1778) );
  INV_GATE U2952 ( .I1(n1774), .O(n1775) );
  NAND_GATE U2953 ( .I1(n1776), .I2(n1775), .O(n1777) );
  NAND_GATE U2954 ( .I1(n1778), .I2(n1777), .O(n2116) );
  NAND_GATE U2955 ( .I1(n2114), .I2(n2116), .O(n2111) );
  NAND_GATE U2956 ( .I1(B[29]), .I2(A[10]), .O(n2104) );
  INV_GATE U2957 ( .I1(n2104), .O(n2098) );
  INV_GATE U2958 ( .I1(n1788), .O(n1785) );
  NAND_GATE U2959 ( .I1(A[9]), .I2(n1848), .O(n1784) );
  NAND_GATE U2960 ( .I1(n1453), .I2(B[31]), .O(n1779) );
  NAND3_GATE U2961 ( .I1(n1452), .I2(n1400), .I3(n1779), .O(n1782) );
  NAND_GATE U2962 ( .I1(A[8]), .I2(n1780), .O(n1781) );
  NAND_GATE U2963 ( .I1(n1782), .I2(n1781), .O(n1783) );
  NAND_GATE U2964 ( .I1(n1784), .I2(n1783), .O(n1786) );
  NAND_GATE U2965 ( .I1(n1785), .I2(n1786), .O(n1790) );
  INV_GATE U2966 ( .I1(n1786), .O(n1787) );
  NAND_GATE U2967 ( .I1(n1788), .I2(n1787), .O(n1789) );
  NAND_GATE U2968 ( .I1(n1790), .I2(n1789), .O(n2097) );
  INV_GATE U2969 ( .I1(n2097), .O(n2100) );
  NAND_GATE U2970 ( .I1(n2098), .I2(n2100), .O(n2095) );
  NAND_GATE U2971 ( .I1(B[29]), .I2(A[9]), .O(n2088) );
  INV_GATE U2972 ( .I1(n2088), .O(n2081) );
  NAND_GATE U2973 ( .I1(n1803), .I2(n1837), .O(n1791) );
  NAND_GATE U2974 ( .I1(A[8]), .I2(n1791), .O(n1795) );
  NAND_GATE U2975 ( .I1(n1452), .I2(B[31]), .O(n1792) );
  NAND_GATE U2976 ( .I1(n1400), .I2(n1792), .O(n1793) );
  NAND_GATE U2977 ( .I1(n1451), .I2(n1793), .O(n1794) );
  NAND_GATE U2978 ( .I1(n1795), .I2(n1794), .O(n1797) );
  NAND_GATE U2979 ( .I1(n1796), .I2(n1797), .O(n1801) );
  INV_GATE U2980 ( .I1(n1797), .O(n1798) );
  NAND_GATE U2981 ( .I1(n1799), .I2(n1798), .O(n1800) );
  NAND_GATE U2982 ( .I1(n1801), .I2(n1800), .O(n2083) );
  NAND_GATE U2983 ( .I1(n2081), .I2(n2083), .O(n2078) );
  NAND_GATE U2984 ( .I1(B[29]), .I2(A[8]), .O(n1977) );
  INV_GATE U2985 ( .I1(n1977), .O(n1971) );
  INV_GATE U2986 ( .I1(n1811), .O(n1808) );
  NAND_GATE U2987 ( .I1(A[7]), .I2(n1848), .O(n1807) );
  NAND_GATE U2988 ( .I1(n1451), .I2(B[31]), .O(n1802) );
  NAND3_GATE U2989 ( .I1(n1450), .I2(n1400), .I3(n1802), .O(n1805) );
  NAND_GATE U2990 ( .I1(A[6]), .I2(n1803), .O(n1804) );
  NAND_GATE U2991 ( .I1(n1805), .I2(n1804), .O(n1806) );
  NAND_GATE U2992 ( .I1(n1807), .I2(n1806), .O(n1809) );
  NAND_GATE U2993 ( .I1(n1808), .I2(n1809), .O(n1813) );
  INV_GATE U2994 ( .I1(n1809), .O(n1810) );
  NAND_GATE U2995 ( .I1(n1811), .I2(n1810), .O(n1812) );
  NAND_GATE U2996 ( .I1(n1813), .I2(n1812), .O(n1970) );
  INV_GATE U2997 ( .I1(n1970), .O(n1973) );
  NAND_GATE U2998 ( .I1(n1971), .I2(n1973), .O(n1968) );
  NAND_GATE U2999 ( .I1(B[29]), .I2(A[7]), .O(n2069) );
  INV_GATE U3000 ( .I1(n2069), .O(n2062) );
  NAND_GATE U3001 ( .I1(n1826), .I2(n1837), .O(n1814) );
  NAND_GATE U3002 ( .I1(A[6]), .I2(n1814), .O(n1818) );
  NAND_GATE U3003 ( .I1(n1450), .I2(B[31]), .O(n1815) );
  NAND_GATE U3004 ( .I1(n1400), .I2(n1815), .O(n1816) );
  NAND_GATE U3005 ( .I1(n1449), .I2(n1816), .O(n1817) );
  NAND_GATE U3006 ( .I1(n1818), .I2(n1817), .O(n1820) );
  NAND_GATE U3007 ( .I1(n1819), .I2(n1820), .O(n1824) );
  INV_GATE U3008 ( .I1(n1820), .O(n1821) );
  NAND_GATE U3009 ( .I1(n1822), .I2(n1821), .O(n1823) );
  NAND_GATE U3010 ( .I1(n1824), .I2(n1823), .O(n2064) );
  NAND_GATE U3011 ( .I1(n2062), .I2(n2064), .O(n2059) );
  NAND_GATE U3012 ( .I1(B[29]), .I2(A[6]), .O(n2052) );
  INV_GATE U3013 ( .I1(n2052), .O(n2047) );
  INV_GATE U3014 ( .I1(n1834), .O(n1831) );
  NAND_GATE U3015 ( .I1(A[5]), .I2(n1848), .O(n1830) );
  NAND_GATE U3016 ( .I1(n1449), .I2(B[31]), .O(n1825) );
  NAND3_GATE U3017 ( .I1(n1448), .I2(n1400), .I3(n1825), .O(n1828) );
  NAND_GATE U3018 ( .I1(A[4]), .I2(n1826), .O(n1827) );
  NAND_GATE U3019 ( .I1(n1828), .I2(n1827), .O(n1829) );
  NAND_GATE U3020 ( .I1(n1830), .I2(n1829), .O(n1832) );
  NAND_GATE U3021 ( .I1(n1831), .I2(n1832), .O(n1836) );
  INV_GATE U3022 ( .I1(n1832), .O(n1833) );
  NAND_GATE U3023 ( .I1(n1834), .I2(n1833), .O(n1835) );
  NAND_GATE U3024 ( .I1(n1836), .I2(n1835), .O(n2048) );
  NAND_GATE U3025 ( .I1(n2047), .I2(n320), .O(n2044) );
  NAND_GATE U3026 ( .I1(B[29]), .I2(A[5]), .O(n1986) );
  INV_GATE U3027 ( .I1(n1986), .O(n1983) );
  NAND_GATE U3028 ( .I1(n1850), .I2(n1837), .O(n1838) );
  NAND_GATE U3029 ( .I1(A[4]), .I2(n1838), .O(n1842) );
  NAND_GATE U3030 ( .I1(n1448), .I2(B[31]), .O(n1839) );
  NAND_GATE U3031 ( .I1(n1400), .I2(n1839), .O(n1840) );
  NAND_GATE U3032 ( .I1(n1447), .I2(n1840), .O(n1841) );
  NAND_GATE U3033 ( .I1(n1842), .I2(n1841), .O(n1843) );
  NAND_GATE U3034 ( .I1(n301), .I2(n1843), .O(n1847) );
  INV_GATE U3035 ( .I1(n1843), .O(n1844) );
  NAND_GATE U3036 ( .I1(n1845), .I2(n1844), .O(n1846) );
  NAND_GATE U3037 ( .I1(n1983), .I2(n1984), .O(n1990) );
  NAND_GATE U3038 ( .I1(B[29]), .I2(A[4]), .O(n2003) );
  INV_GATE U3039 ( .I1(n2003), .O(n2000) );
  NAND_GATE U3040 ( .I1(A[3]), .I2(n1848), .O(n1854) );
  NAND_GATE U3041 ( .I1(n1447), .I2(B[31]), .O(n1849) );
  NAND3_GATE U3042 ( .I1(n1446), .I2(n1400), .I3(n1849), .O(n1852) );
  NAND_GATE U3043 ( .I1(A[2]), .I2(n1850), .O(n1851) );
  NAND_GATE U3044 ( .I1(n1852), .I2(n1851), .O(n1853) );
  NAND_GATE U3045 ( .I1(n1854), .I2(n1853), .O(n1855) );
  NAND_GATE U3046 ( .I1(n1373), .I2(n1855), .O(n1858) );
  NAND_GATE U3047 ( .I1(n2000), .I2(n828), .O(n1996) );
  NAND3_GATE U3048 ( .I1(B[31]), .I2(n1445), .I3(n1442), .O(n1860) );
  NAND3_GATE U3049 ( .I1(B[31]), .I2(n1445), .I3(n1446), .O(n1859) );
  AND_GATE U3050 ( .I1(n1860), .I2(n1859), .O(n1867) );
  NAND_GATE U3051 ( .I1(n1929), .I2(n932), .O(n1862) );
  NAND_GATE U3052 ( .I1(A[2]), .I2(B[30]), .O(n1861) );
  NAND_GATE U3053 ( .I1(n1862), .I2(n1861), .O(n1865) );
  NAND_GATE U3054 ( .I1(B[31]), .I2(n1445), .O(n1864) );
  NAND3_GATE U3055 ( .I1(n1865), .I2(n1864), .I3(n1863), .O(n1866) );
  NAND_GATE U3056 ( .I1(n1867), .I2(n1866), .O(n2013) );
  NAND3_GATE U3057 ( .I1(B[29]), .I2(B[30]), .I3(n1254), .O(n2027) );
  NAND_GATE U3058 ( .I1(B[29]), .I2(A[2]), .O(n2028) );
  NAND3_GATE U3059 ( .I1(A[1]), .I2(n1443), .I3(B[30]), .O(n1869) );
  NAND3_GATE U3060 ( .I1(B[30]), .I2(A[1]), .I3(A[0]), .O(n1868) );
  NAND_GATE U3061 ( .I1(n1869), .I2(n1868), .O(n2030) );
  NAND3_GATE U3062 ( .I1(n2027), .I2(n2032), .I3(n2700), .O(n2011) );
  NAND_GATE U3063 ( .I1(n2013), .I2(n2011), .O(n1872) );
  NAND_GATE U3064 ( .I1(B[29]), .I2(A[3]), .O(n2014) );
  INV_GATE U3065 ( .I1(n2014), .O(n2008) );
  NAND_GATE U3066 ( .I1(n2008), .I2(n2011), .O(n1871) );
  NAND_GATE U3067 ( .I1(n2008), .I2(n2013), .O(n1870) );
  NAND3_GATE U3068 ( .I1(n1872), .I2(n1871), .I3(n1870), .O(n2002) );
  NAND_GATE U3069 ( .I1(n2003), .I2(n940), .O(n1873) );
  NAND_GATE U3070 ( .I1(n2002), .I2(n1873), .O(n1874) );
  NAND_GATE U3071 ( .I1(n1996), .I2(n1874), .O(n1991) );
  NAND_GATE U3072 ( .I1(n1986), .I2(n340), .O(n1875) );
  NAND_GATE U3073 ( .I1(n1991), .I2(n1875), .O(n1876) );
  NAND_GATE U3074 ( .I1(n1990), .I2(n1876), .O(n2049) );
  NAND_GATE U3075 ( .I1(n2052), .I2(n2048), .O(n1877) );
  NAND_GATE U3076 ( .I1(n2049), .I2(n1877), .O(n1878) );
  NAND_GATE U3077 ( .I1(n2044), .I2(n1878), .O(n2065) );
  NAND_GATE U3078 ( .I1(n2069), .I2(n2066), .O(n1879) );
  NAND_GATE U3079 ( .I1(n2065), .I2(n1879), .O(n1880) );
  NAND_GATE U3080 ( .I1(n2059), .I2(n1880), .O(n1972) );
  NAND_GATE U3081 ( .I1(n1977), .I2(n1970), .O(n1881) );
  NAND_GATE U3082 ( .I1(n1972), .I2(n1881), .O(n1882) );
  NAND_GATE U3083 ( .I1(n1968), .I2(n1882), .O(n2084) );
  INV_GATE U3084 ( .I1(n2083), .O(n2085) );
  NAND_GATE U3085 ( .I1(n2088), .I2(n2085), .O(n1883) );
  NAND_GATE U3086 ( .I1(n2084), .I2(n1883), .O(n1884) );
  NAND_GATE U3087 ( .I1(n2078), .I2(n1884), .O(n2099) );
  NAND_GATE U3088 ( .I1(n2104), .I2(n2097), .O(n1885) );
  NAND_GATE U3089 ( .I1(n2099), .I2(n1885), .O(n1886) );
  NAND_GATE U3090 ( .I1(n2095), .I2(n1886), .O(n2117) );
  INV_GATE U3091 ( .I1(n2116), .O(n2118) );
  NAND_GATE U3092 ( .I1(n2121), .I2(n2118), .O(n1887) );
  NAND_GATE U3093 ( .I1(n2117), .I2(n1887), .O(n1888) );
  NAND_GATE U3094 ( .I1(n2111), .I2(n1888), .O(n2132) );
  NAND_GATE U3095 ( .I1(n2137), .I2(n2130), .O(n1889) );
  NAND_GATE U3096 ( .I1(n2132), .I2(n1889), .O(n1890) );
  NAND_GATE U3097 ( .I1(n2128), .I2(n1890), .O(n2150) );
  INV_GATE U3098 ( .I1(n2149), .O(n2151) );
  NAND_GATE U3099 ( .I1(n2154), .I2(n2151), .O(n1891) );
  NAND_GATE U3100 ( .I1(n2150), .I2(n1891), .O(n1892) );
  NAND_GATE U3101 ( .I1(n2144), .I2(n1892), .O(n2165) );
  NAND_GATE U3102 ( .I1(n2170), .I2(n2163), .O(n1893) );
  NAND_GATE U3103 ( .I1(n2165), .I2(n1893), .O(n1894) );
  NAND_GATE U3104 ( .I1(n2161), .I2(n1894), .O(n2183) );
  INV_GATE U3105 ( .I1(n2182), .O(n2184) );
  NAND_GATE U3106 ( .I1(n2187), .I2(n2184), .O(n1895) );
  NAND_GATE U3107 ( .I1(n2183), .I2(n1895), .O(n1896) );
  NAND_GATE U3108 ( .I1(n2177), .I2(n1896), .O(n2198) );
  NAND_GATE U3109 ( .I1(n2203), .I2(n2196), .O(n1897) );
  NAND_GATE U3110 ( .I1(n2198), .I2(n1897), .O(n1898) );
  NAND_GATE U3111 ( .I1(n2194), .I2(n1898), .O(n2216) );
  INV_GATE U3112 ( .I1(n2215), .O(n2217) );
  NAND_GATE U3113 ( .I1(n2220), .I2(n2217), .O(n1899) );
  NAND_GATE U3114 ( .I1(n2216), .I2(n1899), .O(n1900) );
  NAND_GATE U3115 ( .I1(n2210), .I2(n1900), .O(n2231) );
  NAND_GATE U3116 ( .I1(n2236), .I2(n2229), .O(n1901) );
  NAND_GATE U3117 ( .I1(n2231), .I2(n1901), .O(n1902) );
  NAND_GATE U3118 ( .I1(n2227), .I2(n1902), .O(n2249) );
  INV_GATE U3119 ( .I1(n2248), .O(n2250) );
  NAND_GATE U3120 ( .I1(n2253), .I2(n2250), .O(n1903) );
  NAND_GATE U3121 ( .I1(n2249), .I2(n1903), .O(n1904) );
  NAND_GATE U3122 ( .I1(n2243), .I2(n1904), .O(n2264) );
  NAND_GATE U3123 ( .I1(n2269), .I2(n2262), .O(n1905) );
  NAND_GATE U3124 ( .I1(n2264), .I2(n1905), .O(n1906) );
  NAND_GATE U3125 ( .I1(n2260), .I2(n1906), .O(n2282) );
  INV_GATE U3126 ( .I1(n2281), .O(n2283) );
  NAND_GATE U3127 ( .I1(n2286), .I2(n2283), .O(n1907) );
  NAND_GATE U3128 ( .I1(n2282), .I2(n1907), .O(n1908) );
  NAND_GATE U3129 ( .I1(n2276), .I2(n1908), .O(n2297) );
  NAND_GATE U3130 ( .I1(n2302), .I2(n2295), .O(n1909) );
  NAND_GATE U3131 ( .I1(n2297), .I2(n1909), .O(n1910) );
  NAND_GATE U3132 ( .I1(n2293), .I2(n1910), .O(n2315) );
  INV_GATE U3133 ( .I1(n2314), .O(n2316) );
  NAND_GATE U3134 ( .I1(n2319), .I2(n2316), .O(n1911) );
  NAND_GATE U3135 ( .I1(n2315), .I2(n1911), .O(n1912) );
  NAND_GATE U3136 ( .I1(n2309), .I2(n1912), .O(n2330) );
  NAND_GATE U3137 ( .I1(n2335), .I2(n2328), .O(n1913) );
  NAND_GATE U3138 ( .I1(n2330), .I2(n1913), .O(n1914) );
  NAND_GATE U3139 ( .I1(n2326), .I2(n1914), .O(n2348) );
  INV_GATE U3140 ( .I1(n2347), .O(n2349) );
  NAND_GATE U3141 ( .I1(n2352), .I2(n2349), .O(n1915) );
  NAND_GATE U3142 ( .I1(n2348), .I2(n1915), .O(n1916) );
  NAND_GATE U3143 ( .I1(n2342), .I2(n1916), .O(n2363) );
  NAND_GATE U3144 ( .I1(n2368), .I2(n2361), .O(n1917) );
  NAND_GATE U3145 ( .I1(n2363), .I2(n1917), .O(n1918) );
  NAND_GATE U3146 ( .I1(n2359), .I2(n1918), .O(n2381) );
  INV_GATE U3147 ( .I1(n2380), .O(n2382) );
  NAND_GATE U3148 ( .I1(n2385), .I2(n2382), .O(n1919) );
  NAND_GATE U3149 ( .I1(n2381), .I2(n1919), .O(n1920) );
  NAND_GATE U3150 ( .I1(n2375), .I2(n1920), .O(n2396) );
  NAND_GATE U3151 ( .I1(n2401), .I2(n2394), .O(n1921) );
  NAND_GATE U3152 ( .I1(n2396), .I2(n1921), .O(n1922) );
  NAND_GATE U3153 ( .I1(n2392), .I2(n1922), .O(n1959) );
  INV_GATE U3154 ( .I1(n1958), .O(n1960) );
  NAND_GATE U3155 ( .I1(n1963), .I2(n1960), .O(n1923) );
  NAND_GATE U3156 ( .I1(n1959), .I2(n1923), .O(n1924) );
  NAND_GATE U3157 ( .I1(n1953), .I2(n1924), .O(n1943) );
  NAND_GATE U3158 ( .I1(n1948), .I2(n1941), .O(n1925) );
  NAND_GATE U3159 ( .I1(n1943), .I2(n1925), .O(n1927) );
  NAND_GATE U3160 ( .I1(n1441), .I2(A[31]), .O(n1926) );
  NAND3_GATE U3161 ( .I1(n1939), .I2(n1927), .I3(n1926), .O(n2413) );
  NAND_GATE U3162 ( .I1(n2412), .I2(n2413), .O(n1937) );
  NAND_GATE U3163 ( .I1(A[29]), .I2(A[30]), .O(n1928) );
  NAND_GATE U3164 ( .I1(n1929), .I2(n1928), .O(n1935) );
  NAND_GATE U3165 ( .I1(n1475), .I2(n1930), .O(n1933) );
  NAND_GATE U3166 ( .I1(n1442), .I2(n1930), .O(n1931) );
  NAND_GATE U3167 ( .I1(A[31]), .I2(n1931), .O(n1932) );
  NAND_GATE U3168 ( .I1(n1933), .I2(n1932), .O(n1934) );
  NAND_GATE U3169 ( .I1(n1937), .I2(n410), .O(n1938) );
  AND_GATE U3170 ( .I1(n14782), .I2(n1938), .O(\A1[59] ) );
  INV_GATE U3171 ( .I1(n1939), .O(n1940) );
  NAND_GATE U3172 ( .I1(n1940), .I2(n1943), .O(n1952) );
  NAND_GATE U3173 ( .I1(n1942), .I2(n1946), .O(n1950) );
  NAND_GATE U3174 ( .I1(n1944), .I2(n1943), .O(n1945) );
  NAND_GATE U3175 ( .I1(n1946), .I2(n1945), .O(n1947) );
  NAND_GATE U3176 ( .I1(n1948), .I2(n1947), .O(n1949) );
  NAND_GATE U3177 ( .I1(n1950), .I2(n1949), .O(n1951) );
  NAND_GATE U3178 ( .I1(n1952), .I2(n1951), .O(n2418) );
  NAND_GATE U3179 ( .I1(B[28]), .I2(A[30]), .O(n2430) );
  INV_GATE U3180 ( .I1(n2430), .O(n2408) );
  INV_GATE U3181 ( .I1(n1953), .O(n1954) );
  NAND_GATE U3182 ( .I1(n1954), .I2(n1959), .O(n1967) );
  INV_GATE U3183 ( .I1(n1959), .O(n1957) );
  NAND_GATE U3184 ( .I1(n1960), .I2(n1957), .O(n1955) );
  NAND_GATE U3185 ( .I1(n1956), .I2(n1955), .O(n1965) );
  NAND_GATE U3186 ( .I1(n1958), .I2(n1957), .O(n1962) );
  NAND_GATE U3187 ( .I1(n1960), .I2(n1959), .O(n1961) );
  NAND3_GATE U3188 ( .I1(n1963), .I2(n1962), .I3(n1961), .O(n1964) );
  NAND_GATE U3189 ( .I1(n1965), .I2(n1964), .O(n1966) );
  NAND_GATE U3190 ( .I1(n1967), .I2(n1966), .O(n2428) );
  NAND_GATE U3191 ( .I1(n2408), .I2(n2428), .O(n2424) );
  NAND_GATE U3192 ( .I1(B[28]), .I2(A[29]), .O(n2441) );
  INV_GATE U3193 ( .I1(n2441), .O(n2406) );
  NAND_GATE U3194 ( .I1(B[28]), .I2(A[28]), .O(n2452) );
  INV_GATE U3195 ( .I1(n2452), .O(n2390) );
  NAND_GATE U3196 ( .I1(B[28]), .I2(A[27]), .O(n2794) );
  INV_GATE U3197 ( .I1(n2794), .O(n2373) );
  NAND_GATE U3198 ( .I1(B[28]), .I2(A[26]), .O(n2463) );
  INV_GATE U3199 ( .I1(n2463), .O(n2357) );
  NAND_GATE U3200 ( .I1(B[28]), .I2(A[25]), .O(n2474) );
  INV_GATE U3201 ( .I1(n2474), .O(n2340) );
  NAND_GATE U3202 ( .I1(B[28]), .I2(A[24]), .O(n2485) );
  INV_GATE U3203 ( .I1(n2485), .O(n2324) );
  NAND_GATE U3204 ( .I1(B[28]), .I2(A[23]), .O(n2496) );
  INV_GATE U3205 ( .I1(n2496), .O(n2307) );
  NAND_GATE U3206 ( .I1(B[28]), .I2(A[22]), .O(n2507) );
  INV_GATE U3207 ( .I1(n2507), .O(n2291) );
  NAND_GATE U3208 ( .I1(B[28]), .I2(A[21]), .O(n2518) );
  INV_GATE U3209 ( .I1(n2518), .O(n2274) );
  NAND_GATE U3210 ( .I1(B[28]), .I2(A[20]), .O(n2529) );
  INV_GATE U3211 ( .I1(n2529), .O(n2258) );
  NAND_GATE U3212 ( .I1(B[28]), .I2(A[19]), .O(n2540) );
  INV_GATE U3213 ( .I1(n2540), .O(n2241) );
  NAND_GATE U3214 ( .I1(B[28]), .I2(A[18]), .O(n2551) );
  INV_GATE U3215 ( .I1(n2551), .O(n2225) );
  NAND_GATE U3216 ( .I1(B[28]), .I2(A[17]), .O(n2561) );
  INV_GATE U3217 ( .I1(n2561), .O(n2208) );
  NAND_GATE U3218 ( .I1(B[28]), .I2(A[16]), .O(n2572) );
  INV_GATE U3219 ( .I1(n2572), .O(n2192) );
  NAND_GATE U3220 ( .I1(B[28]), .I2(A[15]), .O(n2583) );
  INV_GATE U3221 ( .I1(n2583), .O(n2175) );
  NAND_GATE U3222 ( .I1(B[28]), .I2(A[14]), .O(n2594) );
  INV_GATE U3223 ( .I1(n2594), .O(n2159) );
  NAND_GATE U3224 ( .I1(B[28]), .I2(A[13]), .O(n2605) );
  INV_GATE U3225 ( .I1(n2605), .O(n2142) );
  NAND_GATE U3226 ( .I1(B[28]), .I2(A[12]), .O(n2616) );
  INV_GATE U3227 ( .I1(n2616), .O(n2126) );
  NAND_GATE U3228 ( .I1(B[28]), .I2(A[11]), .O(n2627) );
  INV_GATE U3229 ( .I1(n2627), .O(n2109) );
  NAND_GATE U3230 ( .I1(B[28]), .I2(A[10]), .O(n2638) );
  INV_GATE U3231 ( .I1(n2638), .O(n2093) );
  NAND_GATE U3232 ( .I1(B[28]), .I2(A[9]), .O(n2642) );
  INV_GATE U3233 ( .I1(n2642), .O(n2076) );
  INV_GATE U3234 ( .I1(n1968), .O(n1969) );
  NAND_GATE U3235 ( .I1(n1969), .I2(n1972), .O(n1981) );
  NAND_GATE U3236 ( .I1(n1971), .I2(n1975), .O(n1979) );
  NAND_GATE U3237 ( .I1(n1973), .I2(n1972), .O(n1974) );
  NAND_GATE U3238 ( .I1(n1975), .I2(n1974), .O(n1976) );
  NAND_GATE U3239 ( .I1(n1977), .I2(n1976), .O(n1978) );
  NAND_GATE U3240 ( .I1(n1979), .I2(n1978), .O(n1980) );
  NAND_GATE U3241 ( .I1(n1981), .I2(n1980), .O(n2645) );
  NAND_GATE U3242 ( .I1(n2076), .I2(n2645), .O(n2647) );
  NAND_GATE U3243 ( .I1(B[28]), .I2(A[8]), .O(n2658) );
  INV_GATE U3244 ( .I1(n2658), .O(n2653) );
  NAND_GATE U3245 ( .I1(B[28]), .I2(A[7]), .O(n2667) );
  INV_GATE U3246 ( .I1(n2667), .O(n2669) );
  NAND_GATE U3247 ( .I1(n340), .I2(n813), .O(n1982) );
  NAND_GATE U3248 ( .I1(n1983), .I2(n1982), .O(n1988) );
  NAND_GATE U3249 ( .I1(n1984), .I2(n813), .O(n1985) );
  NAND_GATE U3250 ( .I1(n1986), .I2(n1985), .O(n1987) );
  NAND_GATE U3251 ( .I1(n1988), .I2(n1987), .O(n1995) );
  AND_GATE U3252 ( .I1(n340), .I2(n1991), .O(n1989) );
  NAND_GATE U3253 ( .I1(n1989), .I2(n1988), .O(n1994) );
  INV_GATE U3254 ( .I1(n1990), .O(n1992) );
  NAND_GATE U3255 ( .I1(n1992), .I2(n1991), .O(n1993) );
  NAND3_GATE U3256 ( .I1(n1995), .I2(n1994), .I3(n1993), .O(n2674) );
  INV_GATE U3257 ( .I1(n2002), .O(n2001) );
  NAND_GATE U3258 ( .I1(n940), .I2(n2001), .O(n1999) );
  INV_GATE U3259 ( .I1(n1996), .O(n1997) );
  NAND_GATE U3260 ( .I1(n1997), .I2(n2002), .O(n1998) );
  NAND3_GATE U3261 ( .I1(n2000), .I2(n1999), .I3(n1998), .O(n2007) );
  NAND_GATE U3262 ( .I1(n828), .I2(n2001), .O(n2005) );
  NAND_GATE U3263 ( .I1(n940), .I2(n2002), .O(n2004) );
  NAND3_GATE U3264 ( .I1(n2005), .I2(n2004), .I3(n2003), .O(n2006) );
  NAND_GATE U3265 ( .I1(n2007), .I2(n2006), .O(n2688) );
  NAND3_GATE U3266 ( .I1(n2011), .I2(n349), .I3(n2008), .O(n2010) );
  INV_GATE U3267 ( .I1(n2011), .O(n2012) );
  NAND3_GATE U3268 ( .I1(n2013), .I2(n2012), .I3(n2008), .O(n2009) );
  AND_GATE U3269 ( .I1(n2010), .I2(n2009), .O(n2018) );
  NAND_GATE U3270 ( .I1(n349), .I2(n2011), .O(n2016) );
  NAND_GATE U3271 ( .I1(n2013), .I2(n2012), .O(n2015) );
  NAND3_GATE U3272 ( .I1(n2016), .I2(n2015), .I3(n2014), .O(n2017) );
  NAND_GATE U3273 ( .I1(n2018), .I2(n2017), .O(n2735) );
  NAND_GATE U3274 ( .I1(B[28]), .I2(A[4]), .O(n2736) );
  INV_GATE U3275 ( .I1(n2736), .O(n2738) );
  NAND_GATE U3276 ( .I1(B[28]), .I2(A[3]), .O(n2708) );
  INV_GATE U3277 ( .I1(n2708), .O(n2701) );
  NAND_GATE U3278 ( .I1(B[28]), .I2(A[2]), .O(n2720) );
  INV_GATE U3279 ( .I1(n2720), .O(n2724) );
  NAND_GATE U3280 ( .I1(n1441), .I2(A[0]), .O(n2019) );
  NAND_GATE U3281 ( .I1(n14241), .I2(n2019), .O(n2020) );
  NAND_GATE U3282 ( .I1(B[30]), .I2(n2020), .O(n2716) );
  NAND_GATE U3283 ( .I1(B[29]), .I2(n2021), .O(n2717) );
  NAND_GATE U3284 ( .I1(n2724), .I2(n1281), .O(n2024) );
  NAND3_GATE U3285 ( .I1(B[28]), .I2(B[29]), .I3(n1254), .O(n2719) );
  INV_GATE U3286 ( .I1(n2719), .O(n2723) );
  NAND_GATE U3287 ( .I1(n2716), .I2(n919), .O(n2022) );
  NAND_GATE U3288 ( .I1(n2723), .I2(n2022), .O(n2023) );
  NAND_GATE U3289 ( .I1(n2024), .I2(n2023), .O(n2704) );
  NAND_GATE U3290 ( .I1(n2701), .I2(n2704), .O(n2697) );
  INV_GATE U3291 ( .I1(n2030), .O(n2026) );
  NAND3_GATE U3292 ( .I1(n2026), .I2(n2025), .I3(n2028), .O(n2699) );
  INV_GATE U3293 ( .I1(n2027), .O(n2029) );
  NAND_GATE U3294 ( .I1(n2029), .I2(n2028), .O(n2698) );
  NAND_GATE U3295 ( .I1(n2699), .I2(n2698), .O(n2693) );
  INV_GATE U3296 ( .I1(n2693), .O(n2033) );
  NAND_GATE U3297 ( .I1(n2029), .I2(n2031), .O(n2696) );
  NAND_GATE U3298 ( .I1(n2031), .I2(n2030), .O(n2032) );
  NAND_GATE U3299 ( .I1(n2032), .I2(n2700), .O(n2694) );
  NAND_GATE U3300 ( .I1(n2696), .I2(n2694), .O(n2034) );
  NAND3_GATE U3301 ( .I1(n2033), .I2(n2701), .I3(n2034), .O(n2036) );
  NAND3_GATE U3302 ( .I1(n2034), .I2(n2033), .I3(n2704), .O(n2035) );
  NAND3_GATE U3303 ( .I1(n2697), .I2(n2036), .I3(n2035), .O(n2737) );
  NAND_GATE U3304 ( .I1(n2735), .I2(n2736), .O(n2037) );
  NAND_GATE U3305 ( .I1(n2737), .I2(n2037), .O(n2038) );
  NAND_GATE U3306 ( .I1(n2740), .I2(n2038), .O(n2687) );
  NAND_GATE U3307 ( .I1(n2689), .I2(n2687), .O(n2041) );
  NAND_GATE U3308 ( .I1(B[28]), .I2(A[5]), .O(n2690) );
  INV_GATE U3309 ( .I1(n2690), .O(n2684) );
  NAND_GATE U3310 ( .I1(n2684), .I2(n2687), .O(n2040) );
  NAND_GATE U3311 ( .I1(n2684), .I2(n2689), .O(n2039) );
  NAND3_GATE U3312 ( .I1(n2041), .I2(n2040), .I3(n2039), .O(n2680) );
  NAND_GATE U3313 ( .I1(n2674), .I2(n2680), .O(n2043) );
  NAND_GATE U3314 ( .I1(B[28]), .I2(A[6]), .O(n2677) );
  INV_GATE U3315 ( .I1(n2677), .O(n2679) );
  NAND_GATE U3316 ( .I1(n2679), .I2(n2680), .O(n2042) );
  NAND_GATE U3317 ( .I1(n2679), .I2(n2674), .O(n2678) );
  NAND3_GATE U3318 ( .I1(n2043), .I2(n2042), .I3(n2678), .O(n2670) );
  NAND_GATE U3319 ( .I1(n2669), .I2(n2670), .O(n2058) );
  INV_GATE U3320 ( .I1(n2044), .O(n2045) );
  NAND_GATE U3321 ( .I1(n2045), .I2(n2049), .O(n2056) );
  NAND_GATE U3322 ( .I1(n2048), .I2(n839), .O(n2046) );
  NAND_GATE U3323 ( .I1(n2047), .I2(n2046), .O(n2054) );
  NAND_GATE U3324 ( .I1(n320), .I2(n2049), .O(n2050) );
  NAND_GATE U3325 ( .I1(n2046), .I2(n2050), .O(n2051) );
  NAND_GATE U3326 ( .I1(n2052), .I2(n2051), .O(n2053) );
  NAND_GATE U3327 ( .I1(n2054), .I2(n2053), .O(n2055) );
  NAND_GATE U3328 ( .I1(n2056), .I2(n2055), .O(n2663) );
  NAND_GATE U3329 ( .I1(n2670), .I2(n2663), .O(n2057) );
  NAND_GATE U3330 ( .I1(n2669), .I2(n2663), .O(n2668) );
  NAND3_GATE U3331 ( .I1(n2058), .I2(n2057), .I3(n2668), .O(n2657) );
  NAND_GATE U3332 ( .I1(n2653), .I2(n2657), .O(n2075) );
  INV_GATE U3333 ( .I1(n2059), .O(n2060) );
  NAND_GATE U3334 ( .I1(n2060), .I2(n2065), .O(n2073) );
  INV_GATE U3335 ( .I1(n2065), .O(n2063) );
  NAND_GATE U3336 ( .I1(n2066), .I2(n2063), .O(n2061) );
  NAND_GATE U3337 ( .I1(n2062), .I2(n2061), .O(n2071) );
  NAND_GATE U3338 ( .I1(n2064), .I2(n2063), .O(n2068) );
  NAND_GATE U3339 ( .I1(n2066), .I2(n2065), .O(n2067) );
  NAND3_GATE U3340 ( .I1(n2069), .I2(n2068), .I3(n2067), .O(n2070) );
  NAND_GATE U3341 ( .I1(n2071), .I2(n2070), .O(n2072) );
  NAND_GATE U3342 ( .I1(n2073), .I2(n2072), .O(n2656) );
  NAND_GATE U3343 ( .I1(n2656), .I2(n2657), .O(n2074) );
  NAND_GATE U3344 ( .I1(n2653), .I2(n2656), .O(n2652) );
  NAND3_GATE U3345 ( .I1(n2075), .I2(n2074), .I3(n2652), .O(n2648) );
  NAND_GATE U3346 ( .I1(n2076), .I2(n2648), .O(n2646) );
  NAND_GATE U3347 ( .I1(n2645), .I2(n2648), .O(n2077) );
  NAND3_GATE U3348 ( .I1(n2647), .I2(n2646), .I3(n2077), .O(n2637) );
  NAND_GATE U3349 ( .I1(n2093), .I2(n2637), .O(n2633) );
  INV_GATE U3350 ( .I1(n2078), .O(n2079) );
  NAND_GATE U3351 ( .I1(n2079), .I2(n2084), .O(n2092) );
  INV_GATE U3352 ( .I1(n2084), .O(n2082) );
  NAND_GATE U3353 ( .I1(n2085), .I2(n2082), .O(n2080) );
  NAND_GATE U3354 ( .I1(n2081), .I2(n2080), .O(n2090) );
  NAND_GATE U3355 ( .I1(n2083), .I2(n2082), .O(n2087) );
  NAND_GATE U3356 ( .I1(n2085), .I2(n2084), .O(n2086) );
  NAND3_GATE U3357 ( .I1(n2088), .I2(n2087), .I3(n2086), .O(n2089) );
  NAND_GATE U3358 ( .I1(n2090), .I2(n2089), .O(n2091) );
  NAND_GATE U3359 ( .I1(n2092), .I2(n2091), .O(n2636) );
  NAND_GATE U3360 ( .I1(n2093), .I2(n2636), .O(n2632) );
  NAND_GATE U3361 ( .I1(n2637), .I2(n2636), .O(n2094) );
  NAND3_GATE U3362 ( .I1(n2633), .I2(n2632), .I3(n2094), .O(n2626) );
  NAND_GATE U3363 ( .I1(n2109), .I2(n2626), .O(n2622) );
  INV_GATE U3364 ( .I1(n2095), .O(n2096) );
  NAND_GATE U3365 ( .I1(n2096), .I2(n2099), .O(n2108) );
  NAND_GATE U3366 ( .I1(n2098), .I2(n2102), .O(n2106) );
  NAND_GATE U3367 ( .I1(n2100), .I2(n2099), .O(n2101) );
  NAND_GATE U3368 ( .I1(n2102), .I2(n2101), .O(n2103) );
  NAND_GATE U3369 ( .I1(n2104), .I2(n2103), .O(n2105) );
  NAND_GATE U3370 ( .I1(n2106), .I2(n2105), .O(n2107) );
  NAND_GATE U3371 ( .I1(n2108), .I2(n2107), .O(n2625) );
  NAND_GATE U3372 ( .I1(n2109), .I2(n2625), .O(n2621) );
  NAND_GATE U3373 ( .I1(n2626), .I2(n2625), .O(n2110) );
  NAND3_GATE U3374 ( .I1(n2622), .I2(n2621), .I3(n2110), .O(n2615) );
  NAND_GATE U3375 ( .I1(n2126), .I2(n2615), .O(n2611) );
  INV_GATE U3376 ( .I1(n2111), .O(n2112) );
  NAND_GATE U3377 ( .I1(n2112), .I2(n2117), .O(n2125) );
  INV_GATE U3378 ( .I1(n2117), .O(n2115) );
  NAND_GATE U3379 ( .I1(n2118), .I2(n2115), .O(n2113) );
  NAND_GATE U3380 ( .I1(n2114), .I2(n2113), .O(n2123) );
  NAND_GATE U3381 ( .I1(n2116), .I2(n2115), .O(n2120) );
  NAND_GATE U3382 ( .I1(n2118), .I2(n2117), .O(n2119) );
  NAND3_GATE U3383 ( .I1(n2121), .I2(n2120), .I3(n2119), .O(n2122) );
  NAND_GATE U3384 ( .I1(n2123), .I2(n2122), .O(n2124) );
  NAND_GATE U3385 ( .I1(n2125), .I2(n2124), .O(n2614) );
  NAND_GATE U3386 ( .I1(n2126), .I2(n2614), .O(n2610) );
  NAND_GATE U3387 ( .I1(n2615), .I2(n2614), .O(n2127) );
  NAND3_GATE U3388 ( .I1(n2611), .I2(n2610), .I3(n2127), .O(n2604) );
  NAND_GATE U3389 ( .I1(n2142), .I2(n2604), .O(n2600) );
  INV_GATE U3390 ( .I1(n2128), .O(n2129) );
  NAND_GATE U3391 ( .I1(n2129), .I2(n2132), .O(n2141) );
  NAND_GATE U3392 ( .I1(n2131), .I2(n2135), .O(n2139) );
  NAND_GATE U3393 ( .I1(n2133), .I2(n2132), .O(n2134) );
  NAND_GATE U3394 ( .I1(n2135), .I2(n2134), .O(n2136) );
  NAND_GATE U3395 ( .I1(n2137), .I2(n2136), .O(n2138) );
  NAND_GATE U3396 ( .I1(n2139), .I2(n2138), .O(n2140) );
  NAND_GATE U3397 ( .I1(n2141), .I2(n2140), .O(n2603) );
  NAND_GATE U3398 ( .I1(n2142), .I2(n2603), .O(n2599) );
  NAND_GATE U3399 ( .I1(n2604), .I2(n2603), .O(n2143) );
  NAND3_GATE U3400 ( .I1(n2600), .I2(n2599), .I3(n2143), .O(n2593) );
  NAND_GATE U3401 ( .I1(n2159), .I2(n2593), .O(n2589) );
  INV_GATE U3402 ( .I1(n2144), .O(n2145) );
  NAND_GATE U3403 ( .I1(n2145), .I2(n2150), .O(n2158) );
  INV_GATE U3404 ( .I1(n2150), .O(n2148) );
  NAND_GATE U3405 ( .I1(n2151), .I2(n2148), .O(n2146) );
  NAND_GATE U3406 ( .I1(n2147), .I2(n2146), .O(n2156) );
  NAND_GATE U3407 ( .I1(n2149), .I2(n2148), .O(n2153) );
  NAND_GATE U3408 ( .I1(n2151), .I2(n2150), .O(n2152) );
  NAND3_GATE U3409 ( .I1(n2154), .I2(n2153), .I3(n2152), .O(n2155) );
  NAND_GATE U3410 ( .I1(n2156), .I2(n2155), .O(n2157) );
  NAND_GATE U3411 ( .I1(n2158), .I2(n2157), .O(n2592) );
  NAND_GATE U3412 ( .I1(n2159), .I2(n2592), .O(n2588) );
  NAND_GATE U3413 ( .I1(n2593), .I2(n2592), .O(n2160) );
  NAND3_GATE U3414 ( .I1(n2589), .I2(n2588), .I3(n2160), .O(n2582) );
  NAND_GATE U3415 ( .I1(n2175), .I2(n2582), .O(n2578) );
  INV_GATE U3416 ( .I1(n2161), .O(n2162) );
  NAND_GATE U3417 ( .I1(n2162), .I2(n2165), .O(n2174) );
  NAND_GATE U3418 ( .I1(n2164), .I2(n2168), .O(n2172) );
  NAND_GATE U3419 ( .I1(n2166), .I2(n2165), .O(n2167) );
  NAND_GATE U3420 ( .I1(n2168), .I2(n2167), .O(n2169) );
  NAND_GATE U3421 ( .I1(n2170), .I2(n2169), .O(n2171) );
  NAND_GATE U3422 ( .I1(n2172), .I2(n2171), .O(n2173) );
  NAND_GATE U3423 ( .I1(n2174), .I2(n2173), .O(n2581) );
  NAND_GATE U3424 ( .I1(n2175), .I2(n2581), .O(n2577) );
  NAND_GATE U3425 ( .I1(n2582), .I2(n2581), .O(n2176) );
  NAND3_GATE U3426 ( .I1(n2578), .I2(n2577), .I3(n2176), .O(n2571) );
  NAND_GATE U3427 ( .I1(n2192), .I2(n2571), .O(n2567) );
  INV_GATE U3428 ( .I1(n2177), .O(n2178) );
  NAND_GATE U3429 ( .I1(n2178), .I2(n2183), .O(n2191) );
  INV_GATE U3430 ( .I1(n2183), .O(n2181) );
  NAND_GATE U3431 ( .I1(n2184), .I2(n2181), .O(n2179) );
  NAND_GATE U3432 ( .I1(n2180), .I2(n2179), .O(n2189) );
  NAND_GATE U3433 ( .I1(n2182), .I2(n2181), .O(n2186) );
  NAND_GATE U3434 ( .I1(n2184), .I2(n2183), .O(n2185) );
  NAND3_GATE U3435 ( .I1(n2187), .I2(n2186), .I3(n2185), .O(n2188) );
  NAND_GATE U3436 ( .I1(n2189), .I2(n2188), .O(n2190) );
  NAND_GATE U3437 ( .I1(n2191), .I2(n2190), .O(n2570) );
  NAND_GATE U3438 ( .I1(n2192), .I2(n2570), .O(n2566) );
  NAND_GATE U3439 ( .I1(n2571), .I2(n2570), .O(n2193) );
  NAND3_GATE U3440 ( .I1(n2567), .I2(n2566), .I3(n2193), .O(n2560) );
  NAND_GATE U3441 ( .I1(n2208), .I2(n2560), .O(n2556) );
  INV_GATE U3442 ( .I1(n2194), .O(n2195) );
  NAND_GATE U3443 ( .I1(n2195), .I2(n2198), .O(n2207) );
  NAND_GATE U3444 ( .I1(n2197), .I2(n2201), .O(n2205) );
  NAND_GATE U3445 ( .I1(n2199), .I2(n2198), .O(n2200) );
  NAND_GATE U3446 ( .I1(n2201), .I2(n2200), .O(n2202) );
  NAND_GATE U3447 ( .I1(n2203), .I2(n2202), .O(n2204) );
  NAND_GATE U3448 ( .I1(n2205), .I2(n2204), .O(n2206) );
  NAND_GATE U3449 ( .I1(n2207), .I2(n2206), .O(n2559) );
  NAND_GATE U3450 ( .I1(n2208), .I2(n2559), .O(n2555) );
  NAND_GATE U3451 ( .I1(n2560), .I2(n2559), .O(n2209) );
  NAND3_GATE U3452 ( .I1(n2556), .I2(n2555), .I3(n2209), .O(n2550) );
  NAND_GATE U3453 ( .I1(n2225), .I2(n2550), .O(n2546) );
  INV_GATE U3454 ( .I1(n2210), .O(n2211) );
  NAND_GATE U3455 ( .I1(n2211), .I2(n2216), .O(n2224) );
  INV_GATE U3456 ( .I1(n2216), .O(n2214) );
  NAND_GATE U3457 ( .I1(n2217), .I2(n2214), .O(n2212) );
  NAND_GATE U3458 ( .I1(n2213), .I2(n2212), .O(n2222) );
  NAND_GATE U3459 ( .I1(n2215), .I2(n2214), .O(n2219) );
  NAND_GATE U3460 ( .I1(n2217), .I2(n2216), .O(n2218) );
  NAND3_GATE U3461 ( .I1(n2220), .I2(n2219), .I3(n2218), .O(n2221) );
  NAND_GATE U3462 ( .I1(n2222), .I2(n2221), .O(n2223) );
  NAND_GATE U3463 ( .I1(n2224), .I2(n2223), .O(n2549) );
  NAND_GATE U3464 ( .I1(n2225), .I2(n2549), .O(n2545) );
  NAND_GATE U3465 ( .I1(n2550), .I2(n2549), .O(n2226) );
  NAND3_GATE U3466 ( .I1(n2546), .I2(n2545), .I3(n2226), .O(n2539) );
  NAND_GATE U3467 ( .I1(n2241), .I2(n2539), .O(n2535) );
  INV_GATE U3468 ( .I1(n2227), .O(n2228) );
  NAND_GATE U3469 ( .I1(n2228), .I2(n2231), .O(n2240) );
  NAND_GATE U3470 ( .I1(n2230), .I2(n2234), .O(n2238) );
  NAND_GATE U3471 ( .I1(n2232), .I2(n2231), .O(n2233) );
  NAND_GATE U3472 ( .I1(n2234), .I2(n2233), .O(n2235) );
  NAND_GATE U3473 ( .I1(n2236), .I2(n2235), .O(n2237) );
  NAND_GATE U3474 ( .I1(n2238), .I2(n2237), .O(n2239) );
  NAND_GATE U3475 ( .I1(n2240), .I2(n2239), .O(n2538) );
  NAND_GATE U3476 ( .I1(n2241), .I2(n2538), .O(n2534) );
  NAND_GATE U3477 ( .I1(n2539), .I2(n2538), .O(n2242) );
  NAND3_GATE U3478 ( .I1(n2535), .I2(n2534), .I3(n2242), .O(n2528) );
  NAND_GATE U3479 ( .I1(n2258), .I2(n2528), .O(n2524) );
  INV_GATE U3480 ( .I1(n2243), .O(n2244) );
  NAND_GATE U3481 ( .I1(n2244), .I2(n2249), .O(n2257) );
  INV_GATE U3482 ( .I1(n2249), .O(n2247) );
  NAND_GATE U3483 ( .I1(n2250), .I2(n2247), .O(n2245) );
  NAND_GATE U3484 ( .I1(n2246), .I2(n2245), .O(n2255) );
  NAND_GATE U3485 ( .I1(n2248), .I2(n2247), .O(n2252) );
  NAND_GATE U3486 ( .I1(n2250), .I2(n2249), .O(n2251) );
  NAND3_GATE U3487 ( .I1(n2253), .I2(n2252), .I3(n2251), .O(n2254) );
  NAND_GATE U3488 ( .I1(n2255), .I2(n2254), .O(n2256) );
  NAND_GATE U3489 ( .I1(n2257), .I2(n2256), .O(n2527) );
  NAND_GATE U3490 ( .I1(n2258), .I2(n2527), .O(n2523) );
  NAND_GATE U3491 ( .I1(n2528), .I2(n2527), .O(n2259) );
  NAND3_GATE U3492 ( .I1(n2524), .I2(n2523), .I3(n2259), .O(n2517) );
  NAND_GATE U3493 ( .I1(n2274), .I2(n2517), .O(n2513) );
  INV_GATE U3494 ( .I1(n2260), .O(n2261) );
  NAND_GATE U3495 ( .I1(n2261), .I2(n2264), .O(n2273) );
  NAND_GATE U3496 ( .I1(n2263), .I2(n2267), .O(n2271) );
  NAND_GATE U3497 ( .I1(n2265), .I2(n2264), .O(n2266) );
  NAND_GATE U3498 ( .I1(n2267), .I2(n2266), .O(n2268) );
  NAND_GATE U3499 ( .I1(n2269), .I2(n2268), .O(n2270) );
  NAND_GATE U3500 ( .I1(n2271), .I2(n2270), .O(n2272) );
  NAND_GATE U3501 ( .I1(n2273), .I2(n2272), .O(n2516) );
  NAND_GATE U3502 ( .I1(n2274), .I2(n2516), .O(n2512) );
  NAND_GATE U3503 ( .I1(n2517), .I2(n2516), .O(n2275) );
  NAND3_GATE U3504 ( .I1(n2513), .I2(n2512), .I3(n2275), .O(n2506) );
  NAND_GATE U3505 ( .I1(n2291), .I2(n2506), .O(n2502) );
  INV_GATE U3506 ( .I1(n2276), .O(n2277) );
  NAND_GATE U3507 ( .I1(n2277), .I2(n2282), .O(n2290) );
  INV_GATE U3508 ( .I1(n2282), .O(n2280) );
  NAND_GATE U3509 ( .I1(n2283), .I2(n2280), .O(n2278) );
  NAND_GATE U3510 ( .I1(n2279), .I2(n2278), .O(n2288) );
  NAND_GATE U3511 ( .I1(n2281), .I2(n2280), .O(n2285) );
  NAND_GATE U3512 ( .I1(n2283), .I2(n2282), .O(n2284) );
  NAND3_GATE U3513 ( .I1(n2286), .I2(n2285), .I3(n2284), .O(n2287) );
  NAND_GATE U3514 ( .I1(n2288), .I2(n2287), .O(n2289) );
  NAND_GATE U3515 ( .I1(n2290), .I2(n2289), .O(n2505) );
  NAND_GATE U3516 ( .I1(n2291), .I2(n2505), .O(n2501) );
  NAND_GATE U3517 ( .I1(n2506), .I2(n2505), .O(n2292) );
  NAND3_GATE U3518 ( .I1(n2502), .I2(n2501), .I3(n2292), .O(n2495) );
  NAND_GATE U3519 ( .I1(n2307), .I2(n2495), .O(n2491) );
  INV_GATE U3520 ( .I1(n2293), .O(n2294) );
  NAND_GATE U3521 ( .I1(n2294), .I2(n2297), .O(n2306) );
  NAND_GATE U3522 ( .I1(n2296), .I2(n2300), .O(n2304) );
  NAND_GATE U3523 ( .I1(n2298), .I2(n2297), .O(n2299) );
  NAND_GATE U3524 ( .I1(n2300), .I2(n2299), .O(n2301) );
  NAND_GATE U3525 ( .I1(n2302), .I2(n2301), .O(n2303) );
  NAND_GATE U3526 ( .I1(n2304), .I2(n2303), .O(n2305) );
  NAND_GATE U3527 ( .I1(n2306), .I2(n2305), .O(n2494) );
  NAND_GATE U3528 ( .I1(n2307), .I2(n2494), .O(n2490) );
  NAND_GATE U3529 ( .I1(n2495), .I2(n2494), .O(n2308) );
  NAND3_GATE U3530 ( .I1(n2491), .I2(n2490), .I3(n2308), .O(n2484) );
  NAND_GATE U3531 ( .I1(n2324), .I2(n2484), .O(n2480) );
  INV_GATE U3532 ( .I1(n2309), .O(n2310) );
  NAND_GATE U3533 ( .I1(n2310), .I2(n2315), .O(n2323) );
  INV_GATE U3534 ( .I1(n2315), .O(n2313) );
  NAND_GATE U3535 ( .I1(n2316), .I2(n2313), .O(n2311) );
  NAND_GATE U3536 ( .I1(n2312), .I2(n2311), .O(n2321) );
  NAND_GATE U3537 ( .I1(n2314), .I2(n2313), .O(n2318) );
  NAND_GATE U3538 ( .I1(n2316), .I2(n2315), .O(n2317) );
  NAND3_GATE U3539 ( .I1(n2319), .I2(n2318), .I3(n2317), .O(n2320) );
  NAND_GATE U3540 ( .I1(n2321), .I2(n2320), .O(n2322) );
  NAND_GATE U3541 ( .I1(n2323), .I2(n2322), .O(n2483) );
  NAND_GATE U3542 ( .I1(n2324), .I2(n2483), .O(n2479) );
  NAND_GATE U3543 ( .I1(n2484), .I2(n2483), .O(n2325) );
  NAND3_GATE U3544 ( .I1(n2480), .I2(n2479), .I3(n2325), .O(n2473) );
  NAND_GATE U3545 ( .I1(n2340), .I2(n2473), .O(n2469) );
  INV_GATE U3546 ( .I1(n2326), .O(n2327) );
  NAND_GATE U3547 ( .I1(n2327), .I2(n2330), .O(n2339) );
  NAND_GATE U3548 ( .I1(n2329), .I2(n2333), .O(n2337) );
  NAND_GATE U3549 ( .I1(n2331), .I2(n2330), .O(n2332) );
  NAND_GATE U3550 ( .I1(n2333), .I2(n2332), .O(n2334) );
  NAND_GATE U3551 ( .I1(n2335), .I2(n2334), .O(n2336) );
  NAND_GATE U3552 ( .I1(n2337), .I2(n2336), .O(n2338) );
  NAND_GATE U3553 ( .I1(n2339), .I2(n2338), .O(n2472) );
  NAND_GATE U3554 ( .I1(n2340), .I2(n2472), .O(n2468) );
  NAND_GATE U3555 ( .I1(n2473), .I2(n2472), .O(n2341) );
  NAND3_GATE U3556 ( .I1(n2469), .I2(n2468), .I3(n2341), .O(n2462) );
  NAND_GATE U3557 ( .I1(n2357), .I2(n2462), .O(n2458) );
  INV_GATE U3558 ( .I1(n2342), .O(n2343) );
  NAND_GATE U3559 ( .I1(n2343), .I2(n2348), .O(n2356) );
  INV_GATE U3560 ( .I1(n2348), .O(n2346) );
  NAND_GATE U3561 ( .I1(n2349), .I2(n2346), .O(n2344) );
  NAND_GATE U3562 ( .I1(n2345), .I2(n2344), .O(n2354) );
  NAND_GATE U3563 ( .I1(n2347), .I2(n2346), .O(n2351) );
  NAND_GATE U3564 ( .I1(n2349), .I2(n2348), .O(n2350) );
  NAND3_GATE U3565 ( .I1(n2352), .I2(n2351), .I3(n2350), .O(n2353) );
  NAND_GATE U3566 ( .I1(n2354), .I2(n2353), .O(n2355) );
  NAND_GATE U3567 ( .I1(n2356), .I2(n2355), .O(n2461) );
  NAND_GATE U3568 ( .I1(n2357), .I2(n2461), .O(n2457) );
  NAND_GATE U3569 ( .I1(n2462), .I2(n2461), .O(n2358) );
  NAND3_GATE U3570 ( .I1(n2458), .I2(n2457), .I3(n2358), .O(n2793) );
  NAND_GATE U3571 ( .I1(n2373), .I2(n2793), .O(n2789) );
  INV_GATE U3572 ( .I1(n2359), .O(n2360) );
  NAND_GATE U3573 ( .I1(n2360), .I2(n2363), .O(n2372) );
  NAND_GATE U3574 ( .I1(n2362), .I2(n2366), .O(n2370) );
  NAND_GATE U3575 ( .I1(n2364), .I2(n2363), .O(n2365) );
  NAND_GATE U3576 ( .I1(n2366), .I2(n2365), .O(n2367) );
  NAND_GATE U3577 ( .I1(n2368), .I2(n2367), .O(n2369) );
  NAND_GATE U3578 ( .I1(n2370), .I2(n2369), .O(n2371) );
  NAND_GATE U3579 ( .I1(n2372), .I2(n2371), .O(n2792) );
  NAND_GATE U3580 ( .I1(n2373), .I2(n2792), .O(n2788) );
  NAND_GATE U3581 ( .I1(n2793), .I2(n2792), .O(n2374) );
  NAND3_GATE U3582 ( .I1(n2789), .I2(n2788), .I3(n2374), .O(n2451) );
  NAND_GATE U3583 ( .I1(n2390), .I2(n2451), .O(n2447) );
  INV_GATE U3584 ( .I1(n2375), .O(n2376) );
  NAND_GATE U3585 ( .I1(n2376), .I2(n2381), .O(n2389) );
  INV_GATE U3586 ( .I1(n2381), .O(n2379) );
  NAND_GATE U3587 ( .I1(n2382), .I2(n2379), .O(n2377) );
  NAND_GATE U3588 ( .I1(n2378), .I2(n2377), .O(n2387) );
  NAND_GATE U3589 ( .I1(n2380), .I2(n2379), .O(n2384) );
  NAND_GATE U3590 ( .I1(n2382), .I2(n2381), .O(n2383) );
  NAND3_GATE U3591 ( .I1(n2385), .I2(n2384), .I3(n2383), .O(n2386) );
  NAND_GATE U3592 ( .I1(n2387), .I2(n2386), .O(n2388) );
  NAND_GATE U3593 ( .I1(n2389), .I2(n2388), .O(n2450) );
  NAND_GATE U3594 ( .I1(n2390), .I2(n2450), .O(n2446) );
  NAND_GATE U3595 ( .I1(n2451), .I2(n2450), .O(n2391) );
  NAND3_GATE U3596 ( .I1(n2447), .I2(n2446), .I3(n2391), .O(n2440) );
  NAND_GATE U3597 ( .I1(n2406), .I2(n2440), .O(n2436) );
  INV_GATE U3598 ( .I1(n2392), .O(n2393) );
  NAND_GATE U3599 ( .I1(n2393), .I2(n2396), .O(n2405) );
  NAND_GATE U3600 ( .I1(n2395), .I2(n2399), .O(n2403) );
  NAND_GATE U3601 ( .I1(n2397), .I2(n2396), .O(n2398) );
  NAND_GATE U3602 ( .I1(n2399), .I2(n2398), .O(n2400) );
  NAND_GATE U3603 ( .I1(n2401), .I2(n2400), .O(n2402) );
  NAND_GATE U3604 ( .I1(n2403), .I2(n2402), .O(n2404) );
  NAND_GATE U3605 ( .I1(n2405), .I2(n2404), .O(n2439) );
  NAND_GATE U3606 ( .I1(n2406), .I2(n2439), .O(n2435) );
  NAND_GATE U3607 ( .I1(n2440), .I2(n2439), .O(n2407) );
  NAND3_GATE U3608 ( .I1(n2436), .I2(n2435), .I3(n2407), .O(n2429) );
  NAND_GATE U3609 ( .I1(n2429), .I2(n2428), .O(n2409) );
  NAND_GATE U3610 ( .I1(n2408), .I2(n2429), .O(n2425) );
  AND3_GATE U3611 ( .I1(n2424), .I2(n2409), .I3(n2425), .O(n2420) );
  NAND_GATE U3612 ( .I1(n1440), .I2(A[31]), .O(n2419) );
  NAND_GATE U3613 ( .I1(n2420), .I2(n2419), .O(n2410) );
  NAND_GATE U3614 ( .I1(n2418), .I2(n2410), .O(n2423) );
  INV_GATE U3615 ( .I1(n2413), .O(n2411) );
  NAND_GATE U3616 ( .I1(n2412), .I2(n2411), .O(n2416) );
  INV_GATE U3617 ( .I1(n2412), .O(n2414) );
  NAND_GATE U3618 ( .I1(n2414), .I2(n2413), .O(n2415) );
  NAND_GATE U3619 ( .I1(n2423), .I2(n409), .O(n2417) );
  AND_GATE U3620 ( .I1(n14783), .I2(n2417), .O(\A1[58] ) );
  INV_GATE U3621 ( .I1(n2418), .O(n2421) );
  NAND3_GATE U3622 ( .I1(n2421), .I2(n2420), .I3(n2419), .O(n2422) );
  NAND_GATE U3623 ( .I1(n2423), .I2(n2422), .O(n2806) );
  INV_GATE U3624 ( .I1(n2806), .O(n14785) );
  OR_GATE U3625 ( .I1(n2424), .I2(n2429), .O(n2427) );
  OR_GATE U3626 ( .I1(n2428), .I2(n2425), .O(n2426) );
  AND_GATE U3627 ( .I1(n2427), .I2(n2426), .O(n2434) );
  NAND_GATE U3628 ( .I1(n2429), .I2(n1206), .O(n2431) );
  NAND3_GATE U3629 ( .I1(n2432), .I2(n2431), .I3(n2430), .O(n2433) );
  OR_GATE U3630 ( .I1(n2435), .I2(n2440), .O(n2438) );
  OR_GATE U3631 ( .I1(n2439), .I2(n2436), .O(n2437) );
  AND_GATE U3632 ( .I1(n2438), .I2(n2437), .O(n2445) );
  NAND_GATE U3633 ( .I1(n1205), .I2(n2439), .O(n2443) );
  NAND3_GATE U3634 ( .I1(n2443), .I2(n2442), .I3(n2441), .O(n2444) );
  NAND_GATE U3635 ( .I1(n2445), .I2(n2444), .O(n2814) );
  INV_GATE U3636 ( .I1(n2814), .O(n2817) );
  NAND_GATE U3637 ( .I1(B[27]), .I2(A[30]), .O(n2821) );
  INV_GATE U3638 ( .I1(n2821), .O(n2815) );
  NAND_GATE U3639 ( .I1(n2817), .I2(n2815), .O(n2812) );
  OR_GATE U3640 ( .I1(n2446), .I2(n2451), .O(n2449) );
  OR_GATE U3641 ( .I1(n2450), .I2(n2447), .O(n2448) );
  AND_GATE U3642 ( .I1(n2449), .I2(n2448), .O(n2456) );
  NAND_GATE U3643 ( .I1(n2451), .I2(n1204), .O(n2453) );
  NAND3_GATE U3644 ( .I1(n2454), .I2(n2453), .I3(n2452), .O(n2455) );
  NAND_GATE U3645 ( .I1(n2456), .I2(n2455), .O(n2828) );
  INV_GATE U3646 ( .I1(n2828), .O(n2831) );
  NAND_GATE U3647 ( .I1(B[27]), .I2(A[29]), .O(n2835) );
  INV_GATE U3648 ( .I1(n2835), .O(n2829) );
  NAND_GATE U3649 ( .I1(n2831), .I2(n2829), .O(n2826) );
  NAND_GATE U3650 ( .I1(B[27]), .I2(A[28]), .O(n3257) );
  INV_GATE U3651 ( .I1(n3257), .O(n3251) );
  OR_GATE U3652 ( .I1(n2457), .I2(n2462), .O(n2460) );
  OR_GATE U3653 ( .I1(n2461), .I2(n2458), .O(n2459) );
  AND_GATE U3654 ( .I1(n2460), .I2(n2459), .O(n2467) );
  NAND_GATE U3655 ( .I1(n2462), .I2(n1201), .O(n2464) );
  NAND3_GATE U3656 ( .I1(n2465), .I2(n2464), .I3(n2463), .O(n2466) );
  NAND_GATE U3657 ( .I1(n2467), .I2(n2466), .O(n3234) );
  INV_GATE U3658 ( .I1(n3234), .O(n3237) );
  NAND_GATE U3659 ( .I1(B[27]), .I2(A[27]), .O(n3241) );
  INV_GATE U3660 ( .I1(n3241), .O(n3235) );
  NAND_GATE U3661 ( .I1(n3237), .I2(n3235), .O(n3232) );
  OR_GATE U3662 ( .I1(n2468), .I2(n2473), .O(n2471) );
  OR_GATE U3663 ( .I1(n2472), .I2(n2469), .O(n2470) );
  AND_GATE U3664 ( .I1(n2471), .I2(n2470), .O(n2478) );
  NAND_GATE U3665 ( .I1(n1198), .I2(n2472), .O(n2476) );
  NAND3_GATE U3666 ( .I1(n2476), .I2(n2475), .I3(n2474), .O(n2477) );
  NAND_GATE U3667 ( .I1(n2478), .I2(n2477), .O(n2842) );
  INV_GATE U3668 ( .I1(n2842), .O(n2845) );
  NAND_GATE U3669 ( .I1(B[27]), .I2(A[26]), .O(n2849) );
  INV_GATE U3670 ( .I1(n2849), .O(n2843) );
  NAND_GATE U3671 ( .I1(n2845), .I2(n2843), .O(n2840) );
  OR_GATE U3672 ( .I1(n2479), .I2(n2484), .O(n2482) );
  OR_GATE U3673 ( .I1(n2483), .I2(n2480), .O(n2481) );
  AND_GATE U3674 ( .I1(n2482), .I2(n2481), .O(n2489) );
  NAND_GATE U3675 ( .I1(n2484), .I2(n1194), .O(n2486) );
  NAND3_GATE U3676 ( .I1(n2487), .I2(n2486), .I3(n2485), .O(n2488) );
  NAND_GATE U3677 ( .I1(n2489), .I2(n2488), .O(n3216) );
  INV_GATE U3678 ( .I1(n3216), .O(n3219) );
  NAND_GATE U3679 ( .I1(B[27]), .I2(A[25]), .O(n3223) );
  INV_GATE U3680 ( .I1(n3223), .O(n3217) );
  NAND_GATE U3681 ( .I1(n3219), .I2(n3217), .O(n3214) );
  OR_GATE U3682 ( .I1(n2490), .I2(n2495), .O(n2493) );
  OR_GATE U3683 ( .I1(n2494), .I2(n2491), .O(n2492) );
  AND_GATE U3684 ( .I1(n2493), .I2(n2492), .O(n2500) );
  NAND_GATE U3685 ( .I1(n1185), .I2(n2494), .O(n2498) );
  NAND3_GATE U3686 ( .I1(n2498), .I2(n2497), .I3(n2496), .O(n2499) );
  NAND_GATE U3687 ( .I1(n2500), .I2(n2499), .O(n3200) );
  INV_GATE U3688 ( .I1(n3200), .O(n3203) );
  NAND_GATE U3689 ( .I1(B[27]), .I2(A[24]), .O(n3207) );
  INV_GATE U3690 ( .I1(n3207), .O(n3201) );
  NAND_GATE U3691 ( .I1(n3203), .I2(n3201), .O(n3198) );
  OR_GATE U3692 ( .I1(n2501), .I2(n2506), .O(n2504) );
  OR_GATE U3693 ( .I1(n2505), .I2(n2502), .O(n2503) );
  AND_GATE U3694 ( .I1(n2504), .I2(n2503), .O(n2511) );
  NAND_GATE U3695 ( .I1(n2506), .I2(n1183), .O(n2508) );
  NAND3_GATE U3696 ( .I1(n2509), .I2(n2508), .I3(n2507), .O(n2510) );
  NAND_GATE U3697 ( .I1(n2511), .I2(n2510), .O(n3184) );
  INV_GATE U3698 ( .I1(n3184), .O(n3187) );
  NAND_GATE U3699 ( .I1(B[27]), .I2(A[23]), .O(n3191) );
  INV_GATE U3700 ( .I1(n3191), .O(n3185) );
  NAND_GATE U3701 ( .I1(n3187), .I2(n3185), .O(n3182) );
  OR_GATE U3702 ( .I1(n2512), .I2(n2517), .O(n2515) );
  OR_GATE U3703 ( .I1(n2516), .I2(n2513), .O(n2514) );
  AND_GATE U3704 ( .I1(n2515), .I2(n2514), .O(n2522) );
  NAND_GATE U3705 ( .I1(n1180), .I2(n2516), .O(n2520) );
  NAND3_GATE U3706 ( .I1(n2520), .I2(n2519), .I3(n2518), .O(n2521) );
  NAND_GATE U3707 ( .I1(n2522), .I2(n2521), .O(n3168) );
  INV_GATE U3708 ( .I1(n3168), .O(n3171) );
  NAND_GATE U3709 ( .I1(B[27]), .I2(A[22]), .O(n3175) );
  INV_GATE U3710 ( .I1(n3175), .O(n3169) );
  NAND_GATE U3711 ( .I1(n3171), .I2(n3169), .O(n3166) );
  OR_GATE U3712 ( .I1(n2523), .I2(n2528), .O(n2526) );
  OR_GATE U3713 ( .I1(n2527), .I2(n2524), .O(n2525) );
  AND_GATE U3714 ( .I1(n2526), .I2(n2525), .O(n2533) );
  NAND_GATE U3715 ( .I1(n2528), .I2(n1171), .O(n2530) );
  NAND3_GATE U3716 ( .I1(n2531), .I2(n2530), .I3(n2529), .O(n2532) );
  NAND_GATE U3717 ( .I1(n2533), .I2(n2532), .O(n3152) );
  INV_GATE U3718 ( .I1(n3152), .O(n3155) );
  NAND_GATE U3719 ( .I1(B[27]), .I2(A[21]), .O(n3159) );
  INV_GATE U3720 ( .I1(n3159), .O(n3153) );
  NAND_GATE U3721 ( .I1(n3155), .I2(n3153), .O(n3150) );
  OR_GATE U3722 ( .I1(n2534), .I2(n2539), .O(n2537) );
  OR_GATE U3723 ( .I1(n2538), .I2(n2535), .O(n2536) );
  AND_GATE U3724 ( .I1(n2537), .I2(n2536), .O(n2544) );
  NAND_GATE U3725 ( .I1(n1168), .I2(n2538), .O(n2542) );
  NAND3_GATE U3726 ( .I1(n2542), .I2(n2541), .I3(n2540), .O(n2543) );
  NAND_GATE U3727 ( .I1(n2544), .I2(n2543), .O(n3136) );
  INV_GATE U3728 ( .I1(n3136), .O(n3139) );
  NAND_GATE U3729 ( .I1(B[27]), .I2(A[20]), .O(n3143) );
  INV_GATE U3730 ( .I1(n3143), .O(n3137) );
  NAND_GATE U3731 ( .I1(n3139), .I2(n3137), .O(n3134) );
  OR_GATE U3732 ( .I1(n2545), .I2(n2550), .O(n2548) );
  OR_GATE U3733 ( .I1(n2549), .I2(n2546), .O(n2547) );
  NAND_GATE U3734 ( .I1(n2550), .I2(n1156), .O(n2552) );
  NAND3_GATE U3735 ( .I1(n2553), .I2(n2552), .I3(n2551), .O(n2554) );
  INV_GATE U3736 ( .I1(n3120), .O(n3123) );
  NAND_GATE U3737 ( .I1(B[27]), .I2(A[19]), .O(n3127) );
  INV_GATE U3738 ( .I1(n3127), .O(n3121) );
  NAND_GATE U3739 ( .I1(n3123), .I2(n3121), .O(n3118) );
  OR_GATE U3740 ( .I1(n2555), .I2(n2560), .O(n2558) );
  OR_GATE U3741 ( .I1(n2559), .I2(n2556), .O(n2557) );
  AND_GATE U3742 ( .I1(n2558), .I2(n2557), .O(n2565) );
  NAND_GATE U3743 ( .I1(n1133), .I2(n2559), .O(n2563) );
  NAND3_GATE U3744 ( .I1(n2563), .I2(n2562), .I3(n2561), .O(n2564) );
  NAND_GATE U3745 ( .I1(n2565), .I2(n2564), .O(n3104) );
  INV_GATE U3746 ( .I1(n3104), .O(n3107) );
  NAND_GATE U3747 ( .I1(B[27]), .I2(A[18]), .O(n3111) );
  INV_GATE U3748 ( .I1(n3111), .O(n3105) );
  NAND_GATE U3749 ( .I1(n3107), .I2(n3105), .O(n3102) );
  OR_GATE U3750 ( .I1(n2566), .I2(n2571), .O(n2569) );
  OR_GATE U3751 ( .I1(n2570), .I2(n2567), .O(n2568) );
  AND_GATE U3752 ( .I1(n2569), .I2(n2568), .O(n2576) );
  NAND_GATE U3753 ( .I1(n2571), .I2(n1132), .O(n2573) );
  NAND3_GATE U3754 ( .I1(n2574), .I2(n2573), .I3(n2572), .O(n2575) );
  NAND_GATE U3755 ( .I1(n2576), .I2(n2575), .O(n3088) );
  INV_GATE U3756 ( .I1(n3088), .O(n3091) );
  NAND_GATE U3757 ( .I1(B[27]), .I2(A[17]), .O(n3095) );
  INV_GATE U3758 ( .I1(n3095), .O(n3089) );
  NAND_GATE U3759 ( .I1(n3091), .I2(n3089), .O(n3086) );
  OR_GATE U3760 ( .I1(n2577), .I2(n2582), .O(n2580) );
  OR_GATE U3761 ( .I1(n2581), .I2(n2578), .O(n2579) );
  AND_GATE U3762 ( .I1(n2580), .I2(n2579), .O(n2587) );
  NAND_GATE U3763 ( .I1(n1131), .I2(n2581), .O(n2585) );
  NAND3_GATE U3764 ( .I1(n2585), .I2(n2584), .I3(n2583), .O(n2586) );
  NAND_GATE U3765 ( .I1(n2587), .I2(n2586), .O(n3072) );
  INV_GATE U3766 ( .I1(n3072), .O(n3075) );
  NAND_GATE U3767 ( .I1(B[27]), .I2(A[16]), .O(n3079) );
  INV_GATE U3768 ( .I1(n3079), .O(n3073) );
  NAND_GATE U3769 ( .I1(n3075), .I2(n3073), .O(n3070) );
  OR_GATE U3770 ( .I1(n2588), .I2(n2593), .O(n2591) );
  OR_GATE U3771 ( .I1(n2592), .I2(n2589), .O(n2590) );
  AND_GATE U3772 ( .I1(n2591), .I2(n2590), .O(n2598) );
  NAND_GATE U3773 ( .I1(n2593), .I2(n1152), .O(n2595) );
  NAND3_GATE U3774 ( .I1(n2596), .I2(n2595), .I3(n2594), .O(n2597) );
  NAND_GATE U3775 ( .I1(n2598), .I2(n2597), .O(n3056) );
  INV_GATE U3776 ( .I1(n3056), .O(n3059) );
  NAND_GATE U3777 ( .I1(B[27]), .I2(A[15]), .O(n3063) );
  INV_GATE U3778 ( .I1(n3063), .O(n3057) );
  NAND_GATE U3779 ( .I1(n3059), .I2(n3057), .O(n3054) );
  OR_GATE U3780 ( .I1(n2599), .I2(n2604), .O(n2602) );
  OR_GATE U3781 ( .I1(n2603), .I2(n2600), .O(n2601) );
  AND_GATE U3782 ( .I1(n2602), .I2(n2601), .O(n2609) );
  NAND_GATE U3783 ( .I1(n1153), .I2(n2603), .O(n2607) );
  NAND3_GATE U3784 ( .I1(n2607), .I2(n2606), .I3(n2605), .O(n2608) );
  NAND_GATE U3785 ( .I1(B[27]), .I2(A[14]), .O(n3047) );
  INV_GATE U3786 ( .I1(n3047), .O(n3042) );
  NAND_GATE U3787 ( .I1(n823), .I2(n3042), .O(n3039) );
  OR_GATE U3788 ( .I1(n2610), .I2(n2615), .O(n2613) );
  OR_GATE U3789 ( .I1(n2614), .I2(n2611), .O(n2612) );
  AND_GATE U3790 ( .I1(n2613), .I2(n2612), .O(n2620) );
  NAND_GATE U3791 ( .I1(n2615), .I2(n1154), .O(n2617) );
  NAND3_GATE U3792 ( .I1(n2618), .I2(n2617), .I3(n2616), .O(n2619) );
  NAND_GATE U3793 ( .I1(n2620), .I2(n2619), .O(n3025) );
  INV_GATE U3794 ( .I1(n3025), .O(n3028) );
  NAND_GATE U3795 ( .I1(B[27]), .I2(A[13]), .O(n3032) );
  INV_GATE U3796 ( .I1(n3032), .O(n3026) );
  NAND_GATE U3797 ( .I1(n3028), .I2(n3026), .O(n3023) );
  OR_GATE U3798 ( .I1(n2621), .I2(n2626), .O(n2624) );
  OR_GATE U3799 ( .I1(n2625), .I2(n2622), .O(n2623) );
  AND_GATE U3800 ( .I1(n2624), .I2(n2623), .O(n2631) );
  NAND_GATE U3801 ( .I1(n1130), .I2(n2625), .O(n2629) );
  NAND3_GATE U3802 ( .I1(n2629), .I2(n2628), .I3(n2627), .O(n2630) );
  NAND_GATE U3803 ( .I1(n2631), .I2(n2630), .O(n3013) );
  NAND_GATE U3804 ( .I1(B[27]), .I2(A[12]), .O(n3016) );
  INV_GATE U3805 ( .I1(n3016), .O(n3011) );
  NAND_GATE U3806 ( .I1(n368), .I2(n3011), .O(n3008) );
  OR_GATE U3807 ( .I1(n2632), .I2(n2637), .O(n2635) );
  OR_GATE U3808 ( .I1(n2636), .I2(n2633), .O(n2634) );
  NAND_GATE U3809 ( .I1(n2637), .I2(n1106), .O(n2639) );
  NAND3_GATE U3810 ( .I1(n2640), .I2(n2639), .I3(n2638), .O(n2641) );
  INV_GATE U3811 ( .I1(n2999), .O(n2997) );
  NAND_GATE U3812 ( .I1(B[27]), .I2(A[11]), .O(n3001) );
  INV_GATE U3813 ( .I1(n3001), .O(n2995) );
  NAND_GATE U3814 ( .I1(n2997), .I2(n2995), .O(n2992) );
  NAND_GATE U3815 ( .I1(n1105), .I2(n2648), .O(n2643) );
  NAND3_GATE U3816 ( .I1(n2644), .I2(n2643), .I3(n2642), .O(n2651) );
  OR_GATE U3817 ( .I1(n2646), .I2(n2645), .O(n2650) );
  OR_GATE U3818 ( .I1(n2648), .I2(n2647), .O(n2649) );
  NAND3_GATE U3819 ( .I1(n2651), .I2(n2650), .I3(n2649), .O(n2980) );
  INV_GATE U3820 ( .I1(n2980), .O(n2984) );
  NAND_GATE U3821 ( .I1(B[27]), .I2(A[10]), .O(n2982) );
  INV_GATE U3822 ( .I1(n2982), .O(n2981) );
  NAND_GATE U3823 ( .I1(n2984), .I2(n2981), .O(n2978) );
  OR_GATE U3824 ( .I1(n2657), .I2(n2652), .O(n2655) );
  NAND3_GATE U3825 ( .I1(n2653), .I2(n319), .I3(n2657), .O(n2654) );
  AND_GATE U3826 ( .I1(n2655), .I2(n2654), .O(n2662) );
  NAND_GATE U3827 ( .I1(n319), .I2(n2657), .O(n2659) );
  NAND3_GATE U3828 ( .I1(n2660), .I2(n2659), .I3(n2658), .O(n2661) );
  NAND_GATE U3829 ( .I1(n2662), .I2(n2661), .O(n2855) );
  INV_GATE U3830 ( .I1(n2855), .O(n2854) );
  NAND_GATE U3831 ( .I1(B[27]), .I2(A[9]), .O(n2856) );
  INV_GATE U3832 ( .I1(n2856), .O(n2857) );
  NAND_GATE U3833 ( .I1(n2854), .I2(n2857), .O(n2861) );
  NAND_GATE U3834 ( .I1(n2670), .I2(n840), .O(n2666) );
  INV_GATE U3835 ( .I1(n2670), .O(n2664) );
  NAND_GATE U3836 ( .I1(n2664), .I2(n2663), .O(n2665) );
  NAND3_GATE U3837 ( .I1(n2667), .I2(n2666), .I3(n2665), .O(n2673) );
  OR_GATE U3838 ( .I1(n2668), .I2(n2670), .O(n2672) );
  NAND3_GATE U3839 ( .I1(n840), .I2(n2670), .I3(n2669), .O(n2671) );
  NAND3_GATE U3840 ( .I1(n2673), .I2(n2672), .I3(n2671), .O(n2966) );
  INV_GATE U3841 ( .I1(n2966), .O(n2964) );
  NAND_GATE U3842 ( .I1(B[27]), .I2(A[8]), .O(n2965) );
  INV_GATE U3843 ( .I1(n2965), .O(n2963) );
  NAND_GATE U3844 ( .I1(n2964), .I2(n2963), .O(n2970) );
  NAND_GATE U3845 ( .I1(n897), .I2(n2680), .O(n2676) );
  NAND3_GATE U3846 ( .I1(n2677), .I2(n2676), .I3(n2675), .O(n2683) );
  OR_GATE U3847 ( .I1(n2680), .I2(n2678), .O(n2682) );
  NAND3_GATE U3848 ( .I1(n897), .I2(n2680), .I3(n2679), .O(n2681) );
  NAND3_GATE U3849 ( .I1(n2683), .I2(n2682), .I3(n2681), .O(n2867) );
  NAND_GATE U3850 ( .I1(B[27]), .I2(A[7]), .O(n2866) );
  INV_GATE U3851 ( .I1(n2866), .O(n2869) );
  NAND_GATE U3852 ( .I1(n812), .I2(n2869), .O(n2870) );
  NAND_GATE U3853 ( .I1(B[27]), .I2(A[6]), .O(n2942) );
  INV_GATE U3854 ( .I1(n2942), .O(n2953) );
  NAND3_GATE U3855 ( .I1(n2688), .I2(n2684), .I3(n2687), .O(n2686) );
  NAND3_GATE U3856 ( .I1(n2689), .I2(n2684), .I3(n896), .O(n2685) );
  AND_GATE U3857 ( .I1(n2686), .I2(n2685), .O(n2940) );
  NAND_GATE U3858 ( .I1(n2688), .I2(n2687), .O(n2692) );
  NAND_GATE U3859 ( .I1(n2689), .I2(n896), .O(n2691) );
  NAND3_GATE U3860 ( .I1(n2692), .I2(n2691), .I3(n2690), .O(n2939) );
  NAND_GATE U3861 ( .I1(n2940), .I2(n2939), .O(n2950) );
  NAND_GATE U3862 ( .I1(n2953), .I2(n348), .O(n2946) );
  NAND_GATE U3863 ( .I1(B[27]), .I2(A[5]), .O(n2935) );
  INV_GATE U3864 ( .I1(n2935), .O(n2881) );
  NAND_GATE U3865 ( .I1(B[27]), .I2(A[4]), .O(n2923) );
  INV_GATE U3866 ( .I1(n2923), .O(n2930) );
  OR_GATE U3867 ( .I1(n2694), .I2(n2693), .O(n2695) );
  NAND_GATE U3868 ( .I1(n2696), .I2(n2695), .O(n2705) );
  OR_GATE U3869 ( .I1(n2705), .I2(n2697), .O(n2703) );
  NAND5_GATE U3870 ( .I1(n2701), .I2(n2700), .I3(n2699), .I4(n2698), .I5(n1225), .O(n2702) );
  NAND_GATE U3871 ( .I1(n2703), .I2(n2702), .O(n2709) );
  NAND_GATE U3872 ( .I1(n1225), .I2(n2705), .O(n2707) );
  NAND_GATE U3873 ( .I1(n2930), .I2(n1397), .O(n2732) );
  NAND3_GATE U3874 ( .I1(n2708), .I2(n2923), .I3(n2707), .O(n2730) );
  NAND_GATE U3875 ( .I1(n2923), .I2(n2709), .O(n2729) );
  NAND_GATE U3876 ( .I1(B[27]), .I2(A[3]), .O(n2897) );
  INV_GATE U3877 ( .I1(n2897), .O(n2886) );
  NAND3_GATE U3878 ( .I1(B[27]), .I2(B[28]), .I3(n1254), .O(n2913) );
  INV_GATE U3879 ( .I1(n2913), .O(n2911) );
  NAND_GATE U3880 ( .I1(n1440), .I2(A[0]), .O(n2710) );
  NAND_GATE U3881 ( .I1(n14241), .I2(n2710), .O(n2711) );
  NAND_GATE U3882 ( .I1(B[29]), .I2(n2711), .O(n2907) );
  NAND_GATE U3883 ( .I1(B[28]), .I2(n2712), .O(n2908) );
  NAND_GATE U3884 ( .I1(B[27]), .I2(A[2]), .O(n2912) );
  NAND_GATE U3885 ( .I1(n915), .I2(n2912), .O(n2713) );
  NAND_GATE U3886 ( .I1(n2911), .I2(n2713), .O(n2715) );
  INV_GATE U3887 ( .I1(n2912), .O(n2910) );
  NAND_GATE U3888 ( .I1(n285), .I2(n2910), .O(n2714) );
  NAND_GATE U3889 ( .I1(n2715), .I2(n2714), .O(n2890) );
  NAND_GATE U3890 ( .I1(n2886), .I2(n2890), .O(n2889) );
  NAND3_GATE U3891 ( .I1(n2719), .I2(n2717), .I3(n2716), .O(n2718) );
  NAND_GATE U3892 ( .I1(n2724), .I2(n2718), .O(n2887) );
  NAND3_GATE U3893 ( .I1(n2720), .I2(n2723), .I3(n1281), .O(n2722) );
  NAND3_GATE U3894 ( .I1(n2720), .I2(n2719), .I3(n1339), .O(n2721) );
  AND_GATE U3895 ( .I1(n2722), .I2(n2721), .O(n2888) );
  NAND3_GATE U3896 ( .I1(n2886), .I2(n2887), .I3(n2888), .O(n2728) );
  INV_GATE U3897 ( .I1(n2887), .O(n2725) );
  NAND3_GATE U3898 ( .I1(n2724), .I2(n2723), .I3(n1281), .O(n2891) );
  NAND_GATE U3899 ( .I1(n2725), .I2(n2891), .O(n2726) );
  NAND3_GATE U3900 ( .I1(n2890), .I2(n2726), .I3(n2888), .O(n2727) );
  NAND3_GATE U3901 ( .I1(n2889), .I2(n2728), .I3(n2727), .O(n2922) );
  NAND3_GATE U3902 ( .I1(n2730), .I2(n2729), .I3(n2922), .O(n2731) );
  NAND_GATE U3903 ( .I1(n2732), .I2(n2731), .O(n2885) );
  NAND_GATE U3904 ( .I1(n2881), .I2(n2885), .O(n2952) );
  INV_GATE U3905 ( .I1(n2737), .O(n2734) );
  NAND_GATE U3906 ( .I1(n2735), .I2(n2734), .O(n2733) );
  NAND_GATE U3907 ( .I1(n1269), .I2(n2737), .O(n2744) );
  NAND3_GATE U3908 ( .I1(n2738), .I2(n2733), .I3(n2744), .O(n2880) );
  NAND3_GATE U3909 ( .I1(n2735), .I2(n2736), .I3(n2734), .O(n2742) );
  NAND3_GATE U3910 ( .I1(n907), .I2(n2736), .I3(n2737), .O(n2739) );
  NAND3_GATE U3911 ( .I1(n2880), .I2(n1211), .I3(n2881), .O(n2951) );
  NAND_GATE U3912 ( .I1(n2738), .I2(n2737), .O(n2741) );
  NAND4_GATE U3913 ( .I1(n2742), .I2(n2741), .I3(n2740), .I4(n2739), .O(n2743)
         );
  NAND_GATE U3914 ( .I1(n2744), .I2(n2743), .O(n2884) );
  NAND_GATE U3915 ( .I1(n2885), .I2(n2884), .O(n2949) );
  NAND3_GATE U3916 ( .I1(n2952), .I2(n2951), .I3(n2949), .O(n2947) );
  NAND_GATE U3917 ( .I1(n2942), .I2(n2950), .O(n2745) );
  NAND_GATE U3918 ( .I1(n2947), .I2(n2745), .O(n2746) );
  NAND_GATE U3919 ( .I1(n2966), .I2(n2965), .O(n2748) );
  NAND_GATE U3920 ( .I1(n1265), .I2(n2748), .O(n2749) );
  NAND_GATE U3921 ( .I1(n2970), .I2(n2749), .O(n2862) );
  NAND_GATE U3922 ( .I1(n2855), .I2(n2856), .O(n2750) );
  NAND_GATE U3923 ( .I1(n2862), .I2(n2750), .O(n2751) );
  NAND_GATE U3924 ( .I1(n2861), .I2(n2751), .O(n2983) );
  NAND_GATE U3925 ( .I1(n2980), .I2(n2982), .O(n2752) );
  NAND_GATE U3926 ( .I1(n2983), .I2(n2752), .O(n2753) );
  NAND_GATE U3927 ( .I1(n2978), .I2(n2753), .O(n2996) );
  NAND_GATE U3928 ( .I1(n2999), .I2(n3001), .O(n2754) );
  NAND_GATE U3929 ( .I1(n2996), .I2(n2754), .O(n2755) );
  NAND_GATE U3930 ( .I1(n2992), .I2(n2755), .O(n3012) );
  NAND_GATE U3931 ( .I1(n3013), .I2(n3016), .O(n2756) );
  NAND_GATE U3932 ( .I1(n3012), .I2(n2756), .O(n2757) );
  NAND_GATE U3933 ( .I1(n3008), .I2(n2757), .O(n3027) );
  NAND_GATE U3934 ( .I1(n3025), .I2(n3032), .O(n2758) );
  NAND_GATE U3935 ( .I1(n3027), .I2(n2758), .O(n2759) );
  NAND_GATE U3936 ( .I1(n3023), .I2(n2759), .O(n3043) );
  NAND_GATE U3937 ( .I1(n3041), .I2(n3047), .O(n2760) );
  NAND_GATE U3938 ( .I1(n3043), .I2(n2760), .O(n2761) );
  NAND_GATE U3939 ( .I1(n3039), .I2(n2761), .O(n3058) );
  NAND_GATE U3940 ( .I1(n3056), .I2(n3063), .O(n2762) );
  NAND_GATE U3941 ( .I1(n3058), .I2(n2762), .O(n2763) );
  NAND_GATE U3942 ( .I1(n3054), .I2(n2763), .O(n3074) );
  NAND_GATE U3943 ( .I1(n3072), .I2(n3079), .O(n2764) );
  NAND_GATE U3944 ( .I1(n3074), .I2(n2764), .O(n2765) );
  NAND_GATE U3945 ( .I1(n3070), .I2(n2765), .O(n3090) );
  NAND_GATE U3946 ( .I1(n3088), .I2(n3095), .O(n2766) );
  NAND_GATE U3947 ( .I1(n3090), .I2(n2766), .O(n2767) );
  NAND_GATE U3948 ( .I1(n3086), .I2(n2767), .O(n3106) );
  NAND_GATE U3949 ( .I1(n3104), .I2(n3111), .O(n2768) );
  NAND_GATE U3950 ( .I1(n3106), .I2(n2768), .O(n2769) );
  NAND_GATE U3951 ( .I1(n3102), .I2(n2769), .O(n3122) );
  NAND_GATE U3952 ( .I1(n3120), .I2(n3127), .O(n2770) );
  NAND_GATE U3953 ( .I1(n3122), .I2(n2770), .O(n2771) );
  NAND_GATE U3954 ( .I1(n3118), .I2(n2771), .O(n3138) );
  NAND_GATE U3955 ( .I1(n3136), .I2(n3143), .O(n2772) );
  NAND_GATE U3956 ( .I1(n3138), .I2(n2772), .O(n2773) );
  NAND_GATE U3957 ( .I1(n3134), .I2(n2773), .O(n3154) );
  NAND_GATE U3958 ( .I1(n3152), .I2(n3159), .O(n2774) );
  NAND_GATE U3959 ( .I1(n3154), .I2(n2774), .O(n2775) );
  NAND_GATE U3960 ( .I1(n3150), .I2(n2775), .O(n3170) );
  NAND_GATE U3961 ( .I1(n3168), .I2(n3175), .O(n2776) );
  NAND_GATE U3962 ( .I1(n3170), .I2(n2776), .O(n2777) );
  NAND_GATE U3963 ( .I1(n3166), .I2(n2777), .O(n3186) );
  NAND_GATE U3964 ( .I1(n3184), .I2(n3191), .O(n2778) );
  NAND_GATE U3965 ( .I1(n3186), .I2(n2778), .O(n2779) );
  NAND_GATE U3966 ( .I1(n3182), .I2(n2779), .O(n3202) );
  NAND_GATE U3967 ( .I1(n3200), .I2(n3207), .O(n2780) );
  NAND_GATE U3968 ( .I1(n3202), .I2(n2780), .O(n2781) );
  NAND_GATE U3969 ( .I1(n3198), .I2(n2781), .O(n3218) );
  NAND_GATE U3970 ( .I1(n3216), .I2(n3223), .O(n2782) );
  NAND_GATE U3971 ( .I1(n3218), .I2(n2782), .O(n2783) );
  NAND_GATE U3972 ( .I1(n3214), .I2(n2783), .O(n2844) );
  NAND_GATE U3973 ( .I1(n2842), .I2(n2849), .O(n2784) );
  NAND_GATE U3974 ( .I1(n2844), .I2(n2784), .O(n2785) );
  NAND_GATE U3975 ( .I1(n2840), .I2(n2785), .O(n3236) );
  NAND_GATE U3976 ( .I1(n3234), .I2(n3241), .O(n2786) );
  NAND_GATE U3977 ( .I1(n3236), .I2(n2786), .O(n2787) );
  NAND_GATE U3978 ( .I1(n3232), .I2(n2787), .O(n3253) );
  NAND_GATE U3979 ( .I1(n3251), .I2(n3253), .O(n3248) );
  OR_GATE U3980 ( .I1(n2788), .I2(n2793), .O(n2791) );
  OR_GATE U3981 ( .I1(n2792), .I2(n2789), .O(n2790) );
  AND_GATE U3982 ( .I1(n2791), .I2(n2790), .O(n2798) );
  NAND_GATE U3983 ( .I1(n1202), .I2(n2792), .O(n2796) );
  NAND3_GATE U3984 ( .I1(n2796), .I2(n2795), .I3(n2794), .O(n2797) );
  NAND_GATE U3985 ( .I1(n2798), .I2(n2797), .O(n3249) );
  INV_GATE U3986 ( .I1(n3249), .O(n3252) );
  INV_GATE U3987 ( .I1(n3253), .O(n3250) );
  NAND_GATE U3988 ( .I1(n3257), .I2(n3250), .O(n2799) );
  NAND_GATE U3989 ( .I1(n3252), .I2(n2799), .O(n2800) );
  NAND_GATE U3990 ( .I1(n3248), .I2(n2800), .O(n2830) );
  NAND_GATE U3991 ( .I1(n2828), .I2(n2835), .O(n2801) );
  NAND_GATE U3992 ( .I1(n2830), .I2(n2801), .O(n2802) );
  NAND_GATE U3993 ( .I1(n2826), .I2(n2802), .O(n2816) );
  NAND_GATE U3994 ( .I1(n2814), .I2(n2821), .O(n2803) );
  NAND_GATE U3995 ( .I1(n2816), .I2(n2803), .O(n2805) );
  NAND_GATE U3996 ( .I1(n1439), .I2(A[31]), .O(n2804) );
  NAND3_GATE U3997 ( .I1(n2812), .I2(n2805), .I3(n2804), .O(n2809) );
  NAND_GATE U3998 ( .I1(n408), .I2(n2809), .O(n2811) );
  NAND_GATE U3999 ( .I1(n14785), .I2(n2811), .O(n2808) );
  INV_GATE U4000 ( .I1(n2811), .O(n14784) );
  NAND_GATE U4001 ( .I1(n2806), .I2(n14784), .O(n2807) );
  NAND_GATE U4002 ( .I1(n2808), .I2(n2807), .O(\A1[57] ) );
  NAND_GATE U4003 ( .I1(n2811), .I2(n2810), .O(n3267) );
  INV_GATE U4004 ( .I1(n3267), .O(n14787) );
  INV_GATE U4005 ( .I1(n2812), .O(n2813) );
  NAND_GATE U4006 ( .I1(n2813), .I2(n2816), .O(n2825) );
  NAND_GATE U4007 ( .I1(n2815), .I2(n2819), .O(n2823) );
  NAND_GATE U4008 ( .I1(n2817), .I2(n2816), .O(n2818) );
  NAND_GATE U4009 ( .I1(n2819), .I2(n2818), .O(n2820) );
  NAND_GATE U4010 ( .I1(n2821), .I2(n2820), .O(n2822) );
  NAND_GATE U4011 ( .I1(n2823), .I2(n2822), .O(n2824) );
  NAND_GATE U4012 ( .I1(n2825), .I2(n2824), .O(n3270) );
  NAND_GATE U4013 ( .I1(B[26]), .I2(A[30]), .O(n3282) );
  INV_GATE U4014 ( .I1(n3282), .O(n3264) );
  INV_GATE U4015 ( .I1(n2826), .O(n2827) );
  NAND_GATE U4016 ( .I1(n2827), .I2(n2830), .O(n2839) );
  NAND_GATE U4017 ( .I1(n2829), .I2(n2833), .O(n2837) );
  NAND_GATE U4018 ( .I1(n2831), .I2(n2830), .O(n2832) );
  NAND_GATE U4019 ( .I1(n2833), .I2(n2832), .O(n2834) );
  NAND_GATE U4020 ( .I1(n2835), .I2(n2834), .O(n2836) );
  NAND_GATE U4021 ( .I1(n2837), .I2(n2836), .O(n2838) );
  NAND_GATE U4022 ( .I1(n2839), .I2(n2838), .O(n3280) );
  NAND_GATE U4023 ( .I1(n3264), .I2(n3280), .O(n3276) );
  NAND_GATE U4024 ( .I1(B[26]), .I2(A[29]), .O(n3295) );
  INV_GATE U4025 ( .I1(n3295), .O(n3262) );
  NAND_GATE U4026 ( .I1(B[26]), .I2(A[28]), .O(n3306) );
  INV_GATE U4027 ( .I1(n3306), .O(n3246) );
  NAND_GATE U4028 ( .I1(B[26]), .I2(A[27]), .O(n3319) );
  INV_GATE U4029 ( .I1(n3319), .O(n3230) );
  INV_GATE U4030 ( .I1(n2840), .O(n2841) );
  NAND_GATE U4031 ( .I1(n2841), .I2(n2844), .O(n2853) );
  NAND_GATE U4032 ( .I1(n2843), .I2(n2847), .O(n2851) );
  NAND_GATE U4033 ( .I1(n2845), .I2(n2844), .O(n2846) );
  NAND_GATE U4034 ( .I1(n2847), .I2(n2846), .O(n2848) );
  NAND_GATE U4035 ( .I1(n2849), .I2(n2848), .O(n2850) );
  NAND_GATE U4036 ( .I1(n2851), .I2(n2850), .O(n2852) );
  NAND_GATE U4037 ( .I1(n2853), .I2(n2852), .O(n3316) );
  NAND_GATE U4038 ( .I1(n3230), .I2(n3316), .O(n3312) );
  NAND_GATE U4039 ( .I1(B[26]), .I2(A[26]), .O(n3330) );
  INV_GATE U4040 ( .I1(n3330), .O(n3228) );
  NAND_GATE U4041 ( .I1(B[26]), .I2(A[25]), .O(n3666) );
  INV_GATE U4042 ( .I1(n3666), .O(n3212) );
  NAND_GATE U4043 ( .I1(B[26]), .I2(A[24]), .O(n3341) );
  INV_GATE U4044 ( .I1(n3341), .O(n3196) );
  NAND_GATE U4045 ( .I1(B[26]), .I2(A[23]), .O(n3352) );
  INV_GATE U4046 ( .I1(n3352), .O(n3180) );
  NAND_GATE U4047 ( .I1(B[26]), .I2(A[22]), .O(n3363) );
  INV_GATE U4048 ( .I1(n3363), .O(n3164) );
  NAND_GATE U4049 ( .I1(B[26]), .I2(A[21]), .O(n3374) );
  INV_GATE U4050 ( .I1(n3374), .O(n3148) );
  NAND_GATE U4051 ( .I1(B[26]), .I2(A[20]), .O(n3385) );
  INV_GATE U4052 ( .I1(n3385), .O(n3132) );
  NAND_GATE U4053 ( .I1(B[26]), .I2(A[19]), .O(n3398) );
  INV_GATE U4054 ( .I1(n3398), .O(n3116) );
  NAND_GATE U4055 ( .I1(B[26]), .I2(A[18]), .O(n3409) );
  INV_GATE U4056 ( .I1(n3409), .O(n3100) );
  NAND_GATE U4057 ( .I1(B[26]), .I2(A[17]), .O(n3422) );
  INV_GATE U4058 ( .I1(n3422), .O(n3084) );
  NAND_GATE U4059 ( .I1(B[26]), .I2(A[16]), .O(n3433) );
  INV_GATE U4060 ( .I1(n3433), .O(n3068) );
  NAND_GATE U4061 ( .I1(B[26]), .I2(A[15]), .O(n3445) );
  INV_GATE U4062 ( .I1(n3445), .O(n3052) );
  NAND_GATE U4063 ( .I1(B[26]), .I2(A[14]), .O(n3456) );
  INV_GATE U4064 ( .I1(n3456), .O(n3037) );
  NAND_GATE U4065 ( .I1(B[26]), .I2(A[13]), .O(n3467) );
  INV_GATE U4066 ( .I1(n3467), .O(n3021) );
  NAND_GATE U4067 ( .I1(B[26]), .I2(A[12]), .O(n3478) );
  INV_GATE U4068 ( .I1(n3478), .O(n3006) );
  NAND_GATE U4069 ( .I1(B[26]), .I2(A[11]), .O(n3488) );
  INV_GATE U4070 ( .I1(n3488), .O(n2990) );
  NAND_GATE U4071 ( .I1(B[26]), .I2(A[10]), .O(n3493) );
  INV_GATE U4072 ( .I1(n3493), .O(n2976) );
  NAND_GATE U4073 ( .I1(n2854), .I2(n2862), .O(n2860) );
  NAND_GATE U4074 ( .I1(n2856), .I2(n1398), .O(n2859) );
  NAND3_GATE U4075 ( .I1(n2860), .I2(n2859), .I3(n2858), .O(n2865) );
  INV_GATE U4076 ( .I1(n2861), .O(n2863) );
  NAND_GATE U4077 ( .I1(n2863), .I2(n2862), .O(n2864) );
  NAND_GATE U4078 ( .I1(n2865), .I2(n2864), .O(n3498) );
  NAND_GATE U4079 ( .I1(n2976), .I2(n3498), .O(n3496) );
  NAND3_GATE U4080 ( .I1(n2867), .I2(n2866), .I3(n1375), .O(n2877) );
  NAND3_GATE U4081 ( .I1(n2866), .I2(n2871), .I3(n812), .O(n2876) );
  NAND_GATE U4082 ( .I1(B[26]), .I2(A[8]), .O(n3621) );
  INV_GATE U4083 ( .I1(n3621), .O(n3613) );
  AND3_GATE U4084 ( .I1(n2877), .I2(n2876), .I3(n3613), .O(n2874) );
  NAND_GATE U4085 ( .I1(n2867), .I2(n1375), .O(n2868) );
  NAND_GATE U4086 ( .I1(n2869), .I2(n2868), .O(n2875) );
  INV_GATE U4087 ( .I1(n2875), .O(n2872) );
  NAND_GATE U4088 ( .I1(n2872), .I2(n2879), .O(n2873) );
  NAND_GATE U4089 ( .I1(n2874), .I2(n2873), .O(n3614) );
  NAND3_GATE U4090 ( .I1(n2877), .I2(n2876), .I3(n2875), .O(n2878) );
  NAND_GATE U4091 ( .I1(n2879), .I2(n2878), .O(n3618) );
  NAND_GATE U4092 ( .I1(B[26]), .I2(A[7]), .O(n3516) );
  INV_GATE U4093 ( .I1(n3516), .O(n3518) );
  OR_GATE U4094 ( .I1(n2884), .I2(n2952), .O(n2883) );
  NAND4_GATE U4095 ( .I1(n2881), .I2(n2880), .I3(n1211), .I4(n326), .O(n2882)
         );
  NAND_GATE U4096 ( .I1(n326), .I2(n2884), .O(n2933) );
  NAND3_GATE U4097 ( .I1(n2933), .I2(n2934), .I3(n2935), .O(n3599) );
  NAND_GATE U4098 ( .I1(n1355), .I2(n3599), .O(n3590) );
  INV_GATE U4099 ( .I1(n3590), .O(n3593) );
  NAND_GATE U4100 ( .I1(B[26]), .I2(A[6]), .O(n3592) );
  INV_GATE U4101 ( .I1(n3592), .O(n3605) );
  NAND_GATE U4102 ( .I1(n3593), .I2(n3605), .O(n3589) );
  NAND_GATE U4103 ( .I1(B[26]), .I2(A[4]), .O(n3578) );
  INV_GATE U4104 ( .I1(n3578), .O(n3580) );
  INV_GATE U4105 ( .I1(n2890), .O(n2894) );
  NAND4_GATE U4106 ( .I1(n2886), .I2(n2887), .I3(n2888), .I4(n2894), .O(n2899)
         );
  NAND_GATE U4107 ( .I1(n2888), .I2(n2887), .O(n2892) );
  NAND_GATE U4108 ( .I1(n2891), .I2(n2892), .O(n2893) );
  OR_GATE U4109 ( .I1(n2893), .I2(n2889), .O(n2898) );
  NAND3_GATE U4110 ( .I1(n2892), .I2(n2891), .I3(n2890), .O(n2896) );
  NAND_GATE U4111 ( .I1(n2894), .I2(n2893), .O(n2895) );
  NAND3_GATE U4112 ( .I1(n2897), .I2(n2896), .I3(n2895), .O(n3573) );
  NAND3_GATE U4113 ( .I1(n2899), .I2(n2898), .I3(n3573), .O(n3576) );
  NAND_GATE U4114 ( .I1(n3580), .I2(n304), .O(n2920) );
  NAND_GATE U4115 ( .I1(B[26]), .I2(A[3]), .O(n3569) );
  INV_GATE U4116 ( .I1(n3569), .O(n3559) );
  NAND3_GATE U4117 ( .I1(B[26]), .I2(B[27]), .I3(n1254), .O(n3546) );
  INV_GATE U4118 ( .I1(n3546), .O(n3540) );
  NAND_GATE U4119 ( .I1(n1440), .I2(A[1]), .O(n2900) );
  NAND_GATE U4120 ( .I1(n724), .I2(n2900), .O(n2901) );
  NAND_GATE U4121 ( .I1(B[27]), .I2(n2901), .O(n3547) );
  NAND_GATE U4122 ( .I1(B[26]), .I2(A[2]), .O(n3541) );
  NAND_GATE U4123 ( .I1(n3547), .I2(n3541), .O(n2902) );
  NAND_GATE U4124 ( .I1(n3540), .I2(n2902), .O(n2906) );
  INV_GATE U4125 ( .I1(n3541), .O(n3550) );
  NAND_GATE U4126 ( .I1(n1439), .I2(A[0]), .O(n2903) );
  NAND_GATE U4127 ( .I1(n14241), .I2(n2903), .O(n2904) );
  NAND_GATE U4128 ( .I1(B[28]), .I2(n2904), .O(n3548) );
  NAND_GATE U4129 ( .I1(n3547), .I2(n3548), .O(n3542) );
  NAND_GATE U4130 ( .I1(n3550), .I2(n3542), .O(n2905) );
  NAND_GATE U4131 ( .I1(n2906), .I2(n2905), .O(n3562) );
  NAND_GATE U4132 ( .I1(n3559), .I2(n3562), .O(n3555) );
  NAND3_GATE U4133 ( .I1(n2908), .I2(n2907), .I3(n2913), .O(n2909) );
  NAND_GATE U4134 ( .I1(n2910), .I2(n2909), .O(n3556) );
  NAND3_GATE U4135 ( .I1(n285), .I2(n2910), .I3(n2911), .O(n3563) );
  NAND_GATE U4136 ( .I1(n1348), .I2(n3563), .O(n2915) );
  NAND3_GATE U4137 ( .I1(n2911), .I2(n2912), .I3(n285), .O(n3557) );
  NAND3_GATE U4138 ( .I1(n2913), .I2(n2912), .I3(n915), .O(n3558) );
  NAND_GATE U4139 ( .I1(n3557), .I2(n3558), .O(n2914) );
  INV_GATE U4140 ( .I1(n2914), .O(n3554) );
  NAND3_GATE U4141 ( .I1(n2915), .I2(n3554), .I3(n3562), .O(n2917) );
  NAND3_GATE U4142 ( .I1(n3559), .I2(n2915), .I3(n3554), .O(n2916) );
  NAND3_GATE U4143 ( .I1(n3555), .I2(n2917), .I3(n2916), .O(n3579) );
  NAND_GATE U4144 ( .I1(n3578), .I2(n3576), .O(n2918) );
  NAND_GATE U4145 ( .I1(n3579), .I2(n2918), .O(n2919) );
  NAND_GATE U4146 ( .I1(n2920), .I2(n2919), .O(n3524) );
  NAND_GATE U4147 ( .I1(n2930), .I2(n2922), .O(n2926) );
  INV_GATE U4148 ( .I1(n2926), .O(n2921) );
  NAND_GATE U4149 ( .I1(n1397), .I2(n2921), .O(n2928) );
  NAND3_GATE U4150 ( .I1(n2923), .I2(n2922), .I3(n1397), .O(n2932) );
  NAND3_GATE U4151 ( .I1(n331), .I2(n2924), .I3(n2930), .O(n2925) );
  NAND4_GATE U4152 ( .I1(n2932), .I2(n2931), .I3(n2926), .I4(n2925), .O(n2927)
         );
  NAND_GATE U4153 ( .I1(n2928), .I2(n2927), .O(n3531) );
  NAND_GATE U4154 ( .I1(n3524), .I2(n3531), .O(n3601) );
  NAND_GATE U4155 ( .I1(B[26]), .I2(A[5]), .O(n3527) );
  INV_GATE U4156 ( .I1(n3527), .O(n3530) );
  NAND3_GATE U4157 ( .I1(n2930), .I2(n2929), .I3(n2928), .O(n3529) );
  NAND3_GATE U4158 ( .I1(n3530), .I2(n3529), .I3(n1213), .O(n3597) );
  NAND_GATE U4159 ( .I1(n3530), .I2(n3524), .O(n3598) );
  NAND3_GATE U4160 ( .I1(n3601), .I2(n3597), .I3(n3598), .O(n3594) );
  NAND4_GATE U4161 ( .I1(n2935), .I2(n3592), .I3(n2934), .I4(n2933), .O(n2937)
         );
  NAND_GATE U4162 ( .I1(n3602), .I2(n3592), .O(n2936) );
  NAND3_GATE U4163 ( .I1(n3594), .I2(n2937), .I3(n2936), .O(n2938) );
  NAND_GATE U4164 ( .I1(n3589), .I2(n2938), .O(n3513) );
  NAND_GATE U4165 ( .I1(n3518), .I2(n3513), .O(n3519) );
  NAND3_GATE U4166 ( .I1(n2942), .I2(n348), .I3(n2947), .O(n2957) );
  NAND3_GATE U4167 ( .I1(n2940), .I2(n2939), .I3(n2953), .O(n2945) );
  INV_GATE U4168 ( .I1(n2947), .O(n2941) );
  NAND3_GATE U4169 ( .I1(n2942), .I2(n2950), .I3(n2941), .O(n2956) );
  NAND3_GATE U4170 ( .I1(n2949), .I2(n2951), .I3(n2952), .O(n2943) );
  NAND_GATE U4171 ( .I1(n2953), .I2(n2943), .O(n2944) );
  NAND4_GATE U4172 ( .I1(n2957), .I2(n2945), .I3(n2956), .I4(n2944), .O(n2948)
         );
  NAND_GATE U4173 ( .I1(n2948), .I2(n2954), .O(n3520) );
  NAND_GATE U4174 ( .I1(n3513), .I2(n3520), .O(n2959) );
  NAND4_GATE U4175 ( .I1(n2952), .I2(n2951), .I3(n2950), .I4(n2949), .O(n2955)
         );
  NAND3_GATE U4176 ( .I1(n2955), .I2(n2954), .I3(n2953), .O(n3517) );
  NAND3_GATE U4177 ( .I1(n3518), .I2(n3517), .I3(n1210), .O(n2958) );
  NAND3_GATE U4178 ( .I1(n3519), .I2(n2959), .I3(n2958), .O(n3617) );
  NAND_GATE U4179 ( .I1(n3618), .I2(n3617), .O(n2961) );
  NAND_GATE U4180 ( .I1(n3613), .I2(n3617), .O(n2960) );
  NAND3_GATE U4181 ( .I1(n3614), .I2(n2961), .I3(n2960), .O(n3506) );
  NAND_GATE U4182 ( .I1(n2966), .I2(n1371), .O(n2962) );
  NAND_GATE U4183 ( .I1(n2963), .I2(n2962), .O(n2969) );
  NAND_GATE U4184 ( .I1(n2964), .I2(n1265), .O(n2968) );
  NAND3_GATE U4185 ( .I1(n2966), .I2(n1371), .I3(n2965), .O(n2967) );
  NAND3_GATE U4186 ( .I1(n2969), .I2(n2968), .I3(n2967), .O(n2972) );
  NAND_GATE U4187 ( .I1(n2972), .I2(n2971), .O(n3507) );
  NAND_GATE U4188 ( .I1(n3506), .I2(n3507), .O(n2975) );
  NAND_GATE U4189 ( .I1(B[26]), .I2(A[9]), .O(n3508) );
  INV_GATE U4190 ( .I1(n3508), .O(n3503) );
  NAND_GATE U4191 ( .I1(n3503), .I2(n3507), .O(n2974) );
  NAND_GATE U4192 ( .I1(n3503), .I2(n3506), .O(n2973) );
  NAND3_GATE U4193 ( .I1(n2975), .I2(n2974), .I3(n2973), .O(n3497) );
  NAND_GATE U4194 ( .I1(n3498), .I2(n3497), .O(n2977) );
  NAND_GATE U4195 ( .I1(n2976), .I2(n3497), .O(n3499) );
  NAND3_GATE U4196 ( .I1(n3496), .I2(n2977), .I3(n3499), .O(n3487) );
  NAND_GATE U4197 ( .I1(n2990), .I2(n3487), .O(n3482) );
  INV_GATE U4198 ( .I1(n2978), .O(n2979) );
  NAND_GATE U4199 ( .I1(n2979), .I2(n2983), .O(n2989) );
  NAND_GATE U4200 ( .I1(n2982), .I2(n1391), .O(n2986) );
  NAND_GATE U4201 ( .I1(n2984), .I2(n2983), .O(n2985) );
  NAND3_GATE U4202 ( .I1(n2987), .I2(n2986), .I3(n2985), .O(n2988) );
  NAND_GATE U4203 ( .I1(n2989), .I2(n2988), .O(n3486) );
  NAND_GATE U4204 ( .I1(n2990), .I2(n3486), .O(n3483) );
  NAND_GATE U4205 ( .I1(n3487), .I2(n3486), .O(n2991) );
  NAND_GATE U4206 ( .I1(n3006), .I2(n3477), .O(n3473) );
  INV_GATE U4207 ( .I1(n2992), .O(n2993) );
  NAND_GATE U4208 ( .I1(n2993), .I2(n2996), .O(n3005) );
  INV_GATE U4209 ( .I1(n2996), .O(n2998) );
  NAND_GATE U4210 ( .I1(n2999), .I2(n2998), .O(n2994) );
  NAND_GATE U4211 ( .I1(n2995), .I2(n2994), .O(n3003) );
  NAND_GATE U4212 ( .I1(n2997), .I2(n2996), .O(n3000) );
  NAND_GATE U4213 ( .I1(n3003), .I2(n3002), .O(n3004) );
  NAND_GATE U4214 ( .I1(n3005), .I2(n3004), .O(n3476) );
  NAND_GATE U4215 ( .I1(n3006), .I2(n3476), .O(n3472) );
  NAND_GATE U4216 ( .I1(n3477), .I2(n3476), .O(n3007) );
  NAND3_GATE U4217 ( .I1(n3473), .I2(n3472), .I3(n3007), .O(n3466) );
  NAND_GATE U4218 ( .I1(n3021), .I2(n3466), .O(n3462) );
  INV_GATE U4219 ( .I1(n3008), .O(n3009) );
  NAND_GATE U4220 ( .I1(n3009), .I2(n3012), .O(n3020) );
  NAND_GATE U4221 ( .I1(n3013), .I2(n838), .O(n3010) );
  NAND_GATE U4222 ( .I1(n3011), .I2(n3010), .O(n3018) );
  NAND_GATE U4223 ( .I1(n368), .I2(n3012), .O(n3014) );
  NAND_GATE U4224 ( .I1(n3014), .I2(n3010), .O(n3015) );
  NAND_GATE U4225 ( .I1(n3016), .I2(n3015), .O(n3017) );
  NAND_GATE U4226 ( .I1(n3018), .I2(n3017), .O(n3019) );
  NAND_GATE U4227 ( .I1(n3020), .I2(n3019), .O(n3465) );
  NAND_GATE U4228 ( .I1(n3466), .I2(n3465), .O(n3022) );
  NAND3_GATE U4229 ( .I1(n3462), .I2(n3461), .I3(n3022), .O(n3455) );
  NAND_GATE U4230 ( .I1(n3037), .I2(n3455), .O(n3451) );
  INV_GATE U4231 ( .I1(n3023), .O(n3024) );
  NAND_GATE U4232 ( .I1(n3024), .I2(n3027), .O(n3036) );
  NAND_GATE U4233 ( .I1(n3026), .I2(n3030), .O(n3034) );
  NAND_GATE U4234 ( .I1(n3028), .I2(n3027), .O(n3029) );
  NAND_GATE U4235 ( .I1(n3030), .I2(n3029), .O(n3031) );
  NAND_GATE U4236 ( .I1(n3032), .I2(n3031), .O(n3033) );
  NAND_GATE U4237 ( .I1(n3034), .I2(n3033), .O(n3035) );
  NAND_GATE U4238 ( .I1(n3036), .I2(n3035), .O(n3454) );
  NAND_GATE U4239 ( .I1(n3037), .I2(n3454), .O(n3450) );
  NAND_GATE U4240 ( .I1(n3455), .I2(n3454), .O(n3038) );
  NAND3_GATE U4241 ( .I1(n3451), .I2(n3450), .I3(n3038), .O(n3444) );
  NAND_GATE U4242 ( .I1(n3052), .I2(n3444), .O(n3438) );
  INV_GATE U4243 ( .I1(n3039), .O(n3040) );
  NAND_GATE U4244 ( .I1(n3040), .I2(n3043), .O(n3051) );
  NAND_GATE U4245 ( .I1(n3042), .I2(n3045), .O(n3049) );
  NAND_GATE U4246 ( .I1(n823), .I2(n3043), .O(n3044) );
  NAND_GATE U4247 ( .I1(n3045), .I2(n3044), .O(n3046) );
  NAND_GATE U4248 ( .I1(n3047), .I2(n3046), .O(n3048) );
  NAND_GATE U4249 ( .I1(n3049), .I2(n3048), .O(n3050) );
  NAND_GATE U4250 ( .I1(n3051), .I2(n3050), .O(n3442) );
  NAND_GATE U4251 ( .I1(n3052), .I2(n3442), .O(n3437) );
  NAND_GATE U4252 ( .I1(n3444), .I2(n3442), .O(n3053) );
  NAND3_GATE U4253 ( .I1(n3438), .I2(n3437), .I3(n3053), .O(n3432) );
  NAND_GATE U4254 ( .I1(n3068), .I2(n3432), .O(n3428) );
  INV_GATE U4255 ( .I1(n3054), .O(n3055) );
  NAND_GATE U4256 ( .I1(n3055), .I2(n3058), .O(n3067) );
  NAND_GATE U4257 ( .I1(n3057), .I2(n3061), .O(n3065) );
  NAND_GATE U4258 ( .I1(n3059), .I2(n3058), .O(n3060) );
  NAND_GATE U4259 ( .I1(n3061), .I2(n3060), .O(n3062) );
  NAND_GATE U4260 ( .I1(n3063), .I2(n3062), .O(n3064) );
  NAND_GATE U4261 ( .I1(n3065), .I2(n3064), .O(n3066) );
  NAND_GATE U4262 ( .I1(n3067), .I2(n3066), .O(n3431) );
  NAND_GATE U4263 ( .I1(n3068), .I2(n3431), .O(n3427) );
  NAND_GATE U4264 ( .I1(n3432), .I2(n3431), .O(n3069) );
  NAND3_GATE U4265 ( .I1(n3428), .I2(n3427), .I3(n3069), .O(n3421) );
  NAND_GATE U4266 ( .I1(n3084), .I2(n3421), .O(n3415) );
  INV_GATE U4267 ( .I1(n3070), .O(n3071) );
  NAND_GATE U4268 ( .I1(n3071), .I2(n3074), .O(n3083) );
  NAND_GATE U4269 ( .I1(n3073), .I2(n3077), .O(n3081) );
  NAND_GATE U4270 ( .I1(n3075), .I2(n3074), .O(n3076) );
  NAND_GATE U4271 ( .I1(n3077), .I2(n3076), .O(n3078) );
  NAND_GATE U4272 ( .I1(n3079), .I2(n3078), .O(n3080) );
  NAND_GATE U4273 ( .I1(n3081), .I2(n3080), .O(n3082) );
  NAND_GATE U4274 ( .I1(n3083), .I2(n3082), .O(n3419) );
  NAND_GATE U4275 ( .I1(n3084), .I2(n3419), .O(n3414) );
  NAND_GATE U4276 ( .I1(n3421), .I2(n3419), .O(n3085) );
  NAND3_GATE U4277 ( .I1(n3415), .I2(n3414), .I3(n3085), .O(n3408) );
  NAND_GATE U4278 ( .I1(n3100), .I2(n3408), .O(n3404) );
  INV_GATE U4279 ( .I1(n3086), .O(n3087) );
  NAND_GATE U4280 ( .I1(n3087), .I2(n3090), .O(n3099) );
  NAND_GATE U4281 ( .I1(n3089), .I2(n3093), .O(n3097) );
  NAND_GATE U4282 ( .I1(n3091), .I2(n3090), .O(n3092) );
  NAND_GATE U4283 ( .I1(n3093), .I2(n3092), .O(n3094) );
  NAND_GATE U4284 ( .I1(n3095), .I2(n3094), .O(n3096) );
  NAND_GATE U4285 ( .I1(n3097), .I2(n3096), .O(n3098) );
  NAND_GATE U4286 ( .I1(n3099), .I2(n3098), .O(n3407) );
  NAND_GATE U4287 ( .I1(n3100), .I2(n3407), .O(n3403) );
  NAND_GATE U4288 ( .I1(n3408), .I2(n3407), .O(n3101) );
  NAND3_GATE U4289 ( .I1(n3404), .I2(n3403), .I3(n3101), .O(n3397) );
  NAND_GATE U4290 ( .I1(n3116), .I2(n3397), .O(n3391) );
  INV_GATE U4291 ( .I1(n3102), .O(n3103) );
  NAND_GATE U4292 ( .I1(n3103), .I2(n3106), .O(n3115) );
  NAND_GATE U4293 ( .I1(n3105), .I2(n3109), .O(n3113) );
  NAND_GATE U4294 ( .I1(n3107), .I2(n3106), .O(n3108) );
  NAND_GATE U4295 ( .I1(n3109), .I2(n3108), .O(n3110) );
  NAND_GATE U4296 ( .I1(n3111), .I2(n3110), .O(n3112) );
  NAND_GATE U4297 ( .I1(n3113), .I2(n3112), .O(n3114) );
  NAND_GATE U4298 ( .I1(n3115), .I2(n3114), .O(n3395) );
  NAND_GATE U4299 ( .I1(n3116), .I2(n3395), .O(n3390) );
  NAND_GATE U4300 ( .I1(n3397), .I2(n3395), .O(n3117) );
  NAND3_GATE U4301 ( .I1(n3391), .I2(n3390), .I3(n3117), .O(n3384) );
  NAND_GATE U4302 ( .I1(n3132), .I2(n3384), .O(n3380) );
  INV_GATE U4303 ( .I1(n3118), .O(n3119) );
  NAND_GATE U4304 ( .I1(n3119), .I2(n3122), .O(n3131) );
  NAND_GATE U4305 ( .I1(n3121), .I2(n3125), .O(n3129) );
  NAND_GATE U4306 ( .I1(n3123), .I2(n3122), .O(n3124) );
  NAND_GATE U4307 ( .I1(n3125), .I2(n3124), .O(n3126) );
  NAND_GATE U4308 ( .I1(n3127), .I2(n3126), .O(n3128) );
  NAND_GATE U4309 ( .I1(n3129), .I2(n3128), .O(n3130) );
  NAND_GATE U4310 ( .I1(n3131), .I2(n3130), .O(n3383) );
  NAND_GATE U4311 ( .I1(n3132), .I2(n3383), .O(n3379) );
  NAND_GATE U4312 ( .I1(n3384), .I2(n3383), .O(n3133) );
  NAND3_GATE U4313 ( .I1(n3380), .I2(n3379), .I3(n3133), .O(n3373) );
  NAND_GATE U4314 ( .I1(n3148), .I2(n3373), .O(n3369) );
  INV_GATE U4315 ( .I1(n3134), .O(n3135) );
  NAND_GATE U4316 ( .I1(n3135), .I2(n3138), .O(n3147) );
  NAND_GATE U4317 ( .I1(n3137), .I2(n3141), .O(n3145) );
  NAND_GATE U4318 ( .I1(n3139), .I2(n3138), .O(n3140) );
  NAND_GATE U4319 ( .I1(n3141), .I2(n3140), .O(n3142) );
  NAND_GATE U4320 ( .I1(n3143), .I2(n3142), .O(n3144) );
  NAND_GATE U4321 ( .I1(n3145), .I2(n3144), .O(n3146) );
  NAND_GATE U4322 ( .I1(n3147), .I2(n3146), .O(n3372) );
  NAND_GATE U4323 ( .I1(n3148), .I2(n3372), .O(n3368) );
  NAND_GATE U4324 ( .I1(n3373), .I2(n3372), .O(n3149) );
  NAND3_GATE U4325 ( .I1(n3369), .I2(n3368), .I3(n3149), .O(n3362) );
  NAND_GATE U4326 ( .I1(n3164), .I2(n3362), .O(n3358) );
  INV_GATE U4327 ( .I1(n3150), .O(n3151) );
  NAND_GATE U4328 ( .I1(n3151), .I2(n3154), .O(n3163) );
  NAND_GATE U4329 ( .I1(n3153), .I2(n3157), .O(n3161) );
  NAND_GATE U4330 ( .I1(n3155), .I2(n3154), .O(n3156) );
  NAND_GATE U4331 ( .I1(n3157), .I2(n3156), .O(n3158) );
  NAND_GATE U4332 ( .I1(n3159), .I2(n3158), .O(n3160) );
  NAND_GATE U4333 ( .I1(n3161), .I2(n3160), .O(n3162) );
  NAND_GATE U4334 ( .I1(n3163), .I2(n3162), .O(n3361) );
  NAND_GATE U4335 ( .I1(n3164), .I2(n3361), .O(n3357) );
  NAND_GATE U4336 ( .I1(n3362), .I2(n3361), .O(n3165) );
  NAND3_GATE U4337 ( .I1(n3358), .I2(n3357), .I3(n3165), .O(n3351) );
  NAND_GATE U4338 ( .I1(n3180), .I2(n3351), .O(n3347) );
  INV_GATE U4339 ( .I1(n3166), .O(n3167) );
  NAND_GATE U4340 ( .I1(n3167), .I2(n3170), .O(n3179) );
  NAND_GATE U4341 ( .I1(n3169), .I2(n3173), .O(n3177) );
  NAND_GATE U4342 ( .I1(n3171), .I2(n3170), .O(n3172) );
  NAND_GATE U4343 ( .I1(n3173), .I2(n3172), .O(n3174) );
  NAND_GATE U4344 ( .I1(n3175), .I2(n3174), .O(n3176) );
  NAND_GATE U4345 ( .I1(n3177), .I2(n3176), .O(n3178) );
  NAND_GATE U4346 ( .I1(n3179), .I2(n3178), .O(n3350) );
  NAND_GATE U4347 ( .I1(n3180), .I2(n3350), .O(n3346) );
  NAND_GATE U4348 ( .I1(n3351), .I2(n3350), .O(n3181) );
  NAND3_GATE U4349 ( .I1(n3347), .I2(n3346), .I3(n3181), .O(n3340) );
  NAND_GATE U4350 ( .I1(n3196), .I2(n3340), .O(n3336) );
  INV_GATE U4351 ( .I1(n3182), .O(n3183) );
  NAND_GATE U4352 ( .I1(n3183), .I2(n3186), .O(n3195) );
  NAND_GATE U4353 ( .I1(n3185), .I2(n3189), .O(n3193) );
  NAND_GATE U4354 ( .I1(n3187), .I2(n3186), .O(n3188) );
  NAND_GATE U4355 ( .I1(n3189), .I2(n3188), .O(n3190) );
  NAND_GATE U4356 ( .I1(n3191), .I2(n3190), .O(n3192) );
  NAND_GATE U4357 ( .I1(n3193), .I2(n3192), .O(n3194) );
  NAND_GATE U4358 ( .I1(n3195), .I2(n3194), .O(n3339) );
  NAND_GATE U4359 ( .I1(n3196), .I2(n3339), .O(n3335) );
  NAND_GATE U4360 ( .I1(n3340), .I2(n3339), .O(n3197) );
  NAND3_GATE U4361 ( .I1(n3336), .I2(n3335), .I3(n3197), .O(n3665) );
  NAND_GATE U4362 ( .I1(n3212), .I2(n3665), .O(n3659) );
  INV_GATE U4363 ( .I1(n3198), .O(n3199) );
  NAND_GATE U4364 ( .I1(n3199), .I2(n3202), .O(n3211) );
  NAND_GATE U4365 ( .I1(n3201), .I2(n3205), .O(n3209) );
  NAND_GATE U4366 ( .I1(n3203), .I2(n3202), .O(n3204) );
  NAND_GATE U4367 ( .I1(n3205), .I2(n3204), .O(n3206) );
  NAND_GATE U4368 ( .I1(n3207), .I2(n3206), .O(n3208) );
  NAND_GATE U4369 ( .I1(n3209), .I2(n3208), .O(n3210) );
  NAND_GATE U4370 ( .I1(n3211), .I2(n3210), .O(n3663) );
  NAND_GATE U4371 ( .I1(n3212), .I2(n3663), .O(n3658) );
  NAND_GATE U4372 ( .I1(n3665), .I2(n3663), .O(n3213) );
  NAND3_GATE U4373 ( .I1(n3659), .I2(n3658), .I3(n3213), .O(n3329) );
  NAND_GATE U4374 ( .I1(n3228), .I2(n3329), .O(n3325) );
  INV_GATE U4375 ( .I1(n3214), .O(n3215) );
  NAND_GATE U4376 ( .I1(n3215), .I2(n3218), .O(n3227) );
  NAND_GATE U4377 ( .I1(n3217), .I2(n3221), .O(n3225) );
  NAND_GATE U4378 ( .I1(n3219), .I2(n3218), .O(n3220) );
  NAND_GATE U4379 ( .I1(n3221), .I2(n3220), .O(n3222) );
  NAND_GATE U4380 ( .I1(n3223), .I2(n3222), .O(n3224) );
  NAND_GATE U4381 ( .I1(n3225), .I2(n3224), .O(n3226) );
  NAND_GATE U4382 ( .I1(n3227), .I2(n3226), .O(n3328) );
  NAND_GATE U4383 ( .I1(n3228), .I2(n3328), .O(n3324) );
  NAND_GATE U4384 ( .I1(n3329), .I2(n3328), .O(n3229) );
  NAND3_GATE U4385 ( .I1(n3325), .I2(n3324), .I3(n3229), .O(n3317) );
  NAND_GATE U4386 ( .I1(n3230), .I2(n3317), .O(n3311) );
  NAND_GATE U4387 ( .I1(n3316), .I2(n3317), .O(n3231) );
  NAND3_GATE U4388 ( .I1(n3312), .I2(n3311), .I3(n3231), .O(n3305) );
  NAND_GATE U4389 ( .I1(n3246), .I2(n3305), .O(n3301) );
  INV_GATE U4390 ( .I1(n3232), .O(n3233) );
  NAND_GATE U4391 ( .I1(n3233), .I2(n3236), .O(n3245) );
  NAND_GATE U4392 ( .I1(n3235), .I2(n3239), .O(n3243) );
  NAND_GATE U4393 ( .I1(n3237), .I2(n3236), .O(n3238) );
  NAND_GATE U4394 ( .I1(n3239), .I2(n3238), .O(n3240) );
  NAND_GATE U4395 ( .I1(n3241), .I2(n3240), .O(n3242) );
  NAND_GATE U4396 ( .I1(n3243), .I2(n3242), .O(n3244) );
  NAND_GATE U4397 ( .I1(n3245), .I2(n3244), .O(n3304) );
  NAND_GATE U4398 ( .I1(n3246), .I2(n3304), .O(n3300) );
  NAND_GATE U4399 ( .I1(n3305), .I2(n3304), .O(n3247) );
  NAND3_GATE U4400 ( .I1(n3301), .I2(n3300), .I3(n3247), .O(n3294) );
  NAND_GATE U4401 ( .I1(n3262), .I2(n3294), .O(n3288) );
  OR_GATE U4402 ( .I1(n3249), .I2(n3248), .O(n3261) );
  NAND_GATE U4403 ( .I1(n3250), .I2(n3249), .O(n3255) );
  NAND_GATE U4404 ( .I1(n3251), .I2(n3255), .O(n3259) );
  NAND_GATE U4405 ( .I1(n3253), .I2(n3252), .O(n3254) );
  NAND_GATE U4406 ( .I1(n3255), .I2(n3254), .O(n3256) );
  NAND_GATE U4407 ( .I1(n3257), .I2(n3256), .O(n3258) );
  NAND_GATE U4408 ( .I1(n3259), .I2(n3258), .O(n3260) );
  NAND_GATE U4409 ( .I1(n3261), .I2(n3260), .O(n3292) );
  NAND_GATE U4410 ( .I1(n3262), .I2(n3292), .O(n3287) );
  NAND_GATE U4411 ( .I1(n3294), .I2(n3292), .O(n3263) );
  NAND3_GATE U4412 ( .I1(n3288), .I2(n3287), .I3(n3263), .O(n3281) );
  NAND_GATE U4413 ( .I1(n3281), .I2(n3280), .O(n3265) );
  NAND_GATE U4414 ( .I1(n3264), .I2(n3281), .O(n3277) );
  AND3_GATE U4415 ( .I1(n3276), .I2(n3265), .I3(n3277), .O(n3272) );
  NAND_GATE U4416 ( .I1(n1438), .I2(A[31]), .O(n3271) );
  NAND_GATE U4417 ( .I1(n3272), .I2(n3271), .O(n3266) );
  NAND_GATE U4418 ( .I1(n3270), .I2(n3266), .O(n3275) );
  NAND_GATE U4419 ( .I1(n14787), .I2(n3275), .O(n3269) );
  INV_GATE U4420 ( .I1(n3275), .O(n14786) );
  NAND_GATE U4421 ( .I1(n3267), .I2(n14786), .O(n3268) );
  NAND_GATE U4422 ( .I1(n3269), .I2(n3268), .O(\A1[56] ) );
  INV_GATE U4423 ( .I1(n3270), .O(n3273) );
  NAND3_GATE U4424 ( .I1(n3273), .I2(n3272), .I3(n3271), .O(n3274) );
  NAND_GATE U4425 ( .I1(n3275), .I2(n3274), .O(n3682) );
  INV_GATE U4426 ( .I1(n3682), .O(n14789) );
  OR_GATE U4427 ( .I1(n3276), .I2(n3281), .O(n3279) );
  OR_GATE U4428 ( .I1(n3280), .I2(n3277), .O(n3278) );
  AND_GATE U4429 ( .I1(n3279), .I2(n3278), .O(n3286) );
  NAND_GATE U4430 ( .I1(n1203), .I2(n3280), .O(n3284) );
  NAND3_GATE U4431 ( .I1(n3284), .I2(n3283), .I3(n3282), .O(n3285) );
  NAND_GATE U4432 ( .I1(n3286), .I2(n3285), .O(n3685) );
  OR_GATE U4433 ( .I1(n3287), .I2(n3294), .O(n3290) );
  OR_GATE U4434 ( .I1(n3292), .I2(n3288), .O(n3289) );
  AND_GATE U4435 ( .I1(n3290), .I2(n3289), .O(n3299) );
  INV_GATE U4436 ( .I1(n3294), .O(n3291) );
  NAND_GATE U4437 ( .I1(n3291), .I2(n3292), .O(n3297) );
  INV_GATE U4438 ( .I1(n3292), .O(n3293) );
  NAND_GATE U4439 ( .I1(n3294), .I2(n3293), .O(n3296) );
  NAND3_GATE U4440 ( .I1(n3297), .I2(n3296), .I3(n3295), .O(n3298) );
  NAND_GATE U4441 ( .I1(n3299), .I2(n3298), .O(n3690) );
  INV_GATE U4442 ( .I1(n3690), .O(n3693) );
  NAND_GATE U4443 ( .I1(B[25]), .I2(A[30]), .O(n3697) );
  INV_GATE U4444 ( .I1(n3697), .O(n3691) );
  NAND_GATE U4445 ( .I1(n3693), .I2(n3691), .O(n3688) );
  OR_GATE U4446 ( .I1(n3300), .I2(n3305), .O(n3303) );
  OR_GATE U4447 ( .I1(n3304), .I2(n3301), .O(n3302) );
  AND_GATE U4448 ( .I1(n3303), .I2(n3302), .O(n3310) );
  NAND_GATE U4449 ( .I1(n1200), .I2(n3304), .O(n3308) );
  NAND3_GATE U4450 ( .I1(n3308), .I2(n3307), .I3(n3306), .O(n3309) );
  NAND_GATE U4451 ( .I1(n3310), .I2(n3309), .O(n3704) );
  INV_GATE U4452 ( .I1(n3704), .O(n3707) );
  NAND_GATE U4453 ( .I1(B[25]), .I2(A[29]), .O(n3711) );
  INV_GATE U4454 ( .I1(n3711), .O(n3705) );
  NAND_GATE U4455 ( .I1(n3707), .I2(n3705), .O(n3702) );
  OR_GATE U4456 ( .I1(n3311), .I2(n3316), .O(n3314) );
  OR_GATE U4457 ( .I1(n3317), .I2(n3312), .O(n3313) );
  AND_GATE U4458 ( .I1(n3314), .I2(n3313), .O(n3323) );
  INV_GATE U4459 ( .I1(n3317), .O(n3315) );
  NAND_GATE U4460 ( .I1(n3316), .I2(n3315), .O(n3321) );
  INV_GATE U4461 ( .I1(n3316), .O(n3318) );
  NAND_GATE U4462 ( .I1(n3318), .I2(n3317), .O(n3320) );
  NAND3_GATE U4463 ( .I1(n3321), .I2(n3320), .I3(n3319), .O(n3322) );
  NAND_GATE U4464 ( .I1(n3323), .I2(n3322), .O(n4104) );
  INV_GATE U4465 ( .I1(n4104), .O(n4107) );
  NAND_GATE U4466 ( .I1(B[25]), .I2(A[28]), .O(n4111) );
  INV_GATE U4467 ( .I1(n4111), .O(n4105) );
  NAND_GATE U4468 ( .I1(n4107), .I2(n4105), .O(n4102) );
  OR_GATE U4469 ( .I1(n3324), .I2(n3329), .O(n3327) );
  OR_GATE U4470 ( .I1(n3328), .I2(n3325), .O(n3326) );
  AND_GATE U4471 ( .I1(n3327), .I2(n3326), .O(n3334) );
  NAND_GATE U4472 ( .I1(n1192), .I2(n3328), .O(n3332) );
  NAND3_GATE U4473 ( .I1(n3332), .I2(n3331), .I3(n3330), .O(n3333) );
  NAND_GATE U4474 ( .I1(n3334), .I2(n3333), .O(n4088) );
  INV_GATE U4475 ( .I1(n4088), .O(n4091) );
  NAND_GATE U4476 ( .I1(B[25]), .I2(A[27]), .O(n4095) );
  INV_GATE U4477 ( .I1(n4095), .O(n4089) );
  NAND_GATE U4478 ( .I1(n4091), .I2(n4089), .O(n4086) );
  NAND_GATE U4479 ( .I1(B[25]), .I2(A[26]), .O(n4079) );
  INV_GATE U4480 ( .I1(n4079), .O(n4073) );
  OR_GATE U4481 ( .I1(n3335), .I2(n3340), .O(n3338) );
  OR_GATE U4482 ( .I1(n3339), .I2(n3336), .O(n3337) );
  AND_GATE U4483 ( .I1(n3338), .I2(n3337), .O(n3345) );
  NAND_GATE U4484 ( .I1(n1177), .I2(n3339), .O(n3343) );
  NAND3_GATE U4485 ( .I1(n3343), .I2(n3342), .I3(n3341), .O(n3344) );
  NAND_GATE U4486 ( .I1(n3345), .I2(n3344), .O(n4056) );
  INV_GATE U4487 ( .I1(n4056), .O(n4059) );
  NAND_GATE U4488 ( .I1(B[25]), .I2(A[25]), .O(n4063) );
  INV_GATE U4489 ( .I1(n4063), .O(n4057) );
  NAND_GATE U4490 ( .I1(n4059), .I2(n4057), .O(n4054) );
  OR_GATE U4491 ( .I1(n3346), .I2(n3351), .O(n3349) );
  OR_GATE U4492 ( .I1(n3350), .I2(n3347), .O(n3348) );
  AND_GATE U4493 ( .I1(n3349), .I2(n3348), .O(n3356) );
  NAND_GATE U4494 ( .I1(n1175), .I2(n3350), .O(n3354) );
  NAND3_GATE U4495 ( .I1(n3354), .I2(n3353), .I3(n3352), .O(n3355) );
  NAND_GATE U4496 ( .I1(n3356), .I2(n3355), .O(n3722) );
  INV_GATE U4497 ( .I1(n3722), .O(n3720) );
  NAND_GATE U4498 ( .I1(B[25]), .I2(A[24]), .O(n3718) );
  INV_GATE U4499 ( .I1(n3718), .O(n3724) );
  NAND_GATE U4500 ( .I1(n3720), .I2(n3724), .O(n3716) );
  OR_GATE U4501 ( .I1(n3357), .I2(n3362), .O(n3360) );
  OR_GATE U4502 ( .I1(n3361), .I2(n3358), .O(n3359) );
  AND_GATE U4503 ( .I1(n3360), .I2(n3359), .O(n3367) );
  NAND_GATE U4504 ( .I1(n1167), .I2(n3361), .O(n3365) );
  NAND3_GATE U4505 ( .I1(n3365), .I2(n3364), .I3(n3363), .O(n3366) );
  NAND_GATE U4506 ( .I1(n3367), .I2(n3366), .O(n4038) );
  INV_GATE U4507 ( .I1(n4038), .O(n4041) );
  NAND_GATE U4508 ( .I1(B[25]), .I2(A[23]), .O(n4045) );
  INV_GATE U4509 ( .I1(n4045), .O(n4039) );
  NAND_GATE U4510 ( .I1(n4041), .I2(n4039), .O(n4036) );
  OR_GATE U4511 ( .I1(n3368), .I2(n3373), .O(n3371) );
  OR_GATE U4512 ( .I1(n3372), .I2(n3369), .O(n3370) );
  AND_GATE U4513 ( .I1(n3371), .I2(n3370), .O(n3378) );
  NAND_GATE U4514 ( .I1(n1165), .I2(n3372), .O(n3376) );
  NAND3_GATE U4515 ( .I1(n3376), .I2(n3375), .I3(n3374), .O(n3377) );
  NAND_GATE U4516 ( .I1(n3378), .I2(n3377), .O(n4022) );
  INV_GATE U4517 ( .I1(n4022), .O(n4025) );
  NAND_GATE U4518 ( .I1(B[25]), .I2(A[22]), .O(n4029) );
  INV_GATE U4519 ( .I1(n4029), .O(n4023) );
  NAND_GATE U4520 ( .I1(n4025), .I2(n4023), .O(n4020) );
  OR_GATE U4521 ( .I1(n3379), .I2(n3384), .O(n3382) );
  OR_GATE U4522 ( .I1(n3383), .I2(n3380), .O(n3381) );
  AND_GATE U4523 ( .I1(n3382), .I2(n3381), .O(n3389) );
  NAND_GATE U4524 ( .I1(n1129), .I2(n3383), .O(n3387) );
  NAND3_GATE U4525 ( .I1(n3387), .I2(n3386), .I3(n3385), .O(n3388) );
  NAND_GATE U4526 ( .I1(n3389), .I2(n3388), .O(n4006) );
  INV_GATE U4527 ( .I1(n4006), .O(n4009) );
  NAND_GATE U4528 ( .I1(B[25]), .I2(A[21]), .O(n4013) );
  INV_GATE U4529 ( .I1(n4013), .O(n4007) );
  NAND_GATE U4530 ( .I1(n4009), .I2(n4007), .O(n4004) );
  OR_GATE U4531 ( .I1(n3390), .I2(n3397), .O(n3393) );
  OR_GATE U4532 ( .I1(n3395), .I2(n3391), .O(n3392) );
  AND_GATE U4533 ( .I1(n3393), .I2(n3392), .O(n3402) );
  INV_GATE U4534 ( .I1(n3397), .O(n3394) );
  NAND_GATE U4535 ( .I1(n3394), .I2(n3395), .O(n3400) );
  INV_GATE U4536 ( .I1(n3395), .O(n3396) );
  NAND_GATE U4537 ( .I1(n3397), .I2(n3396), .O(n3399) );
  NAND3_GATE U4538 ( .I1(n3400), .I2(n3399), .I3(n3398), .O(n3401) );
  NAND_GATE U4539 ( .I1(n3402), .I2(n3401), .O(n3990) );
  INV_GATE U4540 ( .I1(n3990), .O(n3993) );
  NAND_GATE U4541 ( .I1(B[25]), .I2(A[20]), .O(n3997) );
  INV_GATE U4542 ( .I1(n3997), .O(n3991) );
  NAND_GATE U4543 ( .I1(n3993), .I2(n3991), .O(n3988) );
  OR_GATE U4544 ( .I1(n3403), .I2(n3408), .O(n3406) );
  OR_GATE U4545 ( .I1(n3407), .I2(n3404), .O(n3405) );
  AND_GATE U4546 ( .I1(n3406), .I2(n3405), .O(n3413) );
  NAND_GATE U4547 ( .I1(n1127), .I2(n3407), .O(n3411) );
  NAND3_GATE U4548 ( .I1(n3411), .I2(n3410), .I3(n3409), .O(n3412) );
  NAND_GATE U4549 ( .I1(n3413), .I2(n3412), .O(n3974) );
  INV_GATE U4550 ( .I1(n3974), .O(n3977) );
  NAND_GATE U4551 ( .I1(B[25]), .I2(A[19]), .O(n3981) );
  INV_GATE U4552 ( .I1(n3981), .O(n3975) );
  NAND_GATE U4553 ( .I1(n3977), .I2(n3975), .O(n3972) );
  OR_GATE U4554 ( .I1(n3414), .I2(n3421), .O(n3417) );
  OR_GATE U4555 ( .I1(n3419), .I2(n3415), .O(n3416) );
  AND_GATE U4556 ( .I1(n3417), .I2(n3416), .O(n3426) );
  INV_GATE U4557 ( .I1(n3421), .O(n3418) );
  NAND_GATE U4558 ( .I1(n3418), .I2(n3419), .O(n3424) );
  INV_GATE U4559 ( .I1(n3419), .O(n3420) );
  NAND_GATE U4560 ( .I1(n3421), .I2(n3420), .O(n3423) );
  NAND3_GATE U4561 ( .I1(n3424), .I2(n3423), .I3(n3422), .O(n3425) );
  NAND_GATE U4562 ( .I1(n3426), .I2(n3425), .O(n3958) );
  INV_GATE U4563 ( .I1(n3958), .O(n3961) );
  NAND_GATE U4564 ( .I1(B[25]), .I2(A[18]), .O(n3965) );
  INV_GATE U4565 ( .I1(n3965), .O(n3959) );
  NAND_GATE U4566 ( .I1(n3961), .I2(n3959), .O(n3956) );
  OR_GATE U4567 ( .I1(n3427), .I2(n3432), .O(n3430) );
  OR_GATE U4568 ( .I1(n3431), .I2(n3428), .O(n3429) );
  NAND_GATE U4569 ( .I1(n1151), .I2(n3431), .O(n3435) );
  NAND3_GATE U4570 ( .I1(n3435), .I2(n3434), .I3(n3433), .O(n3436) );
  NAND_GATE U4571 ( .I1(B[25]), .I2(A[17]), .O(n3949) );
  INV_GATE U4572 ( .I1(n3949), .O(n3944) );
  NAND_GATE U4573 ( .I1(n822), .I2(n3944), .O(n3941) );
  OR_GATE U4574 ( .I1(n3437), .I2(n3444), .O(n3440) );
  OR_GATE U4575 ( .I1(n3442), .I2(n3438), .O(n3439) );
  AND_GATE U4576 ( .I1(n3440), .I2(n3439), .O(n3449) );
  INV_GATE U4577 ( .I1(n3444), .O(n3441) );
  NAND_GATE U4578 ( .I1(n3441), .I2(n3442), .O(n3447) );
  INV_GATE U4579 ( .I1(n3442), .O(n3443) );
  NAND_GATE U4580 ( .I1(n3444), .I2(n3443), .O(n3446) );
  NAND3_GATE U4581 ( .I1(n3447), .I2(n3446), .I3(n3445), .O(n3448) );
  NAND_GATE U4582 ( .I1(n3449), .I2(n3448), .O(n3927) );
  INV_GATE U4583 ( .I1(n3927), .O(n3930) );
  NAND_GATE U4584 ( .I1(B[25]), .I2(A[16]), .O(n3934) );
  INV_GATE U4585 ( .I1(n3934), .O(n3928) );
  NAND_GATE U4586 ( .I1(n3930), .I2(n3928), .O(n3925) );
  OR_GATE U4587 ( .I1(n3450), .I2(n3455), .O(n3453) );
  OR_GATE U4588 ( .I1(n3454), .I2(n3451), .O(n3452) );
  AND_GATE U4589 ( .I1(n3453), .I2(n3452), .O(n3460) );
  NAND_GATE U4590 ( .I1(n321), .I2(n3454), .O(n3458) );
  NAND3_GATE U4591 ( .I1(n3458), .I2(n3457), .I3(n3456), .O(n3459) );
  NAND_GATE U4592 ( .I1(n3460), .I2(n3459), .O(n3911) );
  INV_GATE U4593 ( .I1(n3911), .O(n3914) );
  NAND_GATE U4594 ( .I1(B[25]), .I2(A[15]), .O(n3918) );
  INV_GATE U4595 ( .I1(n3918), .O(n3912) );
  NAND_GATE U4596 ( .I1(n3914), .I2(n3912), .O(n3909) );
  OR_GATE U4597 ( .I1(n3461), .I2(n3466), .O(n3464) );
  OR_GATE U4598 ( .I1(n3465), .I2(n3462), .O(n3463) );
  AND_GATE U4599 ( .I1(n3464), .I2(n3463), .O(n3471) );
  NAND_GATE U4600 ( .I1(n1125), .I2(n3465), .O(n3469) );
  NAND3_GATE U4601 ( .I1(n3469), .I2(n3468), .I3(n3467), .O(n3470) );
  NAND_GATE U4602 ( .I1(n3471), .I2(n3470), .O(n3898) );
  NAND_GATE U4603 ( .I1(B[25]), .I2(A[14]), .O(n3902) );
  INV_GATE U4604 ( .I1(n3902), .O(n3896) );
  NAND_GATE U4605 ( .I1(n837), .I2(n3896), .O(n3894) );
  OR_GATE U4606 ( .I1(n3472), .I2(n3477), .O(n3475) );
  OR_GATE U4607 ( .I1(n3476), .I2(n3473), .O(n3474) );
  NAND_GATE U4608 ( .I1(n370), .I2(n3476), .O(n3480) );
  NAND3_GATE U4609 ( .I1(n3480), .I2(n3479), .I3(n3478), .O(n3481) );
  NAND_GATE U4610 ( .I1(B[25]), .I2(A[13]), .O(n3887) );
  INV_GATE U4611 ( .I1(n3887), .O(n3883) );
  NAND_GATE U4612 ( .I1(n934), .I2(n3883), .O(n3880) );
  NAND_GATE U4613 ( .I1(B[25]), .I2(A[12]), .O(n3867) );
  INV_GATE U4614 ( .I1(n3867), .O(n3870) );
  OR_GATE U4615 ( .I1(n3486), .I2(n3482), .O(n3485) );
  OR_GATE U4616 ( .I1(n3483), .I2(n3487), .O(n3484) );
  AND_GATE U4617 ( .I1(n3485), .I2(n3484), .O(n3492) );
  NAND_GATE U4618 ( .I1(n322), .I2(n3486), .O(n3490) );
  NAND3_GATE U4619 ( .I1(n3490), .I2(n3489), .I3(n3488), .O(n3491) );
  NAND_GATE U4620 ( .I1(n3492), .I2(n3491), .O(n3868) );
  NAND_GATE U4621 ( .I1(n3870), .I2(n902), .O(n3873) );
  NAND_GATE U4622 ( .I1(n3498), .I2(n1104), .O(n3495) );
  NAND3_GATE U4623 ( .I1(n3495), .I2(n3494), .I3(n3493), .O(n3502) );
  OR_GATE U4624 ( .I1(n3497), .I2(n3496), .O(n3501) );
  OR_GATE U4625 ( .I1(n3499), .I2(n3498), .O(n3500) );
  NAND3_GATE U4626 ( .I1(n3502), .I2(n3501), .I3(n3500), .O(n3858) );
  INV_GATE U4627 ( .I1(n3858), .O(n3856) );
  NAND_GATE U4628 ( .I1(B[25]), .I2(A[11]), .O(n3857) );
  NAND_GATE U4629 ( .I1(B[25]), .I2(A[10]), .O(n3844) );
  INV_GATE U4630 ( .I1(n3844), .O(n3843) );
  NAND3_GATE U4631 ( .I1(n3506), .I2(n1267), .I3(n3503), .O(n3505) );
  NAND3_GATE U4632 ( .I1(n3507), .I2(n175), .I3(n3503), .O(n3504) );
  AND_GATE U4633 ( .I1(n3505), .I2(n3504), .O(n3512) );
  NAND_GATE U4634 ( .I1(n3506), .I2(n1267), .O(n3510) );
  NAND_GATE U4635 ( .I1(n175), .I2(n3507), .O(n3509) );
  NAND3_GATE U4636 ( .I1(n3510), .I2(n3509), .I3(n3508), .O(n3511) );
  NAND_GATE U4637 ( .I1(n3512), .I2(n3511), .O(n3845) );
  NAND_GATE U4638 ( .I1(n3843), .I2(n1264), .O(n3849) );
  NAND_GATE U4639 ( .I1(n339), .I2(n3520), .O(n3514) );
  NAND3_GATE U4640 ( .I1(n3516), .I2(n3515), .I3(n3514), .O(n3523) );
  NAND4_GATE U4641 ( .I1(n3518), .I2(n3517), .I3(n1210), .I4(n339), .O(n3522)
         );
  OR_GATE U4642 ( .I1(n3520), .I2(n3519), .O(n3521) );
  NAND3_GATE U4643 ( .I1(n3523), .I2(n3522), .I3(n3521), .O(n3731) );
  NAND_GATE U4644 ( .I1(B[25]), .I2(A[8]), .O(n3732) );
  INV_GATE U4645 ( .I1(n3732), .O(n3825) );
  NAND_GATE U4646 ( .I1(n338), .I2(n3825), .O(n3730) );
  INV_GATE U4647 ( .I1(n3524), .O(n3528) );
  NAND3_GATE U4648 ( .I1(n3527), .I2(n3526), .I3(n3525), .O(n3534) );
  NAND4_GATE U4649 ( .I1(n3530), .I2(n3529), .I3(n1213), .I4(n3528), .O(n3533)
         );
  OR_GATE U4650 ( .I1(n3531), .I2(n3598), .O(n3532) );
  NAND3_GATE U4651 ( .I1(n3534), .I2(n3533), .I3(n3532), .O(n3810) );
  NAND_GATE U4652 ( .I1(B[25]), .I2(A[6]), .O(n4350) );
  INV_GATE U4653 ( .I1(n4350), .O(n4348) );
  NAND_GATE U4654 ( .I1(n312), .I2(n4348), .O(n3588) );
  NAND_GATE U4655 ( .I1(B[25]), .I2(A[5]), .O(n3745) );
  INV_GATE U4656 ( .I1(n3745), .O(n3749) );
  NAND_GATE U4657 ( .I1(B[25]), .I2(A[3]), .O(n3784) );
  INV_GATE U4658 ( .I1(n3784), .O(n3777) );
  NAND_GATE U4659 ( .I1(B[25]), .I2(A[2]), .O(n3767) );
  INV_GATE U4660 ( .I1(n3767), .O(n3772) );
  NAND_GATE U4661 ( .I1(n1438), .I2(A[0]), .O(n3535) );
  NAND_GATE U4662 ( .I1(n14241), .I2(n3535), .O(n3536) );
  NAND_GATE U4663 ( .I1(B[27]), .I2(n3536), .O(n3768) );
  NAND_GATE U4664 ( .I1(n1439), .I2(A[1]), .O(n3537) );
  NAND_GATE U4665 ( .I1(n724), .I2(n3537), .O(n3538) );
  NAND_GATE U4666 ( .I1(B[26]), .I2(n3538), .O(n3769) );
  NAND_GATE U4667 ( .I1(n3768), .I2(n3769), .O(n3765) );
  NAND_GATE U4668 ( .I1(n3772), .I2(n3765), .O(n3778) );
  NAND3_GATE U4669 ( .I1(B[25]), .I2(B[26]), .I3(n1254), .O(n3770) );
  INV_GATE U4670 ( .I1(n3770), .O(n3764) );
  INV_GATE U4671 ( .I1(n3765), .O(n3766) );
  NAND_GATE U4672 ( .I1(n3767), .I2(n3766), .O(n3539) );
  NAND_GATE U4673 ( .I1(n3764), .I2(n3539), .O(n3779) );
  NAND_GATE U4674 ( .I1(n3778), .I2(n3779), .O(n3776) );
  NAND_GATE U4675 ( .I1(n3777), .I2(n3776), .O(n3775) );
  NAND3_GATE U4676 ( .I1(n3540), .I2(n3550), .I3(n3542), .O(n3782) );
  NAND_GATE U4677 ( .I1(n3540), .I2(n3542), .O(n3545) );
  NAND_GATE U4678 ( .I1(n3546), .I2(n3541), .O(n3543) );
  OR_GATE U4679 ( .I1(n3543), .I2(n3542), .O(n3544) );
  AND_GATE U4680 ( .I1(n3545), .I2(n3544), .O(n3780) );
  NAND3_GATE U4681 ( .I1(n3548), .I2(n3547), .I3(n3546), .O(n3549) );
  NAND_GATE U4682 ( .I1(n3550), .I2(n3549), .O(n3781) );
  NAND_GATE U4683 ( .I1(n3780), .I2(n3781), .O(n3551) );
  NAND_GATE U4684 ( .I1(n3782), .I2(n3551), .O(n3788) );
  NAND_GATE U4685 ( .I1(n3776), .I2(n3788), .O(n3553) );
  NAND3_GATE U4686 ( .I1(n3777), .I2(n3781), .I3(n3780), .O(n3552) );
  NAND3_GATE U4687 ( .I1(n3775), .I2(n3553), .I3(n3552), .O(n3803) );
  NAND_GATE U4688 ( .I1(B[25]), .I2(A[4]), .O(n4368) );
  NAND_GATE U4689 ( .I1(n3563), .I2(n3564), .O(n3565) );
  OR_GATE U4690 ( .I1(n3565), .I2(n3555), .O(n3561) );
  INV_GATE U4691 ( .I1(n3562), .O(n3566) );
  NAND5_GATE U4692 ( .I1(n3559), .I2(n3558), .I3(n3566), .I4(n3557), .I5(n3556), .O(n3560) );
  AND_GATE U4693 ( .I1(n3561), .I2(n3560), .O(n3798) );
  NAND3_GATE U4694 ( .I1(n3564), .I2(n3563), .I3(n3562), .O(n3568) );
  NAND_GATE U4695 ( .I1(n3566), .I2(n3565), .O(n3567) );
  NAND3_GATE U4696 ( .I1(n3569), .I2(n3568), .I3(n3567), .O(n3799) );
  NAND_GATE U4697 ( .I1(n3798), .I2(n3799), .O(n4360) );
  NAND_GATE U4698 ( .I1(n4368), .I2(n4360), .O(n3570) );
  NAND_GATE U4699 ( .I1(n3803), .I2(n3570), .O(n3572) );
  INV_GATE U4700 ( .I1(n4368), .O(n4362) );
  NAND_GATE U4701 ( .I1(n4362), .I2(n882), .O(n3571) );
  NAND_GATE U4702 ( .I1(n3572), .I2(n3571), .O(n3743) );
  NAND_GATE U4703 ( .I1(n3749), .I2(n3743), .O(n3750) );
  INV_GATE U4704 ( .I1(n3573), .O(n3574) );
  INV_GATE U4705 ( .I1(n3579), .O(n3577) );
  NAND_GATE U4706 ( .I1(n3574), .I2(n3577), .O(n3575) );
  NAND3_GATE U4707 ( .I1(n3580), .I2(n3579), .I3(n304), .O(n3744) );
  NAND3_GATE U4708 ( .I1(n3575), .I2(n3744), .I3(n3580), .O(n3748) );
  NAND3_GATE U4709 ( .I1(n3578), .I2(n3577), .I3(n3576), .O(n3583) );
  NAND3_GATE U4710 ( .I1(n3578), .I2(n3579), .I3(n304), .O(n3581) );
  NAND3_GATE U4711 ( .I1(n3749), .I2(n3748), .I3(n1215), .O(n3585) );
  NAND_GATE U4712 ( .I1(n3580), .I2(n3579), .O(n3582) );
  NAND4_GATE U4713 ( .I1(n3583), .I2(n3582), .I3(n3581), .I4(n2920), .O(n3742)
         );
  NAND_GATE U4714 ( .I1(n3744), .I2(n3742), .O(n3751) );
  NAND_GATE U4715 ( .I1(n3743), .I2(n3751), .O(n3584) );
  NAND_GATE U4716 ( .I1(n3810), .I2(n4350), .O(n3586) );
  NAND_GATE U4717 ( .I1(n3811), .I2(n3586), .O(n3587) );
  NAND_GATE U4718 ( .I1(n3588), .I2(n3587), .O(n3733) );
  INV_GATE U4719 ( .I1(n3594), .O(n3591) );
  NAND3_GATE U4720 ( .I1(n3592), .I2(n3591), .I3(n3590), .O(n3596) );
  AND_GATE U4721 ( .I1(n3596), .I2(n3595), .O(n3736) );
  INV_GATE U4722 ( .I1(n3599), .O(n3600) );
  NAND3_GATE U4723 ( .I1(n3601), .I2(n413), .I3(n3600), .O(n3604) );
  NAND_GATE U4724 ( .I1(n3602), .I2(n413), .O(n3603) );
  NAND3_GATE U4725 ( .I1(n3605), .I2(n3604), .I3(n3603), .O(n3607) );
  NAND_GATE U4726 ( .I1(n3736), .I2(n3607), .O(n3606) );
  NAND_GATE U4727 ( .I1(n3608), .I2(n3606), .O(n3735) );
  NAND_GATE U4728 ( .I1(n3733), .I2(n3735), .O(n3611) );
  INV_GATE U4729 ( .I1(n3607), .O(n3609) );
  NAND_GATE U4730 ( .I1(n3609), .I2(n3608), .O(n3738) );
  NAND_GATE U4731 ( .I1(B[25]), .I2(A[7]), .O(n3818) );
  INV_GATE U4732 ( .I1(n3818), .O(n3737) );
  NAND3_GATE U4733 ( .I1(n3738), .I2(n3736), .I3(n3737), .O(n3610) );
  NAND_GATE U4734 ( .I1(n3737), .I2(n3733), .O(n3734) );
  NAND_GATE U4735 ( .I1(n3730), .I2(n3612), .O(n3835) );
  NAND_GATE U4736 ( .I1(B[25]), .I2(A[9]), .O(n4454) );
  NAND3_GATE U4737 ( .I1(n3617), .I2(n3613), .I3(n906), .O(n3616) );
  OR_GATE U4738 ( .I1(n3617), .I2(n3614), .O(n3615) );
  AND_GATE U4739 ( .I1(n3616), .I2(n3615), .O(n3623) );
  NAND_GATE U4740 ( .I1(n906), .I2(n3617), .O(n3620) );
  NAND_GATE U4741 ( .I1(n3618), .I2(n328), .O(n3619) );
  NAND3_GATE U4742 ( .I1(n3621), .I2(n3620), .I3(n3619), .O(n3622) );
  NAND_GATE U4743 ( .I1(n4454), .I2(n3836), .O(n3624) );
  NAND_GATE U4744 ( .I1(n3835), .I2(n3624), .O(n3626) );
  INV_GATE U4745 ( .I1(n4454), .O(n3831) );
  NAND_GATE U4746 ( .I1(n3831), .I2(n821), .O(n3625) );
  NAND_GATE U4747 ( .I1(n3844), .I2(n3845), .O(n3627) );
  NAND_GATE U4748 ( .I1(n3850), .I2(n3627), .O(n3628) );
  NAND_GATE U4749 ( .I1(n3858), .I2(n3857), .O(n3629) );
  NAND_GATE U4750 ( .I1(n3867), .I2(n3868), .O(n3630) );
  NAND_GATE U4751 ( .I1(n3874), .I2(n3630), .O(n3631) );
  NAND_GATE U4752 ( .I1(n3873), .I2(n3631), .O(n3884) );
  NAND_GATE U4753 ( .I1(n3884), .I2(n3632), .O(n3633) );
  NAND_GATE U4754 ( .I1(n3880), .I2(n3633), .O(n3897) );
  NAND_GATE U4755 ( .I1(n3898), .I2(n3902), .O(n3634) );
  NAND_GATE U4756 ( .I1(n3897), .I2(n3634), .O(n3635) );
  NAND_GATE U4757 ( .I1(n3894), .I2(n3635), .O(n3913) );
  NAND_GATE U4758 ( .I1(n3911), .I2(n3918), .O(n3636) );
  NAND_GATE U4759 ( .I1(n3913), .I2(n3636), .O(n3637) );
  NAND_GATE U4760 ( .I1(n3909), .I2(n3637), .O(n3929) );
  NAND_GATE U4761 ( .I1(n3927), .I2(n3934), .O(n3638) );
  NAND_GATE U4762 ( .I1(n3929), .I2(n3638), .O(n3639) );
  NAND_GATE U4763 ( .I1(n3925), .I2(n3639), .O(n3945) );
  NAND_GATE U4764 ( .I1(n3943), .I2(n3949), .O(n3640) );
  NAND_GATE U4765 ( .I1(n3945), .I2(n3640), .O(n3641) );
  NAND_GATE U4766 ( .I1(n3941), .I2(n3641), .O(n3960) );
  NAND_GATE U4767 ( .I1(n3958), .I2(n3965), .O(n3642) );
  NAND_GATE U4768 ( .I1(n3960), .I2(n3642), .O(n3643) );
  NAND_GATE U4769 ( .I1(n3956), .I2(n3643), .O(n3976) );
  NAND_GATE U4770 ( .I1(n3974), .I2(n3981), .O(n3644) );
  NAND_GATE U4771 ( .I1(n3976), .I2(n3644), .O(n3645) );
  NAND_GATE U4772 ( .I1(n3972), .I2(n3645), .O(n3992) );
  NAND_GATE U4773 ( .I1(n3990), .I2(n3997), .O(n3646) );
  NAND_GATE U4774 ( .I1(n3992), .I2(n3646), .O(n3647) );
  NAND_GATE U4775 ( .I1(n3988), .I2(n3647), .O(n4008) );
  NAND_GATE U4776 ( .I1(n4006), .I2(n4013), .O(n3648) );
  NAND_GATE U4777 ( .I1(n4008), .I2(n3648), .O(n3649) );
  NAND_GATE U4778 ( .I1(n4004), .I2(n3649), .O(n4024) );
  NAND_GATE U4779 ( .I1(n4022), .I2(n4029), .O(n3650) );
  NAND_GATE U4780 ( .I1(n4024), .I2(n3650), .O(n3651) );
  NAND_GATE U4781 ( .I1(n4020), .I2(n3651), .O(n4040) );
  NAND_GATE U4782 ( .I1(n4038), .I2(n4045), .O(n3652) );
  NAND_GATE U4783 ( .I1(n4040), .I2(n3652), .O(n3653) );
  NAND_GATE U4784 ( .I1(n4036), .I2(n3653), .O(n3719) );
  NAND_GATE U4785 ( .I1(n3722), .I2(n3718), .O(n3654) );
  NAND_GATE U4786 ( .I1(n3719), .I2(n3654), .O(n3655) );
  NAND_GATE U4787 ( .I1(n3716), .I2(n3655), .O(n4058) );
  NAND_GATE U4788 ( .I1(n4056), .I2(n4063), .O(n3656) );
  NAND_GATE U4789 ( .I1(n4058), .I2(n3656), .O(n3657) );
  NAND_GATE U4790 ( .I1(n4054), .I2(n3657), .O(n4075) );
  NAND_GATE U4791 ( .I1(n4073), .I2(n4075), .O(n4070) );
  OR_GATE U4792 ( .I1(n3658), .I2(n3665), .O(n3661) );
  OR_GATE U4793 ( .I1(n3663), .I2(n3659), .O(n3660) );
  AND_GATE U4794 ( .I1(n3661), .I2(n3660), .O(n3670) );
  INV_GATE U4795 ( .I1(n3665), .O(n3662) );
  NAND_GATE U4796 ( .I1(n3662), .I2(n3663), .O(n3668) );
  INV_GATE U4797 ( .I1(n3663), .O(n3664) );
  NAND_GATE U4798 ( .I1(n3665), .I2(n3664), .O(n3667) );
  NAND3_GATE U4799 ( .I1(n3668), .I2(n3667), .I3(n3666), .O(n3669) );
  NAND_GATE U4800 ( .I1(n3670), .I2(n3669), .O(n4071) );
  INV_GATE U4801 ( .I1(n4071), .O(n4074) );
  INV_GATE U4802 ( .I1(n4075), .O(n4072) );
  NAND_GATE U4803 ( .I1(n4079), .I2(n4072), .O(n3671) );
  NAND_GATE U4804 ( .I1(n4074), .I2(n3671), .O(n3672) );
  NAND_GATE U4805 ( .I1(n4070), .I2(n3672), .O(n4090) );
  NAND_GATE U4806 ( .I1(n4088), .I2(n4095), .O(n3673) );
  NAND_GATE U4807 ( .I1(n4090), .I2(n3673), .O(n3674) );
  NAND_GATE U4808 ( .I1(n4086), .I2(n3674), .O(n4106) );
  NAND_GATE U4809 ( .I1(n4104), .I2(n4111), .O(n3675) );
  NAND_GATE U4810 ( .I1(n4106), .I2(n3675), .O(n3676) );
  NAND_GATE U4811 ( .I1(n4102), .I2(n3676), .O(n3706) );
  NAND_GATE U4812 ( .I1(n3704), .I2(n3711), .O(n3677) );
  NAND_GATE U4813 ( .I1(n3706), .I2(n3677), .O(n3678) );
  NAND_GATE U4814 ( .I1(n3702), .I2(n3678), .O(n3692) );
  NAND_GATE U4815 ( .I1(n3690), .I2(n3697), .O(n3679) );
  NAND_GATE U4816 ( .I1(n3692), .I2(n3679), .O(n3681) );
  NAND_GATE U4817 ( .I1(n1437), .I2(A[31]), .O(n3680) );
  NAND_GATE U4818 ( .I1(n14789), .I2(n3687), .O(n3684) );
  INV_GATE U4819 ( .I1(n3687), .O(n14788) );
  NAND_GATE U4820 ( .I1(n3682), .I2(n14788), .O(n3683) );
  NAND_GATE U4821 ( .I1(n3684), .I2(n3683), .O(\A1[55] ) );
  NAND_GATE U4822 ( .I1(n3685), .I2(n407), .O(n3686) );
  NAND_GATE U4823 ( .I1(n3687), .I2(n3686), .O(n4121) );
  INV_GATE U4824 ( .I1(n4121), .O(n14791) );
  INV_GATE U4825 ( .I1(n3688), .O(n3689) );
  NAND_GATE U4826 ( .I1(n3689), .I2(n3692), .O(n3701) );
  NAND_GATE U4827 ( .I1(n3691), .I2(n3695), .O(n3699) );
  NAND_GATE U4828 ( .I1(n3693), .I2(n3692), .O(n3694) );
  NAND_GATE U4829 ( .I1(n3695), .I2(n3694), .O(n3696) );
  NAND_GATE U4830 ( .I1(n3697), .I2(n3696), .O(n3698) );
  NAND_GATE U4831 ( .I1(n3699), .I2(n3698), .O(n3700) );
  NAND_GATE U4832 ( .I1(n3701), .I2(n3700), .O(n4124) );
  NAND_GATE U4833 ( .I1(B[24]), .I2(A[30]), .O(n4136) );
  INV_GATE U4834 ( .I1(n4136), .O(n4118) );
  INV_GATE U4835 ( .I1(n3702), .O(n3703) );
  NAND_GATE U4836 ( .I1(n3703), .I2(n3706), .O(n3715) );
  NAND_GATE U4837 ( .I1(n3705), .I2(n3709), .O(n3713) );
  NAND_GATE U4838 ( .I1(n3707), .I2(n3706), .O(n3708) );
  NAND_GATE U4839 ( .I1(n3709), .I2(n3708), .O(n3710) );
  NAND_GATE U4840 ( .I1(n3711), .I2(n3710), .O(n3712) );
  NAND_GATE U4841 ( .I1(n3713), .I2(n3712), .O(n3714) );
  NAND_GATE U4842 ( .I1(n3715), .I2(n3714), .O(n4134) );
  NAND_GATE U4843 ( .I1(n4118), .I2(n4134), .O(n4130) );
  NAND_GATE U4844 ( .I1(B[24]), .I2(A[29]), .O(n4147) );
  INV_GATE U4845 ( .I1(n4147), .O(n4116) );
  NAND_GATE U4846 ( .I1(B[24]), .I2(A[28]), .O(n4158) );
  INV_GATE U4847 ( .I1(n4158), .O(n4100) );
  NAND_GATE U4848 ( .I1(B[24]), .I2(A[27]), .O(n4169) );
  INV_GATE U4849 ( .I1(n4169), .O(n4084) );
  NAND_GATE U4850 ( .I1(B[24]), .I2(A[26]), .O(n4180) );
  INV_GATE U4851 ( .I1(n4180), .O(n4068) );
  NAND_GATE U4852 ( .I1(B[24]), .I2(A[25]), .O(n4191) );
  INV_GATE U4853 ( .I1(n4191), .O(n4052) );
  INV_GATE U4854 ( .I1(n3716), .O(n3717) );
  NAND_GATE U4855 ( .I1(n3717), .I2(n3719), .O(n3729) );
  INV_GATE U4856 ( .I1(n3719), .O(n3721) );
  NAND3_GATE U4857 ( .I1(n3718), .I2(n3721), .I3(n3722), .O(n3727) );
  NAND_GATE U4858 ( .I1(n3720), .I2(n3719), .O(n3726) );
  NAND_GATE U4859 ( .I1(n3722), .I2(n3721), .O(n3723) );
  NAND_GATE U4860 ( .I1(n3724), .I2(n3723), .O(n3725) );
  NAND3_GATE U4861 ( .I1(n3727), .I2(n3726), .I3(n3725), .O(n3728) );
  NAND_GATE U4862 ( .I1(n3729), .I2(n3728), .O(n4189) );
  NAND_GATE U4863 ( .I1(n4052), .I2(n4189), .O(n4186) );
  NAND_GATE U4864 ( .I1(B[24]), .I2(A[24]), .O(n4202) );
  INV_GATE U4865 ( .I1(n4202), .O(n4050) );
  NAND_GATE U4866 ( .I1(B[24]), .I2(A[23]), .O(n4500) );
  INV_GATE U4867 ( .I1(n4500), .O(n4034) );
  NAND_GATE U4868 ( .I1(B[24]), .I2(A[22]), .O(n4213) );
  INV_GATE U4869 ( .I1(n4213), .O(n4018) );
  NAND_GATE U4870 ( .I1(B[24]), .I2(A[21]), .O(n4224) );
  INV_GATE U4871 ( .I1(n4224), .O(n4002) );
  NAND_GATE U4872 ( .I1(B[24]), .I2(A[20]), .O(n4237) );
  INV_GATE U4873 ( .I1(n4237), .O(n3986) );
  NAND_GATE U4874 ( .I1(B[24]), .I2(A[19]), .O(n4248) );
  INV_GATE U4875 ( .I1(n4248), .O(n3970) );
  NAND_GATE U4876 ( .I1(B[24]), .I2(A[18]), .O(n4259) );
  INV_GATE U4877 ( .I1(n4259), .O(n3954) );
  NAND_GATE U4878 ( .I1(B[24]), .I2(A[17]), .O(n4270) );
  INV_GATE U4879 ( .I1(n4270), .O(n3939) );
  NAND_GATE U4880 ( .I1(B[24]), .I2(A[16]), .O(n4281) );
  INV_GATE U4881 ( .I1(n4281), .O(n3923) );
  NAND_GATE U4882 ( .I1(B[24]), .I2(A[15]), .O(n4292) );
  INV_GATE U4883 ( .I1(n4292), .O(n3907) );
  NAND_GATE U4884 ( .I1(B[24]), .I2(A[14]), .O(n4303) );
  INV_GATE U4885 ( .I1(n4303), .O(n3892) );
  NAND_GATE U4886 ( .I1(B[24]), .I2(A[13]), .O(n4310) );
  INV_GATE U4887 ( .I1(n4310), .O(n3878) );
  NAND_GATE U4888 ( .I1(B[24]), .I2(A[12]), .O(n4326) );
  INV_GATE U4889 ( .I1(n4326), .O(n3864) );
  NAND_GATE U4890 ( .I1(B[24]), .I2(A[11]), .O(n4331) );
  INV_GATE U4891 ( .I1(n4331), .O(n3854) );
  NAND_GATE U4892 ( .I1(B[24]), .I2(A[10]), .O(n4464) );
  INV_GATE U4893 ( .I1(n4464), .O(n4449) );
  NAND_GATE U4894 ( .I1(B[24]), .I2(A[9]), .O(n4442) );
  INV_GATE U4895 ( .I1(n4442), .O(n4340) );
  NAND_GATE U4896 ( .I1(n3731), .I2(n731), .O(n3824) );
  NAND3_GATE U4897 ( .I1(n3825), .I2(n3824), .I3(n3830), .O(n4341) );
  NAND3_GATE U4898 ( .I1(n3731), .I2(n3732), .I3(n731), .O(n3828) );
  NAND3_GATE U4899 ( .I1(n4340), .I2(n4341), .I3(n1212), .O(n4457) );
  NAND_GATE U4900 ( .I1(B[24]), .I2(A[8]), .O(n4582) );
  INV_GATE U4901 ( .I1(n4582), .O(n4580) );
  NAND_GATE U4902 ( .I1(n745), .I2(n3735), .O(n3817) );
  AND3_GATE U4903 ( .I1(n3817), .I2(n3818), .I3(n3816), .O(n3741) );
  OR_GATE U4904 ( .I1(n3735), .I2(n3734), .O(n3740) );
  NAND4_GATE U4905 ( .I1(n3738), .I2(n745), .I3(n3737), .I4(n3736), .O(n3739)
         );
  NAND_GATE U4906 ( .I1(n3740), .I2(n3739), .O(n3819) );
  NAND_GATE U4907 ( .I1(n4580), .I2(n1268), .O(n3823) );
  NAND_GATE U4908 ( .I1(B[24]), .I2(A[7]), .O(n4357) );
  INV_GATE U4909 ( .I1(n4357), .O(n4346) );
  NAND_GATE U4910 ( .I1(B[24]), .I2(A[6]), .O(n4609) );
  INV_GATE U4911 ( .I1(n4609), .O(n4422) );
  NAND_GATE U4912 ( .I1(n883), .I2(n3751), .O(n3747) );
  NAND3_GATE U4913 ( .I1(n3744), .I2(n3743), .I3(n3742), .O(n3746) );
  NAND3_GATE U4914 ( .I1(n3747), .I2(n3746), .I3(n3745), .O(n3754) );
  NAND4_GATE U4915 ( .I1(n3749), .I2(n3748), .I3(n883), .I4(n1215), .O(n3753)
         );
  OR_GATE U4916 ( .I1(n3751), .I2(n3750), .O(n3752) );
  NAND3_GATE U4917 ( .I1(n3754), .I2(n3753), .I3(n3752), .O(n4424) );
  NAND_GATE U4918 ( .I1(n4422), .I2(n4426), .O(n3809) );
  NAND_GATE U4919 ( .I1(B[24]), .I2(A[5]), .O(n4417) );
  INV_GATE U4920 ( .I1(n4417), .O(n3806) );
  NAND_GATE U4921 ( .I1(B[24]), .I2(A[4]), .O(n4616) );
  INV_GATE U4922 ( .I1(n4616), .O(n4403) );
  NAND_GATE U4923 ( .I1(B[24]), .I2(A[3]), .O(n4386) );
  INV_GATE U4924 ( .I1(n4386), .O(n4377) );
  NAND_GATE U4925 ( .I1(B[24]), .I2(A[2]), .O(n4665) );
  NAND_GATE U4926 ( .I1(n1438), .I2(A[1]), .O(n3755) );
  NAND_GATE U4927 ( .I1(n724), .I2(n3755), .O(n3756) );
  NAND_GATE U4928 ( .I1(B[25]), .I2(n3756), .O(n3761) );
  NAND_GATE U4929 ( .I1(n4665), .I2(n3761), .O(n3757) );
  NAND_GATE U4930 ( .I1(n414), .I2(n3757), .O(n3763) );
  INV_GATE U4931 ( .I1(n4665), .O(n4663) );
  NAND_GATE U4932 ( .I1(n1437), .I2(A[0]), .O(n3758) );
  NAND_GATE U4933 ( .I1(n14241), .I2(n3758), .O(n3759) );
  NAND_GATE U4934 ( .I1(B[26]), .I2(n3759), .O(n3760) );
  NAND_GATE U4935 ( .I1(n3761), .I2(n3760), .O(n4393) );
  NAND_GATE U4936 ( .I1(n4663), .I2(n4393), .O(n3762) );
  NAND_GATE U4937 ( .I1(n3763), .I2(n3762), .O(n4383) );
  NAND_GATE U4938 ( .I1(n4377), .I2(n4383), .O(n4373) );
  NAND_GATE U4939 ( .I1(n3765), .I2(n3764), .O(n4375) );
  NAND3_GATE U4940 ( .I1(n3767), .I2(n3770), .I3(n3766), .O(n4376) );
  NAND3_GATE U4941 ( .I1(n3770), .I2(n3769), .I3(n3768), .O(n3771) );
  NAND_GATE U4942 ( .I1(n3772), .I2(n3771), .O(n4374) );
  NAND3_GATE U4943 ( .I1(n4375), .I2(n4376), .I3(n4374), .O(n4382) );
  NAND_GATE U4944 ( .I1(n4384), .I2(n4382), .O(n4380) );
  NAND_GATE U4945 ( .I1(n4383), .I2(n4380), .O(n3774) );
  NAND_GATE U4946 ( .I1(n4377), .I2(n4380), .O(n3773) );
  NAND3_GATE U4947 ( .I1(n4373), .I2(n3774), .I3(n3773), .O(n4406) );
  NAND_GATE U4948 ( .I1(n4403), .I2(n4406), .O(n3797) );
  INV_GATE U4949 ( .I1(n3776), .O(n3789) );
  NAND4_GATE U4950 ( .I1(n3777), .I2(n3781), .I3(n3780), .I4(n3789), .O(n3792)
         );
  NAND3_GATE U4951 ( .I1(n3779), .I2(n3778), .I3(n3784), .O(n3787) );
  NAND3_GATE U4952 ( .I1(n3781), .I2(n3780), .I3(n3784), .O(n3786) );
  INV_GATE U4953 ( .I1(n3782), .O(n3783) );
  NAND_GATE U4954 ( .I1(n3784), .I2(n3783), .O(n3785) );
  NAND3_GATE U4955 ( .I1(n3787), .I2(n3786), .I3(n3785), .O(n3791) );
  NAND_GATE U4956 ( .I1(n3789), .I2(n3788), .O(n3790) );
  NAND_GATE U4957 ( .I1(n3791), .I2(n3790), .O(n3793) );
  NAND3_GATE U4958 ( .I1(n3794), .I2(n3792), .I3(n3793), .O(n4404) );
  NAND_GATE U4959 ( .I1(n4403), .I2(n389), .O(n3796) );
  NAND4_GATE U4960 ( .I1(n3794), .I2(n3793), .I3(n4406), .I4(n3792), .O(n3795)
         );
  NAND3_GATE U4961 ( .I1(n3797), .I2(n3796), .I3(n3795), .O(n4372) );
  NAND3_GATE U4962 ( .I1(n3803), .I2(n4362), .I3(n882), .O(n4365) );
  NAND_GATE U4963 ( .I1(n3803), .I2(n4362), .O(n3801) );
  NAND3_GATE U4964 ( .I1(n3799), .I2(n3798), .I3(n4362), .O(n3800) );
  NAND_GATE U4965 ( .I1(n3801), .I2(n3800), .O(n3802) );
  NAND_GATE U4966 ( .I1(n4365), .I2(n3802), .O(n4370) );
  INV_GATE U4967 ( .I1(n3803), .O(n4361) );
  NAND_GATE U4968 ( .I1(n4361), .I2(n4360), .O(n3805) );
  NAND_GATE U4969 ( .I1(n3803), .I2(n882), .O(n3804) );
  NAND_GATE U4970 ( .I1(n3805), .I2(n3804), .O(n4367) );
  NAND_GATE U4971 ( .I1(n4609), .I2(n4424), .O(n3807) );
  NAND_GATE U4972 ( .I1(n4425), .I2(n3807), .O(n3808) );
  NAND_GATE U4973 ( .I1(n3809), .I2(n3808), .O(n4354) );
  NAND_GATE U4974 ( .I1(n4346), .I2(n4354), .O(n4347) );
  NAND3_GATE U4975 ( .I1(n4348), .I2(n3811), .I3(n312), .O(n4352) );
  NAND3_GATE U4976 ( .I1(n3813), .I2(n4352), .I3(n4348), .O(n4345) );
  NAND_GATE U4977 ( .I1(n3810), .I2(n929), .O(n3813) );
  NAND_GATE U4978 ( .I1(n3813), .I2(n3812), .O(n4349) );
  NAND3_GATE U4979 ( .I1(n4346), .I2(n4345), .I3(n4356), .O(n3815) );
  NAND3_GATE U4980 ( .I1(n4354), .I2(n4345), .I3(n4356), .O(n3814) );
  NAND3_GATE U4981 ( .I1(n4347), .I2(n3815), .I3(n3814), .O(n4434) );
  NAND4_GATE U4982 ( .I1(n4582), .I2(n3818), .I3(n3817), .I4(n3816), .O(n3821)
         );
  NAND_GATE U4983 ( .I1(n4582), .I2(n3819), .O(n3820) );
  NAND3_GATE U4984 ( .I1(n4434), .I2(n3821), .I3(n3820), .O(n3822) );
  NAND_GATE U4985 ( .I1(n3823), .I2(n3822), .O(n4338) );
  NAND_GATE U4986 ( .I1(n3825), .I2(n3824), .O(n3826) );
  NAND3_GATE U4987 ( .I1(n3828), .I2(n3827), .I3(n3826), .O(n3829) );
  NAND_GATE U4988 ( .I1(n3830), .I2(n3829), .O(n4339) );
  NAND_GATE U4989 ( .I1(n4338), .I2(n4339), .O(n4461) );
  NAND_GATE U4990 ( .I1(n4340), .I2(n4338), .O(n4458) );
  NAND3_GATE U4991 ( .I1(n4457), .I2(n4461), .I3(n4458), .O(n4456) );
  NAND_GATE U4992 ( .I1(n4449), .I2(n4456), .O(n3841) );
  NAND3_GATE U4993 ( .I1(n821), .I2(n3831), .I3(n3835), .O(n4452) );
  NAND3_GATE U4994 ( .I1(n3836), .I2(n4454), .I3(n702), .O(n3832) );
  NAND_GATE U4995 ( .I1(n3831), .I2(n3837), .O(n3834) );
  NAND3_GATE U4996 ( .I1(n3832), .I2(n3838), .I3(n3834), .O(n4448) );
  NAND_GATE U4997 ( .I1(n4452), .I2(n4448), .O(n3833) );
  NAND_GATE U4998 ( .I1(n4456), .I2(n3833), .O(n3840) );
  NAND_GATE U4999 ( .I1(n3835), .I2(n821), .O(n3838) );
  NAND_GATE U5000 ( .I1(n702), .I2(n3836), .O(n3837) );
  NAND_GATE U5001 ( .I1(n3838), .I2(n3837), .O(n4453) );
  NAND3_GATE U5002 ( .I1(n4449), .I2(n4460), .I3(n3839), .O(n4447) );
  NAND3_GATE U5003 ( .I1(n3841), .I2(n3840), .I3(n4447), .O(n4332) );
  NAND_GATE U5004 ( .I1(n3854), .I2(n4332), .O(n4334) );
  NAND_GATE U5005 ( .I1(n3845), .I2(n1338), .O(n3842) );
  NAND_GATE U5006 ( .I1(n3843), .I2(n3842), .O(n3848) );
  NAND3_GATE U5007 ( .I1(n3845), .I2(n1338), .I3(n3844), .O(n3847) );
  NAND_GATE U5008 ( .I1(n1264), .I2(n3850), .O(n3846) );
  NAND3_GATE U5009 ( .I1(n3848), .I2(n3847), .I3(n3846), .O(n3853) );
  INV_GATE U5010 ( .I1(n3849), .O(n3851) );
  NAND_GATE U5011 ( .I1(n3851), .I2(n3850), .O(n3852) );
  NAND_GATE U5012 ( .I1(n4332), .I2(n811), .O(n3855) );
  NAND3_GATE U5013 ( .I1(n4334), .I2(n4333), .I3(n3855), .O(n4323) );
  NAND_GATE U5014 ( .I1(n3864), .I2(n4323), .O(n4318) );
  NAND_GATE U5015 ( .I1(n3856), .I2(n894), .O(n3860) );
  NAND3_GATE U5016 ( .I1(n3858), .I2(n1324), .I3(n3857), .O(n3859) );
  NAND3_GATE U5017 ( .I1(n3861), .I2(n3860), .I3(n3859), .O(n3863) );
  NAND_GATE U5018 ( .I1(n1255), .I2(n894), .O(n3862) );
  NAND_GATE U5019 ( .I1(n3863), .I2(n3862), .O(n4322) );
  NAND_GATE U5020 ( .I1(n3864), .I2(n4322), .O(n4319) );
  NAND_GATE U5021 ( .I1(n4323), .I2(n4322), .O(n3865) );
  NAND3_GATE U5022 ( .I1(n4318), .I2(n4319), .I3(n3865), .O(n4311) );
  NAND_GATE U5023 ( .I1(n3878), .I2(n4311), .O(n4313) );
  NAND_GATE U5024 ( .I1(n902), .I2(n3874), .O(n3866) );
  NAND_GATE U5025 ( .I1(n3868), .I2(n895), .O(n3869) );
  NAND_GATE U5026 ( .I1(n3870), .I2(n3869), .O(n3871) );
  NAND_GATE U5027 ( .I1(n3872), .I2(n3871), .O(n3877) );
  INV_GATE U5028 ( .I1(n3873), .O(n3875) );
  NAND_GATE U5029 ( .I1(n3875), .I2(n3874), .O(n3876) );
  NAND_GATE U5030 ( .I1(n3877), .I2(n3876), .O(n4314) );
  NAND_GATE U5031 ( .I1(n3878), .I2(n4314), .O(n4312) );
  NAND_GATE U5032 ( .I1(n4311), .I2(n4314), .O(n3879) );
  NAND3_GATE U5033 ( .I1(n4313), .I2(n4312), .I3(n3879), .O(n4302) );
  NAND_GATE U5034 ( .I1(n3892), .I2(n4302), .O(n4298) );
  INV_GATE U5035 ( .I1(n3880), .O(n3881) );
  NAND_GATE U5036 ( .I1(n3881), .I2(n3884), .O(n3891) );
  NAND_GATE U5037 ( .I1(n3883), .I2(n3882), .O(n3889) );
  NAND_GATE U5038 ( .I1(n934), .I2(n3884), .O(n3885) );
  NAND_GATE U5039 ( .I1(n3885), .I2(n3882), .O(n3886) );
  NAND_GATE U5040 ( .I1(n3887), .I2(n3886), .O(n3888) );
  NAND_GATE U5041 ( .I1(n3889), .I2(n3888), .O(n3890) );
  NAND_GATE U5042 ( .I1(n3891), .I2(n3890), .O(n4301) );
  NAND_GATE U5043 ( .I1(n4302), .I2(n4301), .O(n3893) );
  NAND3_GATE U5044 ( .I1(n4298), .I2(n4297), .I3(n3893), .O(n4291) );
  NAND_GATE U5045 ( .I1(n3907), .I2(n4291), .O(n4287) );
  INV_GATE U5046 ( .I1(n3894), .O(n3895) );
  NAND_GATE U5047 ( .I1(n3895), .I2(n3897), .O(n3906) );
  NAND_GATE U5048 ( .I1(n3896), .I2(n3899), .O(n3904) );
  NAND_GATE U5049 ( .I1(n837), .I2(n3897), .O(n3900) );
  NAND_GATE U5050 ( .I1(n3898), .I2(n1332), .O(n3899) );
  NAND_GATE U5051 ( .I1(n3900), .I2(n3899), .O(n3901) );
  NAND_GATE U5052 ( .I1(n3902), .I2(n3901), .O(n3903) );
  NAND_GATE U5053 ( .I1(n3904), .I2(n3903), .O(n3905) );
  NAND_GATE U5054 ( .I1(n3906), .I2(n3905), .O(n4290) );
  NAND_GATE U5055 ( .I1(n4291), .I2(n4290), .O(n3908) );
  NAND3_GATE U5056 ( .I1(n4287), .I2(n4286), .I3(n3908), .O(n4280) );
  NAND_GATE U5057 ( .I1(n3923), .I2(n4280), .O(n4276) );
  INV_GATE U5058 ( .I1(n3909), .O(n3910) );
  NAND_GATE U5059 ( .I1(n3910), .I2(n3913), .O(n3922) );
  NAND_GATE U5060 ( .I1(n3912), .I2(n3916), .O(n3920) );
  NAND_GATE U5061 ( .I1(n3914), .I2(n3913), .O(n3915) );
  NAND_GATE U5062 ( .I1(n3916), .I2(n3915), .O(n3917) );
  NAND_GATE U5063 ( .I1(n3918), .I2(n3917), .O(n3919) );
  NAND_GATE U5064 ( .I1(n3920), .I2(n3919), .O(n3921) );
  NAND_GATE U5065 ( .I1(n3922), .I2(n3921), .O(n4279) );
  NAND_GATE U5066 ( .I1(n4280), .I2(n4279), .O(n3924) );
  NAND3_GATE U5067 ( .I1(n4276), .I2(n4275), .I3(n3924), .O(n4269) );
  NAND_GATE U5068 ( .I1(n3939), .I2(n4269), .O(n4265) );
  INV_GATE U5069 ( .I1(n3925), .O(n3926) );
  NAND_GATE U5070 ( .I1(n3926), .I2(n3929), .O(n3938) );
  NAND_GATE U5071 ( .I1(n3928), .I2(n3932), .O(n3936) );
  NAND_GATE U5072 ( .I1(n3930), .I2(n3929), .O(n3931) );
  NAND_GATE U5073 ( .I1(n3932), .I2(n3931), .O(n3933) );
  NAND_GATE U5074 ( .I1(n3934), .I2(n3933), .O(n3935) );
  NAND_GATE U5075 ( .I1(n3936), .I2(n3935), .O(n3937) );
  NAND_GATE U5076 ( .I1(n3938), .I2(n3937), .O(n4268) );
  NAND_GATE U5077 ( .I1(n3939), .I2(n4268), .O(n4264) );
  NAND_GATE U5078 ( .I1(n4269), .I2(n4268), .O(n3940) );
  NAND3_GATE U5079 ( .I1(n4265), .I2(n4264), .I3(n3940), .O(n4258) );
  NAND_GATE U5080 ( .I1(n3954), .I2(n4258), .O(n4254) );
  INV_GATE U5081 ( .I1(n3941), .O(n3942) );
  NAND_GATE U5082 ( .I1(n3942), .I2(n3945), .O(n3953) );
  NAND_GATE U5083 ( .I1(n3944), .I2(n3947), .O(n3951) );
  NAND_GATE U5084 ( .I1(n822), .I2(n3945), .O(n3946) );
  NAND_GATE U5085 ( .I1(n3947), .I2(n3946), .O(n3948) );
  NAND_GATE U5086 ( .I1(n3949), .I2(n3948), .O(n3950) );
  NAND_GATE U5087 ( .I1(n3951), .I2(n3950), .O(n3952) );
  NAND_GATE U5088 ( .I1(n3953), .I2(n3952), .O(n4257) );
  NAND_GATE U5089 ( .I1(n3954), .I2(n4257), .O(n4253) );
  NAND_GATE U5090 ( .I1(n4258), .I2(n4257), .O(n3955) );
  NAND3_GATE U5091 ( .I1(n4254), .I2(n4253), .I3(n3955), .O(n4247) );
  NAND_GATE U5092 ( .I1(n3970), .I2(n4247), .O(n4243) );
  INV_GATE U5093 ( .I1(n3956), .O(n3957) );
  NAND_GATE U5094 ( .I1(n3957), .I2(n3960), .O(n3969) );
  NAND_GATE U5095 ( .I1(n3959), .I2(n3963), .O(n3967) );
  NAND_GATE U5096 ( .I1(n3961), .I2(n3960), .O(n3962) );
  NAND_GATE U5097 ( .I1(n3963), .I2(n3962), .O(n3964) );
  NAND_GATE U5098 ( .I1(n3965), .I2(n3964), .O(n3966) );
  NAND_GATE U5099 ( .I1(n3967), .I2(n3966), .O(n3968) );
  NAND_GATE U5100 ( .I1(n3969), .I2(n3968), .O(n4246) );
  NAND_GATE U5101 ( .I1(n3970), .I2(n4246), .O(n4242) );
  NAND_GATE U5102 ( .I1(n4247), .I2(n4246), .O(n3971) );
  NAND3_GATE U5103 ( .I1(n4243), .I2(n4242), .I3(n3971), .O(n4236) );
  NAND_GATE U5104 ( .I1(n3986), .I2(n4236), .O(n4230) );
  INV_GATE U5105 ( .I1(n3972), .O(n3973) );
  NAND_GATE U5106 ( .I1(n3973), .I2(n3976), .O(n3985) );
  NAND_GATE U5107 ( .I1(n3975), .I2(n3979), .O(n3983) );
  NAND_GATE U5108 ( .I1(n3977), .I2(n3976), .O(n3978) );
  NAND_GATE U5109 ( .I1(n3979), .I2(n3978), .O(n3980) );
  NAND_GATE U5110 ( .I1(n3981), .I2(n3980), .O(n3982) );
  NAND_GATE U5111 ( .I1(n3983), .I2(n3982), .O(n3984) );
  NAND_GATE U5112 ( .I1(n3985), .I2(n3984), .O(n4234) );
  NAND_GATE U5113 ( .I1(n3986), .I2(n4234), .O(n4229) );
  NAND_GATE U5114 ( .I1(n4236), .I2(n4234), .O(n3987) );
  NAND3_GATE U5115 ( .I1(n4230), .I2(n4229), .I3(n3987), .O(n4223) );
  NAND_GATE U5116 ( .I1(n4002), .I2(n4223), .O(n4219) );
  INV_GATE U5117 ( .I1(n3988), .O(n3989) );
  NAND_GATE U5118 ( .I1(n3989), .I2(n3992), .O(n4001) );
  NAND_GATE U5119 ( .I1(n3991), .I2(n3995), .O(n3999) );
  NAND_GATE U5120 ( .I1(n3993), .I2(n3992), .O(n3994) );
  NAND_GATE U5121 ( .I1(n3995), .I2(n3994), .O(n3996) );
  NAND_GATE U5122 ( .I1(n3997), .I2(n3996), .O(n3998) );
  NAND_GATE U5123 ( .I1(n3999), .I2(n3998), .O(n4000) );
  NAND_GATE U5124 ( .I1(n4001), .I2(n4000), .O(n4222) );
  NAND_GATE U5125 ( .I1(n4002), .I2(n4222), .O(n4218) );
  NAND_GATE U5126 ( .I1(n4223), .I2(n4222), .O(n4003) );
  NAND3_GATE U5127 ( .I1(n4219), .I2(n4218), .I3(n4003), .O(n4212) );
  NAND_GATE U5128 ( .I1(n4018), .I2(n4212), .O(n4208) );
  INV_GATE U5129 ( .I1(n4004), .O(n4005) );
  NAND_GATE U5130 ( .I1(n4005), .I2(n4008), .O(n4017) );
  NAND_GATE U5131 ( .I1(n4007), .I2(n4011), .O(n4015) );
  NAND_GATE U5132 ( .I1(n4009), .I2(n4008), .O(n4010) );
  NAND_GATE U5133 ( .I1(n4011), .I2(n4010), .O(n4012) );
  NAND_GATE U5134 ( .I1(n4013), .I2(n4012), .O(n4014) );
  NAND_GATE U5135 ( .I1(n4015), .I2(n4014), .O(n4016) );
  NAND_GATE U5136 ( .I1(n4017), .I2(n4016), .O(n4211) );
  NAND_GATE U5137 ( .I1(n4018), .I2(n4211), .O(n4207) );
  NAND_GATE U5138 ( .I1(n4212), .I2(n4211), .O(n4019) );
  NAND3_GATE U5139 ( .I1(n4208), .I2(n4207), .I3(n4019), .O(n4499) );
  NAND_GATE U5140 ( .I1(n4034), .I2(n4499), .O(n4495) );
  INV_GATE U5141 ( .I1(n4020), .O(n4021) );
  NAND_GATE U5142 ( .I1(n4021), .I2(n4024), .O(n4033) );
  NAND_GATE U5143 ( .I1(n4023), .I2(n4027), .O(n4031) );
  NAND_GATE U5144 ( .I1(n4025), .I2(n4024), .O(n4026) );
  NAND_GATE U5145 ( .I1(n4027), .I2(n4026), .O(n4028) );
  NAND_GATE U5146 ( .I1(n4029), .I2(n4028), .O(n4030) );
  NAND_GATE U5147 ( .I1(n4031), .I2(n4030), .O(n4032) );
  NAND_GATE U5148 ( .I1(n4033), .I2(n4032), .O(n4498) );
  NAND_GATE U5149 ( .I1(n4034), .I2(n4498), .O(n4494) );
  NAND_GATE U5150 ( .I1(n4499), .I2(n4498), .O(n4035) );
  NAND3_GATE U5151 ( .I1(n4495), .I2(n4494), .I3(n4035), .O(n4201) );
  NAND_GATE U5152 ( .I1(n4050), .I2(n4201), .O(n4197) );
  INV_GATE U5153 ( .I1(n4036), .O(n4037) );
  NAND_GATE U5154 ( .I1(n4037), .I2(n4040), .O(n4049) );
  NAND_GATE U5155 ( .I1(n4039), .I2(n4043), .O(n4047) );
  NAND_GATE U5156 ( .I1(n4041), .I2(n4040), .O(n4042) );
  NAND_GATE U5157 ( .I1(n4043), .I2(n4042), .O(n4044) );
  NAND_GATE U5158 ( .I1(n4045), .I2(n4044), .O(n4046) );
  NAND_GATE U5159 ( .I1(n4047), .I2(n4046), .O(n4048) );
  NAND_GATE U5160 ( .I1(n4049), .I2(n4048), .O(n4200) );
  NAND_GATE U5161 ( .I1(n4050), .I2(n4200), .O(n4196) );
  NAND_GATE U5162 ( .I1(n4201), .I2(n4200), .O(n4051) );
  NAND3_GATE U5163 ( .I1(n4197), .I2(n4196), .I3(n4051), .O(n4190) );
  NAND_GATE U5164 ( .I1(n4052), .I2(n4190), .O(n4185) );
  NAND_GATE U5165 ( .I1(n4189), .I2(n4190), .O(n4053) );
  NAND3_GATE U5166 ( .I1(n4186), .I2(n4185), .I3(n4053), .O(n4179) );
  NAND_GATE U5167 ( .I1(n4068), .I2(n4179), .O(n4175) );
  INV_GATE U5168 ( .I1(n4054), .O(n4055) );
  NAND_GATE U5169 ( .I1(n4055), .I2(n4058), .O(n4067) );
  NAND_GATE U5170 ( .I1(n4057), .I2(n4061), .O(n4065) );
  NAND_GATE U5171 ( .I1(n4059), .I2(n4058), .O(n4060) );
  NAND_GATE U5172 ( .I1(n4061), .I2(n4060), .O(n4062) );
  NAND_GATE U5173 ( .I1(n4063), .I2(n4062), .O(n4064) );
  NAND_GATE U5174 ( .I1(n4065), .I2(n4064), .O(n4066) );
  NAND_GATE U5175 ( .I1(n4067), .I2(n4066), .O(n4178) );
  NAND_GATE U5176 ( .I1(n4068), .I2(n4178), .O(n4174) );
  NAND_GATE U5177 ( .I1(n4179), .I2(n4178), .O(n4069) );
  NAND3_GATE U5178 ( .I1(n4175), .I2(n4174), .I3(n4069), .O(n4168) );
  NAND_GATE U5179 ( .I1(n4084), .I2(n4168), .O(n4164) );
  OR_GATE U5180 ( .I1(n4071), .I2(n4070), .O(n4083) );
  NAND_GATE U5181 ( .I1(n4072), .I2(n4071), .O(n4077) );
  NAND_GATE U5182 ( .I1(n4073), .I2(n4077), .O(n4081) );
  NAND_GATE U5183 ( .I1(n4075), .I2(n4074), .O(n4076) );
  NAND_GATE U5184 ( .I1(n4077), .I2(n4076), .O(n4078) );
  NAND_GATE U5185 ( .I1(n4079), .I2(n4078), .O(n4080) );
  NAND_GATE U5186 ( .I1(n4081), .I2(n4080), .O(n4082) );
  NAND_GATE U5187 ( .I1(n4083), .I2(n4082), .O(n4167) );
  NAND_GATE U5188 ( .I1(n4084), .I2(n4167), .O(n4163) );
  NAND_GATE U5189 ( .I1(n4168), .I2(n4167), .O(n4085) );
  NAND3_GATE U5190 ( .I1(n4164), .I2(n4163), .I3(n4085), .O(n4157) );
  NAND_GATE U5191 ( .I1(n4100), .I2(n4157), .O(n4153) );
  INV_GATE U5192 ( .I1(n4086), .O(n4087) );
  NAND_GATE U5193 ( .I1(n4087), .I2(n4090), .O(n4099) );
  NAND_GATE U5194 ( .I1(n4089), .I2(n4093), .O(n4097) );
  NAND_GATE U5195 ( .I1(n4091), .I2(n4090), .O(n4092) );
  NAND_GATE U5196 ( .I1(n4093), .I2(n4092), .O(n4094) );
  NAND_GATE U5197 ( .I1(n4095), .I2(n4094), .O(n4096) );
  NAND_GATE U5198 ( .I1(n4097), .I2(n4096), .O(n4098) );
  NAND_GATE U5199 ( .I1(n4099), .I2(n4098), .O(n4156) );
  NAND_GATE U5200 ( .I1(n4100), .I2(n4156), .O(n4152) );
  NAND_GATE U5201 ( .I1(n4157), .I2(n4156), .O(n4101) );
  NAND3_GATE U5202 ( .I1(n4153), .I2(n4152), .I3(n4101), .O(n4146) );
  NAND_GATE U5203 ( .I1(n4116), .I2(n4146), .O(n4142) );
  INV_GATE U5204 ( .I1(n4102), .O(n4103) );
  NAND_GATE U5205 ( .I1(n4103), .I2(n4106), .O(n4115) );
  NAND_GATE U5206 ( .I1(n4105), .I2(n4109), .O(n4113) );
  NAND_GATE U5207 ( .I1(n4107), .I2(n4106), .O(n4108) );
  NAND_GATE U5208 ( .I1(n4109), .I2(n4108), .O(n4110) );
  NAND_GATE U5209 ( .I1(n4111), .I2(n4110), .O(n4112) );
  NAND_GATE U5210 ( .I1(n4113), .I2(n4112), .O(n4114) );
  NAND_GATE U5211 ( .I1(n4115), .I2(n4114), .O(n4145) );
  NAND_GATE U5212 ( .I1(n4116), .I2(n4145), .O(n4141) );
  NAND_GATE U5213 ( .I1(n4146), .I2(n4145), .O(n4117) );
  NAND3_GATE U5214 ( .I1(n4142), .I2(n4141), .I3(n4117), .O(n4135) );
  NAND_GATE U5215 ( .I1(n4135), .I2(n4134), .O(n4119) );
  NAND_GATE U5216 ( .I1(n4118), .I2(n4135), .O(n4131) );
  AND3_GATE U5217 ( .I1(n4130), .I2(n4119), .I3(n4131), .O(n4126) );
  NAND_GATE U5218 ( .I1(n1436), .I2(A[31]), .O(n4125) );
  NAND_GATE U5219 ( .I1(n4126), .I2(n4125), .O(n4120) );
  NAND_GATE U5220 ( .I1(n4124), .I2(n4120), .O(n4129) );
  NAND_GATE U5221 ( .I1(n14791), .I2(n4129), .O(n4123) );
  INV_GATE U5222 ( .I1(n4129), .O(n14790) );
  NAND_GATE U5223 ( .I1(n4121), .I2(n14790), .O(n4122) );
  NAND_GATE U5224 ( .I1(n4123), .I2(n4122), .O(\A1[54] ) );
  INV_GATE U5225 ( .I1(n4124), .O(n4127) );
  NAND3_GATE U5226 ( .I1(n4127), .I2(n4126), .I3(n4125), .O(n4128) );
  NAND_GATE U5227 ( .I1(n4129), .I2(n4128), .O(n4520) );
  INV_GATE U5228 ( .I1(n4520), .O(n14793) );
  OR_GATE U5229 ( .I1(n4130), .I2(n4135), .O(n4133) );
  OR_GATE U5230 ( .I1(n4134), .I2(n4131), .O(n4132) );
  AND_GATE U5231 ( .I1(n4133), .I2(n4132), .O(n4140) );
  NAND_GATE U5232 ( .I1(n4135), .I2(n1199), .O(n4137) );
  NAND3_GATE U5233 ( .I1(n4138), .I2(n4137), .I3(n4136), .O(n4139) );
  OR_GATE U5234 ( .I1(n4141), .I2(n4146), .O(n4144) );
  OR_GATE U5235 ( .I1(n4145), .I2(n4142), .O(n4143) );
  AND_GATE U5236 ( .I1(n4144), .I2(n4143), .O(n4151) );
  NAND_GATE U5237 ( .I1(n4146), .I2(n1197), .O(n4148) );
  NAND3_GATE U5238 ( .I1(n4149), .I2(n4148), .I3(n4147), .O(n4150) );
  NAND_GATE U5239 ( .I1(n4151), .I2(n4150), .O(n4528) );
  INV_GATE U5240 ( .I1(n4528), .O(n4531) );
  NAND_GATE U5241 ( .I1(B[23]), .I2(A[30]), .O(n4535) );
  INV_GATE U5242 ( .I1(n4535), .O(n4529) );
  NAND_GATE U5243 ( .I1(n4531), .I2(n4529), .O(n4526) );
  OR_GATE U5244 ( .I1(n4152), .I2(n4157), .O(n4155) );
  OR_GATE U5245 ( .I1(n4156), .I2(n4153), .O(n4154) );
  AND_GATE U5246 ( .I1(n4155), .I2(n4154), .O(n4162) );
  NAND_GATE U5247 ( .I1(n1188), .I2(n4156), .O(n4160) );
  NAND3_GATE U5248 ( .I1(n4160), .I2(n4159), .I3(n4158), .O(n4161) );
  NAND_GATE U5249 ( .I1(n4162), .I2(n4161), .O(n4543) );
  INV_GATE U5250 ( .I1(n4543), .O(n4546) );
  NAND_GATE U5251 ( .I1(B[23]), .I2(A[29]), .O(n4550) );
  INV_GATE U5252 ( .I1(n4550), .O(n4544) );
  NAND_GATE U5253 ( .I1(n4546), .I2(n4544), .O(n4540) );
  OR_GATE U5254 ( .I1(n4163), .I2(n4168), .O(n4166) );
  OR_GATE U5255 ( .I1(n4167), .I2(n4164), .O(n4165) );
  AND_GATE U5256 ( .I1(n4166), .I2(n4165), .O(n4173) );
  NAND_GATE U5257 ( .I1(n1182), .I2(n4167), .O(n4171) );
  NAND3_GATE U5258 ( .I1(n4171), .I2(n4170), .I3(n4169), .O(n4172) );
  NAND_GATE U5259 ( .I1(n4173), .I2(n4172), .O(n4967) );
  INV_GATE U5260 ( .I1(n4967), .O(n4970) );
  NAND_GATE U5261 ( .I1(B[23]), .I2(A[28]), .O(n4974) );
  INV_GATE U5262 ( .I1(n4974), .O(n4968) );
  NAND_GATE U5263 ( .I1(n4970), .I2(n4968), .O(n4965) );
  OR_GATE U5264 ( .I1(n4174), .I2(n4179), .O(n4177) );
  OR_GATE U5265 ( .I1(n4178), .I2(n4175), .O(n4176) );
  AND_GATE U5266 ( .I1(n4177), .I2(n4176), .O(n4184) );
  NAND_GATE U5267 ( .I1(n1178), .I2(n4178), .O(n4182) );
  NAND3_GATE U5268 ( .I1(n4182), .I2(n4181), .I3(n4180), .O(n4183) );
  NAND_GATE U5269 ( .I1(n4184), .I2(n4183), .O(n4951) );
  INV_GATE U5270 ( .I1(n4951), .O(n4954) );
  NAND_GATE U5271 ( .I1(B[23]), .I2(A[27]), .O(n4958) );
  INV_GATE U5272 ( .I1(n4958), .O(n4952) );
  NAND_GATE U5273 ( .I1(n4954), .I2(n4952), .O(n4949) );
  OR_GATE U5274 ( .I1(n4185), .I2(n4189), .O(n4188) );
  OR_GATE U5275 ( .I1(n4190), .I2(n4186), .O(n4187) );
  AND_GATE U5276 ( .I1(n4188), .I2(n4187), .O(n4195) );
  NAND_GATE U5277 ( .I1(n1172), .I2(n4190), .O(n4192) );
  NAND3_GATE U5278 ( .I1(n4193), .I2(n4192), .I3(n4191), .O(n4194) );
  NAND_GATE U5279 ( .I1(n4195), .I2(n4194), .O(n4935) );
  INV_GATE U5280 ( .I1(n4935), .O(n4938) );
  NAND_GATE U5281 ( .I1(B[23]), .I2(A[26]), .O(n4942) );
  INV_GATE U5282 ( .I1(n4942), .O(n4936) );
  NAND_GATE U5283 ( .I1(n4938), .I2(n4936), .O(n4933) );
  OR_GATE U5284 ( .I1(n4196), .I2(n4201), .O(n4199) );
  OR_GATE U5285 ( .I1(n4200), .I2(n4197), .O(n4198) );
  AND_GATE U5286 ( .I1(n4199), .I2(n4198), .O(n4206) );
  NAND_GATE U5287 ( .I1(n1164), .I2(n4200), .O(n4204) );
  NAND3_GATE U5288 ( .I1(n4204), .I2(n4203), .I3(n4202), .O(n4205) );
  NAND_GATE U5289 ( .I1(n4206), .I2(n4205), .O(n4919) );
  INV_GATE U5290 ( .I1(n4919), .O(n4922) );
  NAND_GATE U5291 ( .I1(B[23]), .I2(A[25]), .O(n4926) );
  INV_GATE U5292 ( .I1(n4926), .O(n4920) );
  NAND_GATE U5293 ( .I1(n4922), .I2(n4920), .O(n4917) );
  NAND_GATE U5294 ( .I1(B[23]), .I2(A[24]), .O(n4910) );
  INV_GATE U5295 ( .I1(n4910), .O(n4904) );
  OR_GATE U5296 ( .I1(n4207), .I2(n4212), .O(n4210) );
  OR_GATE U5297 ( .I1(n4211), .I2(n4208), .O(n4209) );
  AND_GATE U5298 ( .I1(n4210), .I2(n4209), .O(n4217) );
  NAND_GATE U5299 ( .I1(n1123), .I2(n4211), .O(n4215) );
  NAND3_GATE U5300 ( .I1(n4215), .I2(n4214), .I3(n4213), .O(n4216) );
  NAND_GATE U5301 ( .I1(n4217), .I2(n4216), .O(n4887) );
  INV_GATE U5302 ( .I1(n4887), .O(n4890) );
  NAND_GATE U5303 ( .I1(B[23]), .I2(A[23]), .O(n4894) );
  INV_GATE U5304 ( .I1(n4894), .O(n4888) );
  NAND_GATE U5305 ( .I1(n4890), .I2(n4888), .O(n4885) );
  OR_GATE U5306 ( .I1(n4218), .I2(n4223), .O(n4221) );
  OR_GATE U5307 ( .I1(n4222), .I2(n4219), .O(n4220) );
  AND_GATE U5308 ( .I1(n4221), .I2(n4220), .O(n4228) );
  NAND_GATE U5309 ( .I1(n1121), .I2(n4222), .O(n4226) );
  NAND3_GATE U5310 ( .I1(n4226), .I2(n4225), .I3(n4224), .O(n4227) );
  NAND_GATE U5311 ( .I1(n4228), .I2(n4227), .O(n4557) );
  INV_GATE U5312 ( .I1(n4557), .O(n4560) );
  NAND_GATE U5313 ( .I1(B[23]), .I2(A[22]), .O(n4564) );
  INV_GATE U5314 ( .I1(n4564), .O(n4558) );
  NAND_GATE U5315 ( .I1(n4560), .I2(n4558), .O(n4555) );
  OR_GATE U5316 ( .I1(n4229), .I2(n4236), .O(n4232) );
  OR_GATE U5317 ( .I1(n4234), .I2(n4230), .O(n4231) );
  AND_GATE U5318 ( .I1(n4232), .I2(n4231), .O(n4241) );
  INV_GATE U5319 ( .I1(n4236), .O(n4233) );
  NAND_GATE U5320 ( .I1(n4233), .I2(n4234), .O(n4239) );
  INV_GATE U5321 ( .I1(n4234), .O(n4235) );
  NAND_GATE U5322 ( .I1(n4236), .I2(n4235), .O(n4238) );
  NAND3_GATE U5323 ( .I1(n4239), .I2(n4238), .I3(n4237), .O(n4240) );
  NAND_GATE U5324 ( .I1(n4241), .I2(n4240), .O(n4869) );
  INV_GATE U5325 ( .I1(n4869), .O(n4872) );
  NAND_GATE U5326 ( .I1(B[23]), .I2(A[21]), .O(n4876) );
  INV_GATE U5327 ( .I1(n4876), .O(n4870) );
  NAND_GATE U5328 ( .I1(n4872), .I2(n4870), .O(n4867) );
  OR_GATE U5329 ( .I1(n4242), .I2(n4247), .O(n4245) );
  OR_GATE U5330 ( .I1(n4246), .I2(n4243), .O(n4244) );
  AND_GATE U5331 ( .I1(n4245), .I2(n4244), .O(n4252) );
  NAND_GATE U5332 ( .I1(n1148), .I2(n4246), .O(n4250) );
  NAND3_GATE U5333 ( .I1(n4250), .I2(n4249), .I3(n4248), .O(n4251) );
  NAND_GATE U5334 ( .I1(n4252), .I2(n4251), .O(n4853) );
  INV_GATE U5335 ( .I1(n4853), .O(n4856) );
  NAND_GATE U5336 ( .I1(B[23]), .I2(A[20]), .O(n4860) );
  INV_GATE U5337 ( .I1(n4860), .O(n4854) );
  NAND_GATE U5338 ( .I1(n4856), .I2(n4854), .O(n4851) );
  OR_GATE U5339 ( .I1(n4253), .I2(n4258), .O(n4256) );
  OR_GATE U5340 ( .I1(n4257), .I2(n4254), .O(n4255) );
  AND_GATE U5341 ( .I1(n4256), .I2(n4255), .O(n4263) );
  NAND_GATE U5342 ( .I1(n1149), .I2(n4257), .O(n4261) );
  NAND3_GATE U5343 ( .I1(n4261), .I2(n4260), .I3(n4259), .O(n4262) );
  NAND_GATE U5344 ( .I1(n4263), .I2(n4262), .O(n4837) );
  INV_GATE U5345 ( .I1(n4837), .O(n4840) );
  NAND_GATE U5346 ( .I1(B[23]), .I2(A[19]), .O(n4844) );
  INV_GATE U5347 ( .I1(n4844), .O(n4838) );
  NAND_GATE U5348 ( .I1(n4840), .I2(n4838), .O(n4835) );
  OR_GATE U5349 ( .I1(n4264), .I2(n4269), .O(n4267) );
  OR_GATE U5350 ( .I1(n4268), .I2(n4265), .O(n4266) );
  AND_GATE U5351 ( .I1(n4267), .I2(n4266), .O(n4274) );
  NAND_GATE U5352 ( .I1(n723), .I2(n4268), .O(n4272) );
  NAND3_GATE U5353 ( .I1(n4272), .I2(n4271), .I3(n4270), .O(n4273) );
  NAND_GATE U5354 ( .I1(B[23]), .I2(A[18]), .O(n4828) );
  INV_GATE U5355 ( .I1(n4828), .O(n4823) );
  NAND_GATE U5356 ( .I1(n801), .I2(n4823), .O(n4820) );
  OR_GATE U5357 ( .I1(n4275), .I2(n4280), .O(n4278) );
  OR_GATE U5358 ( .I1(n4279), .I2(n4276), .O(n4277) );
  AND_GATE U5359 ( .I1(n4278), .I2(n4277), .O(n4285) );
  NAND_GATE U5360 ( .I1(n1124), .I2(n4279), .O(n4283) );
  NAND3_GATE U5361 ( .I1(n4283), .I2(n4282), .I3(n4281), .O(n4284) );
  NAND_GATE U5362 ( .I1(n4285), .I2(n4284), .O(n4807) );
  NAND_GATE U5363 ( .I1(B[23]), .I2(A[17]), .O(n4813) );
  INV_GATE U5364 ( .I1(n4813), .O(n4808) );
  NAND_GATE U5365 ( .I1(n313), .I2(n4808), .O(n4805) );
  OR_GATE U5366 ( .I1(n4290), .I2(n4287), .O(n4288) );
  AND_GATE U5367 ( .I1(n4289), .I2(n4288), .O(n4296) );
  NAND_GATE U5368 ( .I1(n1116), .I2(n4290), .O(n4294) );
  NAND3_GATE U5369 ( .I1(n4294), .I2(n4293), .I3(n4292), .O(n4295) );
  NAND_GATE U5370 ( .I1(n4296), .I2(n4295), .O(n4797) );
  NAND_GATE U5371 ( .I1(B[23]), .I2(A[16]), .O(n4800) );
  INV_GATE U5372 ( .I1(n4800), .O(n4794) );
  OR_GATE U5373 ( .I1(n4297), .I2(n4302), .O(n4300) );
  OR_GATE U5374 ( .I1(n4301), .I2(n4298), .O(n4299) );
  AND_GATE U5375 ( .I1(n4300), .I2(n4299), .O(n4307) );
  NAND_GATE U5376 ( .I1(n1094), .I2(n4301), .O(n4305) );
  NAND3_GATE U5377 ( .I1(n4305), .I2(n4304), .I3(n4303), .O(n4306) );
  NAND_GATE U5378 ( .I1(n4307), .I2(n4306), .O(n4781) );
  NAND_GATE U5379 ( .I1(B[23]), .I2(A[15]), .O(n4785) );
  INV_GATE U5380 ( .I1(n4785), .O(n4779) );
  NAND_GATE U5381 ( .I1(B[23]), .I2(A[14]), .O(n4569) );
  INV_GATE U5382 ( .I1(n4569), .O(n4572) );
  NAND_GATE U5383 ( .I1(n1394), .I2(n4314), .O(n4309) );
  NAND3_GATE U5384 ( .I1(n4310), .I2(n4309), .I3(n4308), .O(n4317) );
  OR_GATE U5385 ( .I1(n4312), .I2(n4311), .O(n4316) );
  OR_GATE U5386 ( .I1(n4314), .I2(n4313), .O(n4315) );
  NAND3_GATE U5387 ( .I1(n4317), .I2(n4316), .I3(n4315), .O(n4570) );
  NAND_GATE U5388 ( .I1(n4572), .I2(n903), .O(n4575) );
  NAND_GATE U5389 ( .I1(B[23]), .I2(A[13]), .O(n4765) );
  INV_GATE U5390 ( .I1(n4765), .O(n4761) );
  OR_GATE U5391 ( .I1(n4322), .I2(n4318), .O(n4321) );
  OR_GATE U5392 ( .I1(n4319), .I2(n4323), .O(n4320) );
  AND_GATE U5393 ( .I1(n4321), .I2(n4320), .O(n4328) );
  NAND_GATE U5394 ( .I1(n333), .I2(n4322), .O(n4325) );
  NAND3_GATE U5395 ( .I1(n4326), .I2(n4325), .I3(n4324), .O(n4327) );
  NAND_GATE U5396 ( .I1(n4328), .I2(n4327), .O(n4762) );
  NAND_GATE U5397 ( .I1(n4761), .I2(n905), .O(n4768) );
  NAND_GATE U5398 ( .I1(B[23]), .I2(A[12]), .O(n4750) );
  INV_GATE U5399 ( .I1(n4750), .O(n4745) );
  NAND_GATE U5400 ( .I1(n4332), .I2(n1266), .O(n4330) );
  NAND3_GATE U5401 ( .I1(n4331), .I2(n4330), .I3(n4329), .O(n4337) );
  OR_GATE U5402 ( .I1(n4333), .I2(n4332), .O(n4336) );
  OR_GATE U5403 ( .I1(n811), .I2(n4334), .O(n4335) );
  NAND3_GATE U5404 ( .I1(n4337), .I2(n4336), .I3(n4335), .O(n4746) );
  NAND_GATE U5405 ( .I1(n4745), .I2(n810), .O(n4753) );
  NAND_GATE U5406 ( .I1(B[23]), .I2(A[10]), .O(n4720) );
  INV_GATE U5407 ( .I1(n4720), .O(n4727) );
  NAND_GATE U5408 ( .I1(n303), .I2(n4339), .O(n4440) );
  AND3_GATE U5409 ( .I1(n4440), .I2(n4442), .I3(n4441), .O(n4344) );
  OR_GATE U5410 ( .I1(n4339), .I2(n4458), .O(n4343) );
  NAND4_GATE U5411 ( .I1(n4341), .I2(n1212), .I3(n4340), .I4(n303), .O(n4342)
         );
  NAND_GATE U5412 ( .I1(n4343), .I2(n4342), .O(n4439) );
  OR_GATE U5413 ( .I1(n4344), .I2(n4439), .O(n4722) );
  INV_GATE U5414 ( .I1(n4722), .O(n4718) );
  NAND_GATE U5415 ( .I1(n4727), .I2(n4718), .O(n4446) );
  NAND_GATE U5416 ( .I1(B[23]), .I2(A[9]), .O(n4596) );
  INV_GATE U5417 ( .I1(n4596), .O(n4588) );
  NAND_GATE U5418 ( .I1(B[23]), .I2(A[8]), .O(n5202) );
  INV_GATE U5419 ( .I1(n5202), .O(n4709) );
  NAND4_GATE U5420 ( .I1(n4346), .I2(n4345), .I3(n4356), .I4(n386), .O(n4701)
         );
  NAND_GATE U5421 ( .I1(n4350), .I2(n4349), .O(n4356) );
  NAND_GATE U5422 ( .I1(n4352), .I2(n746), .O(n4355) );
  NAND_GATE U5423 ( .I1(n4356), .I2(n4355), .O(n4353) );
  NAND_GATE U5424 ( .I1(n4354), .I2(n4353), .O(n4359) );
  NAND3_GATE U5425 ( .I1(n4356), .I2(n4355), .I3(n386), .O(n4358) );
  NAND3_GATE U5426 ( .I1(n4359), .I2(n4358), .I3(n4357), .O(n4700) );
  NAND_GATE U5427 ( .I1(n4709), .I2(n1301), .O(n4432) );
  NAND_GATE U5428 ( .I1(B[23]), .I2(A[7]), .O(n4614) );
  INV_GATE U5429 ( .I1(n4614), .O(n4606) );
  NAND_GATE U5430 ( .I1(B[23]), .I2(A[6]), .O(n4687) );
  INV_GATE U5431 ( .I1(n4687), .O(n5298) );
  NAND_GATE U5432 ( .I1(n4362), .I2(n3805), .O(n4364) );
  NAND_GATE U5433 ( .I1(n4368), .I2(n4367), .O(n4363) );
  NAND_GATE U5434 ( .I1(n4364), .I2(n4363), .O(n4366) );
  NAND3_GATE U5435 ( .I1(n4366), .I2(n4365), .I3(n1256), .O(n4413) );
  INV_GATE U5436 ( .I1(n4372), .O(n4369) );
  NAND3_GATE U5437 ( .I1(n4369), .I2(n4363), .I3(n1216), .O(n4412) );
  NAND3_GATE U5438 ( .I1(n4369), .I2(n4370), .I3(n4363), .O(n4415) );
  NAND_GATE U5439 ( .I1(n4370), .I2(n4363), .O(n4371) );
  NAND_GATE U5440 ( .I1(n4372), .I2(n4371), .O(n4416) );
  NAND3_GATE U5441 ( .I1(n4417), .I2(n4415), .I3(n4416), .O(n5299) );
  NAND_GATE U5442 ( .I1(n1214), .I2(n5299), .O(n4688) );
  INV_GATE U5443 ( .I1(n4688), .O(n4691) );
  NAND_GATE U5444 ( .I1(n5298), .I2(n4691), .O(n4421) );
  NAND_GATE U5445 ( .I1(B[23]), .I2(A[5]), .O(n4627) );
  INV_GATE U5446 ( .I1(n4627), .O(n4409) );
  NAND_GATE U5447 ( .I1(B[23]), .I2(A[4]), .O(n5273) );
  OR_GATE U5448 ( .I1(n4380), .I2(n4373), .O(n4379) );
  INV_GATE U5449 ( .I1(n4383), .O(n4381) );
  NAND5_GATE U5450 ( .I1(n4377), .I2(n4376), .I3(n4381), .I4(n4375), .I5(n4374), .O(n4378) );
  NAND_GATE U5451 ( .I1(n4379), .I2(n4378), .O(n4398) );
  NAND_GATE U5452 ( .I1(n5273), .I2(n4398), .O(n4397) );
  NAND_GATE U5453 ( .I1(n4381), .I2(n4380), .O(n4399) );
  NAND3_GATE U5454 ( .I1(n4384), .I2(n4383), .I3(n4382), .O(n4385) );
  AND_GATE U5455 ( .I1(n4386), .I2(n4385), .O(n4400) );
  NAND3_GATE U5456 ( .I1(n5273), .I2(n4399), .I3(n4400), .O(n4396) );
  NAND_GATE U5457 ( .I1(B[23]), .I2(A[3]), .O(n4659) );
  INV_GATE U5458 ( .I1(n4659), .O(n4671) );
  NAND_GATE U5459 ( .I1(B[23]), .I2(A[2]), .O(n4647) );
  INV_GATE U5460 ( .I1(n4647), .O(n4645) );
  NAND_GATE U5461 ( .I1(n1436), .I2(A[0]), .O(n4387) );
  NAND_GATE U5462 ( .I1(n14241), .I2(n4387), .O(n4388) );
  NAND_GATE U5463 ( .I1(B[25]), .I2(n4388), .O(n4642) );
  NAND_GATE U5464 ( .I1(n1437), .I2(A[1]), .O(n4389) );
  NAND_GATE U5465 ( .I1(n724), .I2(n4389), .O(n4390) );
  NAND_GATE U5466 ( .I1(B[24]), .I2(n4390), .O(n4643) );
  NAND_GATE U5467 ( .I1(n4642), .I2(n4643), .O(n4650) );
  NAND_GATE U5468 ( .I1(n4645), .I2(n4650), .O(n4641) );
  NAND3_GATE U5469 ( .I1(B[23]), .I2(B[24]), .I3(n1254), .O(n4646) );
  INV_GATE U5470 ( .I1(n4646), .O(n4649) );
  NAND_GATE U5471 ( .I1(n4647), .I2(n4643), .O(n4391) );
  NAND_GATE U5472 ( .I1(n4649), .I2(n4391), .O(n4392) );
  NAND_GATE U5473 ( .I1(n4641), .I2(n4392), .O(n4657) );
  NAND_GATE U5474 ( .I1(n4671), .I2(n4657), .O(n4667) );
  NAND_GATE U5475 ( .I1(n414), .I2(n4393), .O(n4669) );
  NAND3_GATE U5476 ( .I1(n4662), .I2(n4669), .I3(n4663), .O(n4673) );
  NAND_GATE U5477 ( .I1(n4662), .I2(n4669), .O(n4664) );
  NAND3_GATE U5478 ( .I1(n4657), .I2(n4673), .I3(n4658), .O(n4395) );
  NAND3_GATE U5479 ( .I1(n4671), .I2(n4673), .I3(n4658), .O(n4394) );
  NAND3_GATE U5480 ( .I1(n4667), .I2(n4395), .I3(n4394), .O(n5270) );
  NAND3_GATE U5481 ( .I1(n4397), .I2(n4396), .I3(n5270), .O(n4402) );
  INV_GATE U5482 ( .I1(n5273), .O(n5261) );
  INV_GATE U5483 ( .I1(n4398), .O(n5262) );
  NAND_GATE U5484 ( .I1(n4400), .I2(n4399), .O(n5263) );
  NAND_GATE U5485 ( .I1(n5262), .I2(n5263), .O(n5268) );
  NAND_GATE U5486 ( .I1(n5261), .I2(n676), .O(n4401) );
  NAND_GATE U5487 ( .I1(n4402), .I2(n4401), .O(n4624) );
  NAND_GATE U5488 ( .I1(n4409), .I2(n4624), .O(n4619) );
  INV_GATE U5489 ( .I1(n4406), .O(n4405) );
  NAND3_GATE U5490 ( .I1(n4403), .I2(n4406), .I3(n389), .O(n4620) );
  NAND_GATE U5491 ( .I1(n760), .I2(n4620), .O(n4626) );
  NAND_GATE U5492 ( .I1(n4405), .I2(n4404), .O(n4408) );
  NAND_GATE U5493 ( .I1(n4406), .I2(n389), .O(n4407) );
  NAND_GATE U5494 ( .I1(n4408), .I2(n4407), .O(n4615) );
  NAND3_GATE U5495 ( .I1(n4624), .I2(n4626), .I3(n4617), .O(n4411) );
  NAND_GATE U5496 ( .I1(n4617), .I2(n1217), .O(n4410) );
  NAND3_GATE U5497 ( .I1(n4619), .I2(n4411), .I3(n4410), .O(n4689) );
  NAND_GATE U5498 ( .I1(n4413), .I2(n4412), .O(n4414) );
  NAND_GATE U5499 ( .I1(n4687), .I2(n4414), .O(n4419) );
  NAND4_GATE U5500 ( .I1(n4417), .I2(n4416), .I3(n4687), .I4(n4415), .O(n4418)
         );
  NAND3_GATE U5501 ( .I1(n4689), .I2(n4419), .I3(n4418), .O(n4420) );
  NAND_GATE U5502 ( .I1(n4421), .I2(n4420), .O(n4611) );
  NAND_GATE U5503 ( .I1(n4606), .I2(n4611), .O(n4603) );
  INV_GATE U5504 ( .I1(n4425), .O(n4423) );
  NAND_GATE U5505 ( .I1(n4422), .I2(n4428), .O(n4602) );
  NAND3_GATE U5506 ( .I1(n4422), .I2(n4425), .I3(n4426), .O(n4607) );
  NAND_GATE U5507 ( .I1(n4424), .I2(n4423), .O(n4428) );
  NAND_GATE U5508 ( .I1(n4426), .I2(n4425), .O(n4427) );
  NAND_GATE U5509 ( .I1(n4428), .I2(n4427), .O(n4608) );
  NAND3_GATE U5510 ( .I1(n4606), .I2(n4605), .I3(n4601), .O(n4430) );
  NAND3_GATE U5511 ( .I1(n4611), .I2(n4605), .I3(n4601), .O(n4429) );
  NAND3_GATE U5512 ( .I1(n4603), .I2(n4430), .I3(n4429), .O(n4705) );
  NAND4_GATE U5513 ( .I1(n4701), .I2(n4702), .I3(n4705), .I4(n4700), .O(n4431)
         );
  NAND_GATE U5514 ( .I1(n4709), .I2(n4705), .O(n4704) );
  NAND3_GATE U5515 ( .I1(n4432), .I2(n4431), .I3(n4704), .O(n4592) );
  NAND_GATE U5516 ( .I1(n4588), .I2(n4592), .O(n4584) );
  INV_GATE U5517 ( .I1(n4434), .O(n4433) );
  NAND3_GATE U5518 ( .I1(n4580), .I2(n4434), .I3(n1268), .O(n4586) );
  NAND3_GATE U5519 ( .I1(n4436), .I2(n4586), .I3(n4580), .O(n4594) );
  NAND_GATE U5520 ( .I1(n744), .I2(n4433), .O(n4436) );
  NAND_GATE U5521 ( .I1(n1268), .I2(n4434), .O(n4435) );
  NAND_GATE U5522 ( .I1(n4436), .I2(n4435), .O(n4581) );
  NAND_GATE U5523 ( .I1(n4582), .I2(n4581), .O(n4593) );
  NAND3_GATE U5524 ( .I1(n4588), .I2(n4594), .I3(n4593), .O(n4438) );
  NAND3_GATE U5525 ( .I1(n4594), .I2(n4593), .I3(n4592), .O(n4437) );
  NAND3_GATE U5526 ( .I1(n4584), .I2(n4438), .I3(n4437), .O(n4719) );
  NAND_GATE U5527 ( .I1(n4720), .I2(n4439), .O(n4444) );
  NAND4_GATE U5528 ( .I1(n4442), .I2(n4441), .I3(n4720), .I4(n4440), .O(n4443)
         );
  NAND3_GATE U5529 ( .I1(n4719), .I2(n4444), .I3(n4443), .O(n4445) );
  NAND_GATE U5530 ( .I1(B[23]), .I2(A[11]), .O(n5174) );
  OR_GATE U5531 ( .I1(n4447), .I2(n4456), .O(n4451) );
  NAND4_GATE U5532 ( .I1(n4452), .I2(n4449), .I3(n4448), .I4(n4456), .O(n4450)
         );
  AND_GATE U5533 ( .I1(n4451), .I2(n4450), .O(n4466) );
  NAND_GATE U5534 ( .I1(n4452), .I2(n1280), .O(n4460) );
  NAND_GATE U5535 ( .I1(n4454), .I2(n4453), .O(n4459) );
  NAND_GATE U5536 ( .I1(n4460), .I2(n4459), .O(n4455) );
  NAND_GATE U5537 ( .I1(n4456), .I2(n4455), .O(n4463) );
  NAND5_GATE U5538 ( .I1(n4461), .I2(n4460), .I3(n4459), .I4(n4458), .I5(n4457), .O(n4462) );
  NAND3_GATE U5539 ( .I1(n4464), .I2(n4463), .I3(n4462), .O(n4465) );
  NAND_GATE U5540 ( .I1(n4466), .I2(n4465), .O(n4736) );
  NAND_GATE U5541 ( .I1(n5174), .I2(n4736), .O(n4467) );
  NAND_GATE U5542 ( .I1(n308), .I2(n4467), .O(n4469) );
  INV_GATE U5543 ( .I1(n5174), .O(n4738) );
  INV_GATE U5544 ( .I1(n4736), .O(n4737) );
  NAND_GATE U5545 ( .I1(n4738), .I2(n4737), .O(n4468) );
  NAND_GATE U5546 ( .I1(n4469), .I2(n4468), .O(n4754) );
  NAND_GATE U5547 ( .I1(n4750), .I2(n4746), .O(n4470) );
  NAND_GATE U5548 ( .I1(n4754), .I2(n4470), .O(n4471) );
  NAND_GATE U5549 ( .I1(n4753), .I2(n4471), .O(n4769) );
  NAND_GATE U5550 ( .I1(n4765), .I2(n4762), .O(n4472) );
  NAND_GATE U5551 ( .I1(n4769), .I2(n4472), .O(n4473) );
  NAND_GATE U5552 ( .I1(n4768), .I2(n4473), .O(n4576) );
  NAND_GATE U5553 ( .I1(n4569), .I2(n4570), .O(n4474) );
  NAND_GATE U5554 ( .I1(n4576), .I2(n4474), .O(n4475) );
  NAND_GATE U5555 ( .I1(n4781), .I2(n4785), .O(n4476) );
  NAND_GATE U5556 ( .I1(n4780), .I2(n4476), .O(n4477) );
  NAND_GATE U5557 ( .I1(n4777), .I2(n4477), .O(n4795) );
  NAND_GATE U5558 ( .I1(n4797), .I2(n4800), .O(n4478) );
  NAND_GATE U5559 ( .I1(n4795), .I2(n4478), .O(n4479) );
  NAND_GATE U5560 ( .I1(n4792), .I2(n4479), .O(n4809) );
  NAND_GATE U5561 ( .I1(n4807), .I2(n4813), .O(n4480) );
  NAND_GATE U5562 ( .I1(n4809), .I2(n4480), .O(n4481) );
  NAND_GATE U5563 ( .I1(n4805), .I2(n4481), .O(n4824) );
  NAND_GATE U5564 ( .I1(n4822), .I2(n4828), .O(n4482) );
  NAND_GATE U5565 ( .I1(n4824), .I2(n4482), .O(n4483) );
  NAND_GATE U5566 ( .I1(n4820), .I2(n4483), .O(n4839) );
  NAND_GATE U5567 ( .I1(n4837), .I2(n4844), .O(n4484) );
  NAND_GATE U5568 ( .I1(n4839), .I2(n4484), .O(n4485) );
  NAND_GATE U5569 ( .I1(n4835), .I2(n4485), .O(n4855) );
  NAND_GATE U5570 ( .I1(n4853), .I2(n4860), .O(n4486) );
  NAND_GATE U5571 ( .I1(n4855), .I2(n4486), .O(n4487) );
  NAND_GATE U5572 ( .I1(n4851), .I2(n4487), .O(n4871) );
  NAND_GATE U5573 ( .I1(n4869), .I2(n4876), .O(n4488) );
  NAND_GATE U5574 ( .I1(n4871), .I2(n4488), .O(n4489) );
  NAND_GATE U5575 ( .I1(n4867), .I2(n4489), .O(n4559) );
  NAND_GATE U5576 ( .I1(n4557), .I2(n4564), .O(n4490) );
  NAND_GATE U5577 ( .I1(n4559), .I2(n4490), .O(n4491) );
  NAND_GATE U5578 ( .I1(n4555), .I2(n4491), .O(n4889) );
  NAND_GATE U5579 ( .I1(n4887), .I2(n4894), .O(n4492) );
  NAND_GATE U5580 ( .I1(n4889), .I2(n4492), .O(n4493) );
  NAND_GATE U5581 ( .I1(n4885), .I2(n4493), .O(n4906) );
  NAND_GATE U5582 ( .I1(n4904), .I2(n4906), .O(n4901) );
  OR_GATE U5583 ( .I1(n4494), .I2(n4499), .O(n4497) );
  OR_GATE U5584 ( .I1(n4498), .I2(n4495), .O(n4496) );
  AND_GATE U5585 ( .I1(n4497), .I2(n4496), .O(n4504) );
  NAND_GATE U5586 ( .I1(n1150), .I2(n4498), .O(n4502) );
  NAND3_GATE U5587 ( .I1(n4502), .I2(n4501), .I3(n4500), .O(n4503) );
  NAND_GATE U5588 ( .I1(n4504), .I2(n4503), .O(n4902) );
  INV_GATE U5589 ( .I1(n4902), .O(n4905) );
  INV_GATE U5590 ( .I1(n4906), .O(n4903) );
  NAND_GATE U5591 ( .I1(n4910), .I2(n4903), .O(n4505) );
  NAND_GATE U5592 ( .I1(n4905), .I2(n4505), .O(n4506) );
  NAND_GATE U5593 ( .I1(n4901), .I2(n4506), .O(n4921) );
  NAND_GATE U5594 ( .I1(n4919), .I2(n4926), .O(n4507) );
  NAND_GATE U5595 ( .I1(n4921), .I2(n4507), .O(n4508) );
  NAND_GATE U5596 ( .I1(n4917), .I2(n4508), .O(n4937) );
  NAND_GATE U5597 ( .I1(n4935), .I2(n4942), .O(n4509) );
  NAND_GATE U5598 ( .I1(n4937), .I2(n4509), .O(n4510) );
  NAND_GATE U5599 ( .I1(n4933), .I2(n4510), .O(n4953) );
  NAND_GATE U5600 ( .I1(n4951), .I2(n4958), .O(n4511) );
  NAND_GATE U5601 ( .I1(n4953), .I2(n4511), .O(n4512) );
  NAND_GATE U5602 ( .I1(n4949), .I2(n4512), .O(n4969) );
  NAND_GATE U5603 ( .I1(n4967), .I2(n4974), .O(n4513) );
  NAND_GATE U5604 ( .I1(n4969), .I2(n4513), .O(n4514) );
  NAND_GATE U5605 ( .I1(n4965), .I2(n4514), .O(n4545) );
  NAND_GATE U5606 ( .I1(n4543), .I2(n4550), .O(n4515) );
  NAND_GATE U5607 ( .I1(n4545), .I2(n4515), .O(n4516) );
  NAND_GATE U5608 ( .I1(n4540), .I2(n4516), .O(n4530) );
  NAND_GATE U5609 ( .I1(n4528), .I2(n4535), .O(n4517) );
  NAND_GATE U5610 ( .I1(n4530), .I2(n4517), .O(n4519) );
  NAND_GATE U5611 ( .I1(n1435), .I2(A[31]), .O(n4518) );
  NAND3_GATE U5612 ( .I1(n4526), .I2(n4519), .I3(n4518), .O(n4523) );
  NAND_GATE U5613 ( .I1(n406), .I2(n4523), .O(n4525) );
  NAND_GATE U5614 ( .I1(n14793), .I2(n4525), .O(n4522) );
  INV_GATE U5615 ( .I1(n4525), .O(n14792) );
  NAND_GATE U5616 ( .I1(n4520), .I2(n14792), .O(n4521) );
  NAND_GATE U5617 ( .I1(n4522), .I2(n4521), .O(\A1[53] ) );
  NAND_GATE U5618 ( .I1(n4525), .I2(n4524), .O(n4984) );
  INV_GATE U5619 ( .I1(n4984), .O(n14795) );
  INV_GATE U5620 ( .I1(n4526), .O(n4527) );
  NAND_GATE U5621 ( .I1(n4527), .I2(n4530), .O(n4539) );
  NAND_GATE U5622 ( .I1(n4529), .I2(n4533), .O(n4537) );
  NAND_GATE U5623 ( .I1(n4531), .I2(n4530), .O(n4532) );
  NAND_GATE U5624 ( .I1(n4533), .I2(n4532), .O(n4534) );
  NAND_GATE U5625 ( .I1(n4535), .I2(n4534), .O(n4536) );
  NAND_GATE U5626 ( .I1(n4537), .I2(n4536), .O(n4538) );
  NAND_GATE U5627 ( .I1(n4539), .I2(n4538), .O(n4987) );
  NAND_GATE U5628 ( .I1(B[22]), .I2(A[30]), .O(n4999) );
  INV_GATE U5629 ( .I1(n4999), .O(n4981) );
  INV_GATE U5630 ( .I1(n4540), .O(n4541) );
  NAND_GATE U5631 ( .I1(n4541), .I2(n4545), .O(n4554) );
  INV_GATE U5632 ( .I1(n4545), .O(n4542) );
  NAND_GATE U5633 ( .I1(n4543), .I2(n4542), .O(n4548) );
  NAND_GATE U5634 ( .I1(n4544), .I2(n4548), .O(n4552) );
  NAND_GATE U5635 ( .I1(n4546), .I2(n4545), .O(n4547) );
  NAND_GATE U5636 ( .I1(n4548), .I2(n4547), .O(n4549) );
  NAND_GATE U5637 ( .I1(n4550), .I2(n4549), .O(n4551) );
  NAND_GATE U5638 ( .I1(n4552), .I2(n4551), .O(n4553) );
  NAND_GATE U5639 ( .I1(n4554), .I2(n4553), .O(n4997) );
  NAND_GATE U5640 ( .I1(n4981), .I2(n4997), .O(n4993) );
  NAND_GATE U5641 ( .I1(B[22]), .I2(A[29]), .O(n5010) );
  INV_GATE U5642 ( .I1(n5010), .O(n4979) );
  NAND_GATE U5643 ( .I1(B[22]), .I2(A[28]), .O(n5021) );
  INV_GATE U5644 ( .I1(n5021), .O(n4963) );
  NAND_GATE U5645 ( .I1(B[22]), .I2(A[27]), .O(n5032) );
  INV_GATE U5646 ( .I1(n5032), .O(n4947) );
  NAND_GATE U5647 ( .I1(B[22]), .I2(A[26]), .O(n5042) );
  INV_GATE U5648 ( .I1(n5042), .O(n4931) );
  NAND_GATE U5649 ( .I1(B[22]), .I2(A[25]), .O(n5052) );
  INV_GATE U5650 ( .I1(n5052), .O(n4915) );
  NAND_GATE U5651 ( .I1(B[22]), .I2(A[24]), .O(n5062) );
  INV_GATE U5652 ( .I1(n5062), .O(n4899) );
  NAND_GATE U5653 ( .I1(B[22]), .I2(A[23]), .O(n5073) );
  INV_GATE U5654 ( .I1(n5073), .O(n4883) );
  INV_GATE U5655 ( .I1(n4555), .O(n4556) );
  NAND_GATE U5656 ( .I1(n4556), .I2(n4559), .O(n4568) );
  NAND_GATE U5657 ( .I1(n4558), .I2(n4562), .O(n4566) );
  NAND_GATE U5658 ( .I1(n4560), .I2(n4559), .O(n4561) );
  NAND_GATE U5659 ( .I1(n4562), .I2(n4561), .O(n4563) );
  NAND_GATE U5660 ( .I1(n4564), .I2(n4563), .O(n4565) );
  NAND_GATE U5661 ( .I1(n4566), .I2(n4565), .O(n4567) );
  NAND_GATE U5662 ( .I1(n4568), .I2(n4567), .O(n5071) );
  NAND_GATE U5663 ( .I1(n4883), .I2(n5071), .O(n5068) );
  NAND_GATE U5664 ( .I1(B[22]), .I2(A[22]), .O(n5084) );
  INV_GATE U5665 ( .I1(n5084), .O(n4881) );
  NAND_GATE U5666 ( .I1(B[22]), .I2(A[21]), .O(n5377) );
  INV_GATE U5667 ( .I1(n5377), .O(n4865) );
  NAND_GATE U5668 ( .I1(B[22]), .I2(A[20]), .O(n5095) );
  INV_GATE U5669 ( .I1(n5095), .O(n4849) );
  NAND_GATE U5670 ( .I1(B[22]), .I2(A[19]), .O(n5106) );
  INV_GATE U5671 ( .I1(n5106), .O(n4833) );
  NAND_GATE U5672 ( .I1(B[22]), .I2(A[18]), .O(n5117) );
  INV_GATE U5673 ( .I1(n5117), .O(n4818) );
  NAND_GATE U5674 ( .I1(B[22]), .I2(A[17]), .O(n5122) );
  INV_GATE U5675 ( .I1(n5122), .O(n4803) );
  NAND_GATE U5676 ( .I1(B[22]), .I2(A[16]), .O(n5132) );
  INV_GATE U5677 ( .I1(n5132), .O(n4790) );
  NAND_GATE U5678 ( .I1(B[22]), .I2(A[15]), .O(n5143) );
  INV_GATE U5679 ( .I1(n5143), .O(n4775) );
  NAND_GATE U5680 ( .I1(n4572), .I2(n4571), .O(n4573) );
  NAND_GATE U5681 ( .I1(n4574), .I2(n4573), .O(n4579) );
  INV_GATE U5682 ( .I1(n4575), .O(n4577) );
  NAND_GATE U5683 ( .I1(n4577), .I2(n4576), .O(n4578) );
  NAND_GATE U5684 ( .I1(n4579), .I2(n4578), .O(n5144) );
  NAND_GATE U5685 ( .I1(n4775), .I2(n5144), .O(n5146) );
  NAND_GATE U5686 ( .I1(B[22]), .I2(A[14]), .O(n5153) );
  INV_GATE U5687 ( .I1(n5153), .O(n4773) );
  NAND_GATE U5688 ( .I1(B[22]), .I2(A[13]), .O(n5170) );
  INV_GATE U5689 ( .I1(n5170), .O(n4758) );
  NAND_GATE U5690 ( .I1(B[22]), .I2(A[12]), .O(n5180) );
  INV_GATE U5691 ( .I1(n5180), .O(n4739) );
  NAND_GATE U5692 ( .I1(B[22]), .I2(A[11]), .O(n5189) );
  INV_GATE U5693 ( .I1(n5189), .O(n4731) );
  NAND_GATE U5694 ( .I1(B[22]), .I2(A[10]), .O(n5467) );
  INV_GATE U5695 ( .I1(n5467), .O(n5345) );
  NAND_GATE U5696 ( .I1(n4580), .I2(n4436), .O(n4583) );
  NAND_GATE U5697 ( .I1(n4583), .I2(n4593), .O(n4587) );
  INV_GATE U5698 ( .I1(n4584), .O(n4585) );
  NAND3_GATE U5699 ( .I1(n4587), .I2(n4586), .I3(n4585), .O(n4590) );
  INV_GATE U5700 ( .I1(n4592), .O(n4595) );
  NAND4_GATE U5701 ( .I1(n4588), .I2(n4594), .I3(n4595), .I4(n4593), .O(n4589)
         );
  AND_GATE U5702 ( .I1(n4590), .I2(n4589), .O(n4600) );
  NAND_GATE U5703 ( .I1(n4594), .I2(n4593), .O(n4591) );
  NAND_GATE U5704 ( .I1(n4592), .I2(n4591), .O(n4598) );
  NAND3_GATE U5705 ( .I1(n4595), .I2(n4594), .I3(n4593), .O(n4597) );
  NAND3_GATE U5706 ( .I1(n4598), .I2(n4597), .I3(n4596), .O(n4599) );
  NAND_GATE U5707 ( .I1(n4600), .I2(n4599), .O(n5340) );
  NAND_GATE U5708 ( .I1(n5345), .I2(n5343), .O(n4717) );
  NAND_GATE U5709 ( .I1(B[22]), .I2(A[9]), .O(n5201) );
  INV_GATE U5710 ( .I1(n5201), .O(n5204) );
  NAND_GATE U5711 ( .I1(B[22]), .I2(A[8]), .O(n5324) );
  INV_GATE U5712 ( .I1(n5324), .O(n5325) );
  NAND_GATE U5713 ( .I1(n4609), .I2(n4608), .O(n4601) );
  INV_GATE U5714 ( .I1(n4611), .O(n4604) );
  NAND4_GATE U5715 ( .I1(n4606), .I2(n4605), .I3(n4604), .I4(n4601), .O(n5326)
         );
  NAND_GATE U5716 ( .I1(n4605), .I2(n4601), .O(n4610) );
  OR_GATE U5717 ( .I1(n4610), .I2(n4611), .O(n4613) );
  NAND_GATE U5718 ( .I1(n4611), .I2(n4610), .O(n4612) );
  NAND3_GATE U5719 ( .I1(n4614), .I2(n4613), .I3(n4612), .O(n5329) );
  NAND3_GATE U5720 ( .I1(n5327), .I2(n5326), .I3(n5329), .O(n5321) );
  NAND_GATE U5721 ( .I1(n5325), .I2(n881), .O(n4699) );
  NAND_GATE U5722 ( .I1(B[22]), .I2(A[7]), .O(n5306) );
  INV_GATE U5723 ( .I1(n5306), .O(n5310) );
  NAND_GATE U5724 ( .I1(B[22]), .I2(A[6]), .O(n5287) );
  INV_GATE U5725 ( .I1(n5287), .O(n5293) );
  INV_GATE U5726 ( .I1(n4624), .O(n4625) );
  NAND3_GATE U5727 ( .I1(n4625), .I2(n4617), .I3(n1217), .O(n4632) );
  NAND_GATE U5728 ( .I1(n4616), .I2(n4615), .O(n4617) );
  NAND_GATE U5729 ( .I1(n4618), .I2(n4617), .O(n4622) );
  INV_GATE U5730 ( .I1(n4619), .O(n4621) );
  NAND3_GATE U5731 ( .I1(n4622), .I2(n4621), .I3(n4620), .O(n4631) );
  NAND_GATE U5732 ( .I1(n4626), .I2(n4617), .O(n4623) );
  NAND_GATE U5733 ( .I1(n4624), .I2(n4623), .O(n4629) );
  NAND3_GATE U5734 ( .I1(n4626), .I2(n4617), .I3(n4625), .O(n4628) );
  NAND3_GATE U5735 ( .I1(n4629), .I2(n4628), .I3(n4627), .O(n4630) );
  NAND3_GATE U5736 ( .I1(n4632), .I2(n4631), .I3(n4630), .O(n5290) );
  NAND_GATE U5737 ( .I1(B[22]), .I2(A[5]), .O(n5280) );
  INV_GATE U5738 ( .I1(n5280), .O(n5281) );
  NAND_GATE U5739 ( .I1(B[22]), .I2(A[4]), .O(n5520) );
  INV_GATE U5740 ( .I1(n5520), .O(n5221) );
  NAND_GATE U5741 ( .I1(B[22]), .I2(A[3]), .O(n5232) );
  INV_GATE U5742 ( .I1(n5232), .O(n5223) );
  NAND_GATE U5743 ( .I1(B[22]), .I2(A[2]), .O(n5536) );
  INV_GATE U5744 ( .I1(n5536), .O(n5242) );
  NAND_GATE U5745 ( .I1(n1435), .I2(A[0]), .O(n4633) );
  NAND_GATE U5746 ( .I1(n14241), .I2(n4633), .O(n4634) );
  NAND_GATE U5747 ( .I1(B[24]), .I2(n4634), .O(n4637) );
  NAND_GATE U5748 ( .I1(n1436), .I2(A[1]), .O(n4635) );
  NAND_GATE U5749 ( .I1(n724), .I2(n4635), .O(n4636) );
  NAND_GATE U5750 ( .I1(B[23]), .I2(n4636), .O(n4638) );
  NAND_GATE U5751 ( .I1(n4637), .I2(n4638), .O(n5237) );
  NAND_GATE U5752 ( .I1(n5242), .I2(n5237), .O(n5243) );
  NAND3_GATE U5753 ( .I1(B[22]), .I2(B[23]), .I3(n1254), .O(n5240) );
  INV_GATE U5754 ( .I1(n5240), .O(n5244) );
  NAND_GATE U5755 ( .I1(n5536), .I2(n4638), .O(n4639) );
  NAND_GATE U5756 ( .I1(n5244), .I2(n4639), .O(n4640) );
  NAND_GATE U5757 ( .I1(n5243), .I2(n4640), .O(n5230) );
  NAND_GATE U5758 ( .I1(n5223), .I2(n5230), .O(n5224) );
  NAND3_GATE U5759 ( .I1(n4643), .I2(n4642), .I3(n4646), .O(n4644) );
  NAND_GATE U5760 ( .I1(n4645), .I2(n4644), .O(n4653) );
  NAND_GATE U5761 ( .I1(n4647), .I2(n4646), .O(n4648) );
  OR_GATE U5762 ( .I1(n4648), .I2(n4650), .O(n4652) );
  NAND_GATE U5763 ( .I1(n4650), .I2(n4649), .O(n4651) );
  NAND3_GATE U5764 ( .I1(n4653), .I2(n4652), .I3(n4651), .O(n5229) );
  NAND_GATE U5765 ( .I1(n5231), .I2(n5229), .O(n5227) );
  NAND_GATE U5766 ( .I1(n5230), .I2(n5227), .O(n4655) );
  NAND_GATE U5767 ( .I1(n5223), .I2(n5227), .O(n4654) );
  NAND3_GATE U5768 ( .I1(n5224), .I2(n4655), .I3(n4654), .O(n5220) );
  NAND_GATE U5769 ( .I1(n5221), .I2(n5220), .O(n4678) );
  NAND_GATE U5770 ( .I1(n4665), .I2(n4664), .O(n4658) );
  NAND_GATE U5771 ( .I1(n4673), .I2(n4658), .O(n4656) );
  NAND_GATE U5772 ( .I1(n4657), .I2(n4656), .O(n4661) );
  INV_GATE U5773 ( .I1(n4657), .O(n4672) );
  NAND3_GATE U5774 ( .I1(n4658), .I2(n4673), .I3(n4672), .O(n4660) );
  NAND3_GATE U5775 ( .I1(n4661), .I2(n4660), .I3(n4659), .O(n5214) );
  NAND_GATE U5776 ( .I1(n4663), .I2(n4662), .O(n4666) );
  NAND_GATE U5777 ( .I1(n4666), .I2(n4658), .O(n4670) );
  INV_GATE U5778 ( .I1(n4667), .O(n4668) );
  NAND3_GATE U5779 ( .I1(n4670), .I2(n4669), .I3(n4668), .O(n4674) );
  NAND4_GATE U5780 ( .I1(n4673), .I2(n4672), .I3(n4671), .I4(n4658), .O(n4675)
         );
  NAND3_GATE U5781 ( .I1(n5214), .I2(n1296), .I3(n5221), .O(n4677) );
  NAND4_GATE U5782 ( .I1(n4675), .I2(n5214), .I3(n5220), .I4(n4674), .O(n4676)
         );
  NAND3_GATE U5783 ( .I1(n4678), .I2(n4677), .I3(n4676), .O(n5277) );
  NAND_GATE U5784 ( .I1(n5281), .I2(n5277), .O(n5283) );
  NAND3_GATE U5785 ( .I1(n5270), .I2(n5261), .I3(n676), .O(n5267) );
  NAND_GATE U5786 ( .I1(n5270), .I2(n676), .O(n4681) );
  INV_GATE U5787 ( .I1(n5270), .O(n5269) );
  NAND3_GATE U5788 ( .I1(n5273), .I2(n5268), .I3(n5269), .O(n4680) );
  NAND_GATE U5789 ( .I1(n5261), .I2(n5271), .O(n4679) );
  NAND3_GATE U5790 ( .I1(n4681), .I2(n4680), .I3(n4679), .O(n4682) );
  NAND_GATE U5791 ( .I1(n5267), .I2(n4682), .O(n5284) );
  NAND_GATE U5792 ( .I1(n5277), .I2(n5284), .O(n4684) );
  NAND_GATE U5793 ( .I1(n5281), .I2(n5284), .O(n4683) );
  NAND3_GATE U5794 ( .I1(n5283), .I2(n4684), .I3(n4683), .O(n5288) );
  NAND_GATE U5795 ( .I1(n5287), .I2(n5290), .O(n4685) );
  NAND_GATE U5796 ( .I1(n5288), .I2(n4685), .O(n4686) );
  NAND_GATE U5797 ( .I1(n5310), .I2(n758), .O(n5311) );
  NAND3_GATE U5798 ( .I1(n4687), .I2(n728), .I3(n4688), .O(n5303) );
  AND_GATE U5799 ( .I1(n5303), .I2(n5301), .O(n4693) );
  NAND_GATE U5800 ( .I1(n4688), .I2(n728), .O(n4694) );
  NAND_GATE U5801 ( .I1(n5298), .I2(n4689), .O(n5302) );
  INV_GATE U5802 ( .I1(n5302), .O(n4690) );
  NAND_GATE U5803 ( .I1(n4691), .I2(n4690), .O(n5305) );
  NAND3_GATE U5804 ( .I1(n5298), .I2(n4694), .I3(n5305), .O(n4692) );
  NAND3_GATE U5805 ( .I1(n758), .I2(n4693), .I3(n4692), .O(n4696) );
  NAND3_GATE U5806 ( .I1(n5298), .I2(n5305), .I3(n4694), .O(n5309) );
  NAND3_GATE U5807 ( .I1(n5310), .I2(n4693), .I3(n5309), .O(n4695) );
  NAND3_GATE U5808 ( .I1(n5311), .I2(n4696), .I3(n4695), .O(n5323) );
  NAND_GATE U5809 ( .I1(n5324), .I2(n5321), .O(n4697) );
  NAND_GATE U5810 ( .I1(n5323), .I2(n4697), .O(n4698) );
  NAND_GATE U5811 ( .I1(n4699), .I2(n4698), .O(n5198) );
  NAND_GATE U5812 ( .I1(n5204), .I2(n5198), .O(n5209) );
  NAND4_GATE U5813 ( .I1(n4702), .I2(n4701), .I3(n4709), .I4(n4700), .O(n4703)
         );
  NAND3_GATE U5814 ( .I1(n5202), .I2(n4705), .I3(n1301), .O(n4708) );
  INV_GATE U5815 ( .I1(n4705), .O(n5203) );
  NAND4_GATE U5816 ( .I1(n4704), .I2(n4703), .I3(n4708), .I4(n4707), .O(n4706)
         );
  NAND_GATE U5817 ( .I1(n1301), .I2(n1221), .O(n4710) );
  NAND_GATE U5818 ( .I1(n4706), .I2(n4710), .O(n5210) );
  NAND_GATE U5819 ( .I1(n5198), .I2(n5210), .O(n4714) );
  NAND_GATE U5820 ( .I1(n5203), .I2(n387), .O(n4711) );
  NAND3_GATE U5821 ( .I1(n4711), .I2(n4710), .I3(n4709), .O(n4712) );
  NAND3_GATE U5822 ( .I1(n5204), .I2(n1223), .I3(n4712), .O(n4713) );
  NAND3_GATE U5823 ( .I1(n5209), .I2(n4714), .I3(n4713), .O(n5344) );
  NAND_GATE U5824 ( .I1(n5467), .I2(n5340), .O(n4715) );
  NAND_GATE U5825 ( .I1(n5344), .I2(n4715), .O(n4716) );
  NAND_GATE U5826 ( .I1(n4717), .I2(n4716), .O(n5188) );
  NAND_GATE U5827 ( .I1(n4731), .I2(n5188), .O(n5193) );
  NAND3_GATE U5828 ( .I1(n4727), .I2(n4719), .I3(n4718), .O(n4728) );
  INV_GATE U5829 ( .I1(n4719), .O(n4721) );
  NAND_GATE U5830 ( .I1(n4722), .I2(n4721), .O(n4729) );
  NAND_GATE U5831 ( .I1(n4727), .I2(n4729), .O(n4723) );
  NAND3_GATE U5832 ( .I1(n4722), .I2(n4721), .I3(n4720), .O(n4725) );
  NAND3_GATE U5833 ( .I1(n4726), .I2(n4723), .I3(n4725), .O(n4724) );
  NAND_GATE U5834 ( .I1(n4728), .I2(n4724), .O(n5194) );
  NAND_GATE U5835 ( .I1(n5188), .I2(n5194), .O(n4733) );
  NAND3_GATE U5836 ( .I1(n4729), .I2(n4728), .I3(n4727), .O(n4730) );
  AND_GATE U5837 ( .I1(n4731), .I2(n4730), .O(n5192) );
  NAND_GATE U5838 ( .I1(n1222), .I2(n5192), .O(n4732) );
  NAND3_GATE U5839 ( .I1(n5193), .I2(n4733), .I3(n4732), .O(n5181) );
  NAND_GATE U5840 ( .I1(n4739), .I2(n5181), .O(n5183) );
  NAND_GATE U5841 ( .I1(n1303), .I2(n4736), .O(n4735) );
  NAND_GATE U5842 ( .I1(n4735), .I2(n4734), .O(n5173) );
  NAND3_GATE U5843 ( .I1(n308), .I2(n4738), .I3(n4737), .O(n4742) );
  NAND_GATE U5844 ( .I1(n730), .I2(n4742), .O(n5176) );
  NAND3_GATE U5845 ( .I1(n5175), .I2(n5176), .I3(n4739), .O(n5182) );
  NAND_GATE U5846 ( .I1(n4740), .I2(n5175), .O(n4741) );
  NAND_GATE U5847 ( .I1(n4742), .I2(n4741), .O(n5184) );
  NAND_GATE U5848 ( .I1(n5181), .I2(n5184), .O(n4743) );
  NAND3_GATE U5849 ( .I1(n5183), .I2(n5182), .I3(n4743), .O(n5167) );
  NAND_GATE U5850 ( .I1(n4758), .I2(n5167), .O(n5162) );
  NAND_GATE U5851 ( .I1(n4746), .I2(n311), .O(n4744) );
  NAND_GATE U5852 ( .I1(n4745), .I2(n4744), .O(n4752) );
  NAND_GATE U5853 ( .I1(n810), .I2(n4754), .O(n4747) );
  NAND_GATE U5854 ( .I1(n4748), .I2(n4747), .O(n4749) );
  NAND_GATE U5855 ( .I1(n4750), .I2(n4749), .O(n4751) );
  NAND_GATE U5856 ( .I1(n4752), .I2(n4751), .O(n4757) );
  INV_GATE U5857 ( .I1(n4753), .O(n4755) );
  NAND_GATE U5858 ( .I1(n4755), .I2(n4754), .O(n4756) );
  NAND_GATE U5859 ( .I1(n4757), .I2(n4756), .O(n5166) );
  NAND_GATE U5860 ( .I1(n5167), .I2(n5166), .O(n4759) );
  NAND3_GATE U5861 ( .I1(n5162), .I2(n5161), .I3(n4759), .O(n5154) );
  NAND_GATE U5862 ( .I1(n4773), .I2(n5154), .O(n5156) );
  NAND_GATE U5863 ( .I1(n4761), .I2(n4760), .O(n4767) );
  NAND_GATE U5864 ( .I1(n905), .I2(n4769), .O(n4763) );
  NAND_GATE U5865 ( .I1(n4763), .I2(n4760), .O(n4764) );
  NAND_GATE U5866 ( .I1(n4765), .I2(n4764), .O(n4766) );
  NAND_GATE U5867 ( .I1(n4767), .I2(n4766), .O(n4772) );
  INV_GATE U5868 ( .I1(n4768), .O(n4770) );
  NAND_GATE U5869 ( .I1(n4770), .I2(n4769), .O(n4771) );
  NAND_GATE U5870 ( .I1(n4772), .I2(n4771), .O(n5157) );
  NAND_GATE U5871 ( .I1(n4773), .I2(n5157), .O(n5155) );
  NAND_GATE U5872 ( .I1(n5154), .I2(n5157), .O(n4774) );
  NAND_GATE U5873 ( .I1(n5144), .I2(n5147), .O(n4776) );
  NAND_GATE U5874 ( .I1(n4790), .I2(n893), .O(n5136) );
  INV_GATE U5875 ( .I1(n4777), .O(n4778) );
  NAND_GATE U5876 ( .I1(n4778), .I2(n4780), .O(n4789) );
  NAND_GATE U5877 ( .I1(n4779), .I2(n4782), .O(n4787) );
  NAND_GATE U5878 ( .I1(n4781), .I2(n1349), .O(n4782) );
  NAND_GATE U5879 ( .I1(n4783), .I2(n4782), .O(n4784) );
  NAND_GATE U5880 ( .I1(n4785), .I2(n4784), .O(n4786) );
  NAND_GATE U5881 ( .I1(n4787), .I2(n4786), .O(n4788) );
  NAND_GATE U5882 ( .I1(n4789), .I2(n4788), .O(n5137) );
  NAND_GATE U5883 ( .I1(n4790), .I2(n5137), .O(n5135) );
  NAND_GATE U5884 ( .I1(n893), .I2(n5137), .O(n4791) );
  NAND3_GATE U5885 ( .I1(n5136), .I2(n5135), .I3(n4791), .O(n5125) );
  NAND_GATE U5886 ( .I1(n4803), .I2(n5125), .O(n5127) );
  NAND_GATE U5887 ( .I1(n220), .I2(n4795), .O(n4802) );
  INV_GATE U5888 ( .I1(n4795), .O(n4796) );
  NAND_GATE U5889 ( .I1(n4797), .I2(n4796), .O(n4793) );
  NAND_GATE U5890 ( .I1(n4794), .I2(n4793), .O(n4801) );
  NAND_GATE U5891 ( .I1(n4798), .I2(n4793), .O(n4799) );
  NAND_GATE U5892 ( .I1(n4803), .I2(n5128), .O(n5126) );
  NAND_GATE U5893 ( .I1(n5125), .I2(n5128), .O(n4804) );
  NAND3_GATE U5894 ( .I1(n5127), .I2(n5126), .I3(n4804), .O(n5116) );
  NAND_GATE U5895 ( .I1(n4818), .I2(n5116), .O(n5112) );
  INV_GATE U5896 ( .I1(n4805), .O(n4806) );
  NAND_GATE U5897 ( .I1(n4806), .I2(n4809), .O(n4817) );
  NAND_GATE U5898 ( .I1(n4808), .I2(n4811), .O(n4815) );
  NAND_GATE U5899 ( .I1(n313), .I2(n4809), .O(n4810) );
  NAND_GATE U5900 ( .I1(n4811), .I2(n4810), .O(n4812) );
  NAND_GATE U5901 ( .I1(n4813), .I2(n4812), .O(n4814) );
  NAND_GATE U5902 ( .I1(n4815), .I2(n4814), .O(n4816) );
  NAND_GATE U5903 ( .I1(n4817), .I2(n4816), .O(n5115) );
  NAND_GATE U5904 ( .I1(n5116), .I2(n5115), .O(n4819) );
  NAND3_GATE U5905 ( .I1(n5112), .I2(n5111), .I3(n4819), .O(n5105) );
  NAND_GATE U5906 ( .I1(n4833), .I2(n5105), .O(n5101) );
  INV_GATE U5907 ( .I1(n4820), .O(n4821) );
  NAND_GATE U5908 ( .I1(n4821), .I2(n4824), .O(n4832) );
  NAND_GATE U5909 ( .I1(n4823), .I2(n4826), .O(n4830) );
  NAND_GATE U5910 ( .I1(n801), .I2(n4824), .O(n4825) );
  NAND_GATE U5911 ( .I1(n4826), .I2(n4825), .O(n4827) );
  NAND_GATE U5912 ( .I1(n4828), .I2(n4827), .O(n4829) );
  NAND_GATE U5913 ( .I1(n4830), .I2(n4829), .O(n4831) );
  NAND_GATE U5914 ( .I1(n4832), .I2(n4831), .O(n5104) );
  NAND_GATE U5915 ( .I1(n4833), .I2(n5104), .O(n5100) );
  NAND_GATE U5916 ( .I1(n5105), .I2(n5104), .O(n4834) );
  NAND3_GATE U5917 ( .I1(n5101), .I2(n5100), .I3(n4834), .O(n5094) );
  NAND_GATE U5918 ( .I1(n4849), .I2(n5094), .O(n5090) );
  INV_GATE U5919 ( .I1(n4835), .O(n4836) );
  NAND_GATE U5920 ( .I1(n4836), .I2(n4839), .O(n4848) );
  NAND_GATE U5921 ( .I1(n4838), .I2(n4842), .O(n4846) );
  NAND_GATE U5922 ( .I1(n4840), .I2(n4839), .O(n4841) );
  NAND_GATE U5923 ( .I1(n4842), .I2(n4841), .O(n4843) );
  NAND_GATE U5924 ( .I1(n4844), .I2(n4843), .O(n4845) );
  NAND_GATE U5925 ( .I1(n4846), .I2(n4845), .O(n4847) );
  NAND_GATE U5926 ( .I1(n4848), .I2(n4847), .O(n5093) );
  NAND_GATE U5927 ( .I1(n5094), .I2(n5093), .O(n4850) );
  NAND3_GATE U5928 ( .I1(n5090), .I2(n5089), .I3(n4850), .O(n5376) );
  NAND_GATE U5929 ( .I1(n4865), .I2(n5376), .O(n5372) );
  INV_GATE U5930 ( .I1(n4851), .O(n4852) );
  NAND_GATE U5931 ( .I1(n4852), .I2(n4855), .O(n4864) );
  NAND_GATE U5932 ( .I1(n4854), .I2(n4858), .O(n4862) );
  NAND_GATE U5933 ( .I1(n4856), .I2(n4855), .O(n4857) );
  NAND_GATE U5934 ( .I1(n4858), .I2(n4857), .O(n4859) );
  NAND_GATE U5935 ( .I1(n4860), .I2(n4859), .O(n4861) );
  NAND_GATE U5936 ( .I1(n4862), .I2(n4861), .O(n4863) );
  NAND_GATE U5937 ( .I1(n4864), .I2(n4863), .O(n5375) );
  NAND_GATE U5938 ( .I1(n4865), .I2(n5375), .O(n5371) );
  NAND_GATE U5939 ( .I1(n5376), .I2(n5375), .O(n4866) );
  NAND3_GATE U5940 ( .I1(n5372), .I2(n5371), .I3(n4866), .O(n5083) );
  NAND_GATE U5941 ( .I1(n4881), .I2(n5083), .O(n5079) );
  INV_GATE U5942 ( .I1(n4867), .O(n4868) );
  NAND_GATE U5943 ( .I1(n4868), .I2(n4871), .O(n4880) );
  NAND_GATE U5944 ( .I1(n4870), .I2(n4874), .O(n4878) );
  NAND_GATE U5945 ( .I1(n4872), .I2(n4871), .O(n4873) );
  NAND_GATE U5946 ( .I1(n4874), .I2(n4873), .O(n4875) );
  NAND_GATE U5947 ( .I1(n4876), .I2(n4875), .O(n4877) );
  NAND_GATE U5948 ( .I1(n4878), .I2(n4877), .O(n4879) );
  NAND_GATE U5949 ( .I1(n4880), .I2(n4879), .O(n5082) );
  NAND_GATE U5950 ( .I1(n4881), .I2(n5082), .O(n5078) );
  NAND_GATE U5951 ( .I1(n5083), .I2(n5082), .O(n4882) );
  NAND3_GATE U5952 ( .I1(n5079), .I2(n5078), .I3(n4882), .O(n5072) );
  NAND_GATE U5953 ( .I1(n4883), .I2(n5072), .O(n5067) );
  NAND_GATE U5954 ( .I1(n5071), .I2(n5072), .O(n4884) );
  NAND3_GATE U5955 ( .I1(n5068), .I2(n5067), .I3(n4884), .O(n5061) );
  NAND_GATE U5956 ( .I1(n4899), .I2(n5061), .O(n5057) );
  INV_GATE U5957 ( .I1(n4885), .O(n4886) );
  NAND_GATE U5958 ( .I1(n4886), .I2(n4889), .O(n4898) );
  NAND_GATE U5959 ( .I1(n4888), .I2(n4892), .O(n4896) );
  NAND_GATE U5960 ( .I1(n4890), .I2(n4889), .O(n4891) );
  NAND_GATE U5961 ( .I1(n4892), .I2(n4891), .O(n4893) );
  NAND_GATE U5962 ( .I1(n4894), .I2(n4893), .O(n4895) );
  NAND_GATE U5963 ( .I1(n4896), .I2(n4895), .O(n4897) );
  NAND_GATE U5964 ( .I1(n4898), .I2(n4897), .O(n5060) );
  NAND_GATE U5965 ( .I1(n4899), .I2(n5060), .O(n5056) );
  NAND_GATE U5966 ( .I1(n5061), .I2(n5060), .O(n4900) );
  NAND3_GATE U5967 ( .I1(n5057), .I2(n5056), .I3(n4900), .O(n5051) );
  NAND_GATE U5968 ( .I1(n4915), .I2(n5051), .O(n5047) );
  OR_GATE U5969 ( .I1(n4902), .I2(n4901), .O(n4914) );
  NAND_GATE U5970 ( .I1(n4903), .I2(n4902), .O(n4908) );
  NAND_GATE U5971 ( .I1(n4904), .I2(n4908), .O(n4912) );
  NAND_GATE U5972 ( .I1(n4906), .I2(n4905), .O(n4907) );
  NAND_GATE U5973 ( .I1(n4908), .I2(n4907), .O(n4909) );
  NAND_GATE U5974 ( .I1(n4910), .I2(n4909), .O(n4911) );
  NAND_GATE U5975 ( .I1(n4912), .I2(n4911), .O(n4913) );
  NAND_GATE U5976 ( .I1(n4914), .I2(n4913), .O(n5050) );
  NAND_GATE U5977 ( .I1(n4915), .I2(n5050), .O(n5046) );
  NAND_GATE U5978 ( .I1(n5051), .I2(n5050), .O(n4916) );
  NAND3_GATE U5979 ( .I1(n5047), .I2(n5046), .I3(n4916), .O(n5041) );
  NAND_GATE U5980 ( .I1(n4931), .I2(n5041), .O(n5037) );
  INV_GATE U5981 ( .I1(n4917), .O(n4918) );
  NAND_GATE U5982 ( .I1(n4918), .I2(n4921), .O(n4930) );
  NAND_GATE U5983 ( .I1(n4920), .I2(n4924), .O(n4928) );
  NAND_GATE U5984 ( .I1(n4922), .I2(n4921), .O(n4923) );
  NAND_GATE U5985 ( .I1(n4924), .I2(n4923), .O(n4925) );
  NAND_GATE U5986 ( .I1(n4926), .I2(n4925), .O(n4927) );
  NAND_GATE U5987 ( .I1(n4928), .I2(n4927), .O(n4929) );
  NAND_GATE U5988 ( .I1(n4930), .I2(n4929), .O(n5040) );
  NAND_GATE U5989 ( .I1(n4931), .I2(n5040), .O(n5036) );
  NAND_GATE U5990 ( .I1(n5041), .I2(n5040), .O(n4932) );
  NAND3_GATE U5991 ( .I1(n5037), .I2(n5036), .I3(n4932), .O(n5031) );
  NAND_GATE U5992 ( .I1(n4947), .I2(n5031), .O(n5027) );
  INV_GATE U5993 ( .I1(n4933), .O(n4934) );
  NAND_GATE U5994 ( .I1(n4934), .I2(n4937), .O(n4946) );
  NAND_GATE U5995 ( .I1(n4936), .I2(n4940), .O(n4944) );
  NAND_GATE U5996 ( .I1(n4938), .I2(n4937), .O(n4939) );
  NAND_GATE U5997 ( .I1(n4940), .I2(n4939), .O(n4941) );
  NAND_GATE U5998 ( .I1(n4942), .I2(n4941), .O(n4943) );
  NAND_GATE U5999 ( .I1(n4944), .I2(n4943), .O(n4945) );
  NAND_GATE U6000 ( .I1(n4946), .I2(n4945), .O(n5030) );
  NAND_GATE U6001 ( .I1(n4947), .I2(n5030), .O(n5026) );
  NAND_GATE U6002 ( .I1(n5031), .I2(n5030), .O(n4948) );
  NAND3_GATE U6003 ( .I1(n5027), .I2(n5026), .I3(n4948), .O(n5020) );
  NAND_GATE U6004 ( .I1(n4963), .I2(n5020), .O(n5016) );
  INV_GATE U6005 ( .I1(n4949), .O(n4950) );
  NAND_GATE U6006 ( .I1(n4950), .I2(n4953), .O(n4962) );
  NAND_GATE U6007 ( .I1(n4952), .I2(n4956), .O(n4960) );
  NAND_GATE U6008 ( .I1(n4954), .I2(n4953), .O(n4955) );
  NAND_GATE U6009 ( .I1(n4956), .I2(n4955), .O(n4957) );
  NAND_GATE U6010 ( .I1(n4958), .I2(n4957), .O(n4959) );
  NAND_GATE U6011 ( .I1(n4960), .I2(n4959), .O(n4961) );
  NAND_GATE U6012 ( .I1(n4962), .I2(n4961), .O(n5019) );
  NAND_GATE U6013 ( .I1(n4963), .I2(n5019), .O(n5015) );
  NAND_GATE U6014 ( .I1(n5020), .I2(n5019), .O(n4964) );
  NAND3_GATE U6015 ( .I1(n5016), .I2(n5015), .I3(n4964), .O(n5009) );
  NAND_GATE U6016 ( .I1(n4979), .I2(n5009), .O(n5005) );
  INV_GATE U6017 ( .I1(n4965), .O(n4966) );
  NAND_GATE U6018 ( .I1(n4966), .I2(n4969), .O(n4978) );
  NAND_GATE U6019 ( .I1(n4968), .I2(n4972), .O(n4976) );
  NAND_GATE U6020 ( .I1(n4970), .I2(n4969), .O(n4971) );
  NAND_GATE U6021 ( .I1(n4972), .I2(n4971), .O(n4973) );
  NAND_GATE U6022 ( .I1(n4974), .I2(n4973), .O(n4975) );
  NAND_GATE U6023 ( .I1(n4976), .I2(n4975), .O(n4977) );
  NAND_GATE U6024 ( .I1(n4978), .I2(n4977), .O(n5008) );
  NAND_GATE U6025 ( .I1(n4979), .I2(n5008), .O(n5004) );
  NAND_GATE U6026 ( .I1(n5009), .I2(n5008), .O(n4980) );
  NAND3_GATE U6027 ( .I1(n5005), .I2(n5004), .I3(n4980), .O(n4998) );
  NAND_GATE U6028 ( .I1(n4998), .I2(n4997), .O(n4982) );
  NAND_GATE U6029 ( .I1(n4981), .I2(n4998), .O(n4994) );
  AND3_GATE U6030 ( .I1(n4993), .I2(n4982), .I3(n4994), .O(n4989) );
  NAND_GATE U6031 ( .I1(n1434), .I2(A[31]), .O(n4988) );
  NAND_GATE U6032 ( .I1(n4989), .I2(n4988), .O(n4983) );
  NAND_GATE U6033 ( .I1(n4987), .I2(n4983), .O(n4992) );
  NAND_GATE U6034 ( .I1(n14795), .I2(n4992), .O(n4986) );
  INV_GATE U6035 ( .I1(n4992), .O(n14794) );
  NAND_GATE U6036 ( .I1(n4984), .I2(n14794), .O(n4985) );
  NAND_GATE U6037 ( .I1(n4986), .I2(n4985), .O(\A1[52] ) );
  INV_GATE U6038 ( .I1(n4987), .O(n4990) );
  NAND3_GATE U6039 ( .I1(n4990), .I2(n4989), .I3(n4988), .O(n4991) );
  NAND_GATE U6040 ( .I1(n4992), .I2(n4991), .O(n5401) );
  INV_GATE U6041 ( .I1(n5401), .O(n14797) );
  OR_GATE U6042 ( .I1(n4993), .I2(n4998), .O(n4996) );
  OR_GATE U6043 ( .I1(n4997), .I2(n4994), .O(n4995) );
  AND_GATE U6044 ( .I1(n4996), .I2(n4995), .O(n5003) );
  NAND_GATE U6045 ( .I1(n1190), .I2(n4997), .O(n5001) );
  NAND3_GATE U6046 ( .I1(n5001), .I2(n5000), .I3(n4999), .O(n5002) );
  NAND_GATE U6047 ( .I1(n5003), .I2(n5002), .O(n5404) );
  OR_GATE U6048 ( .I1(n5004), .I2(n5009), .O(n5007) );
  OR_GATE U6049 ( .I1(n5008), .I2(n5005), .O(n5006) );
  AND_GATE U6050 ( .I1(n5007), .I2(n5006), .O(n5014) );
  NAND_GATE U6051 ( .I1(n5009), .I2(n1181), .O(n5011) );
  NAND3_GATE U6052 ( .I1(n5012), .I2(n5011), .I3(n5010), .O(n5013) );
  NAND_GATE U6053 ( .I1(n5014), .I2(n5013), .O(n5409) );
  INV_GATE U6054 ( .I1(n5409), .O(n5412) );
  NAND_GATE U6055 ( .I1(B[21]), .I2(A[30]), .O(n5416) );
  INV_GATE U6056 ( .I1(n5416), .O(n5410) );
  NAND_GATE U6057 ( .I1(n5412), .I2(n5410), .O(n5407) );
  OR_GATE U6058 ( .I1(n5015), .I2(n5020), .O(n5018) );
  OR_GATE U6059 ( .I1(n5019), .I2(n5016), .O(n5017) );
  AND_GATE U6060 ( .I1(n5018), .I2(n5017), .O(n5025) );
  NAND_GATE U6061 ( .I1(n5020), .I2(n1174), .O(n5022) );
  NAND3_GATE U6062 ( .I1(n5023), .I2(n5022), .I3(n5021), .O(n5024) );
  NAND_GATE U6063 ( .I1(n5025), .I2(n5024), .O(n5423) );
  INV_GATE U6064 ( .I1(n5423), .O(n5426) );
  NAND_GATE U6065 ( .I1(B[21]), .I2(A[29]), .O(n5430) );
  INV_GATE U6066 ( .I1(n5430), .O(n5424) );
  NAND_GATE U6067 ( .I1(n5426), .I2(n5424), .O(n5421) );
  OR_GATE U6068 ( .I1(n5026), .I2(n5031), .O(n5029) );
  OR_GATE U6069 ( .I1(n5030), .I2(n5027), .O(n5028) );
  NAND_GATE U6070 ( .I1(n5031), .I2(n1169), .O(n5033) );
  NAND3_GATE U6071 ( .I1(n5034), .I2(n5033), .I3(n5032), .O(n5035) );
  INV_GATE U6072 ( .I1(n5813), .O(n5816) );
  NAND_GATE U6073 ( .I1(B[21]), .I2(A[28]), .O(n5820) );
  INV_GATE U6074 ( .I1(n5820), .O(n5814) );
  NAND_GATE U6075 ( .I1(n5816), .I2(n5814), .O(n5811) );
  OR_GATE U6076 ( .I1(n5036), .I2(n5041), .O(n5039) );
  OR_GATE U6077 ( .I1(n5040), .I2(n5037), .O(n5038) );
  NAND_GATE U6078 ( .I1(n1122), .I2(n5040), .O(n5044) );
  NAND3_GATE U6079 ( .I1(n5044), .I2(n5043), .I3(n5042), .O(n5045) );
  INV_GATE U6080 ( .I1(n5797), .O(n5800) );
  NAND_GATE U6081 ( .I1(B[21]), .I2(A[27]), .O(n5804) );
  INV_GATE U6082 ( .I1(n5804), .O(n5798) );
  NAND_GATE U6083 ( .I1(n5800), .I2(n5798), .O(n5794) );
  OR_GATE U6084 ( .I1(n5046), .I2(n5051), .O(n5049) );
  OR_GATE U6085 ( .I1(n5050), .I2(n5047), .O(n5048) );
  NAND_GATE U6086 ( .I1(n1146), .I2(n5050), .O(n5054) );
  NAND3_GATE U6087 ( .I1(n5054), .I2(n5053), .I3(n5052), .O(n5055) );
  INV_GATE U6088 ( .I1(n5780), .O(n5783) );
  NAND_GATE U6089 ( .I1(B[21]), .I2(A[26]), .O(n5787) );
  INV_GATE U6090 ( .I1(n5787), .O(n5781) );
  NAND_GATE U6091 ( .I1(n5783), .I2(n5781), .O(n5778) );
  OR_GATE U6092 ( .I1(n5056), .I2(n5061), .O(n5059) );
  OR_GATE U6093 ( .I1(n5060), .I2(n5057), .O(n5058) );
  AND_GATE U6094 ( .I1(n5059), .I2(n5058), .O(n5066) );
  NAND_GATE U6095 ( .I1(n1145), .I2(n5060), .O(n5064) );
  NAND3_GATE U6096 ( .I1(n5064), .I2(n5063), .I3(n5062), .O(n5065) );
  NAND_GATE U6097 ( .I1(n5066), .I2(n5065), .O(n5764) );
  INV_GATE U6098 ( .I1(n5764), .O(n5767) );
  NAND_GATE U6099 ( .I1(B[21]), .I2(A[25]), .O(n5771) );
  INV_GATE U6100 ( .I1(n5771), .O(n5765) );
  NAND_GATE U6101 ( .I1(n5767), .I2(n5765), .O(n5762) );
  OR_GATE U6102 ( .I1(n5067), .I2(n5071), .O(n5070) );
  OR_GATE U6103 ( .I1(n5072), .I2(n5068), .O(n5069) );
  AND_GATE U6104 ( .I1(n5070), .I2(n5069), .O(n5077) );
  NAND_GATE U6105 ( .I1(n5071), .I2(n1161), .O(n5075) );
  NAND3_GATE U6106 ( .I1(n5075), .I2(n5074), .I3(n5073), .O(n5076) );
  NAND_GATE U6107 ( .I1(n5077), .I2(n5076), .O(n5748) );
  INV_GATE U6108 ( .I1(n5748), .O(n5751) );
  NAND_GATE U6109 ( .I1(B[21]), .I2(A[24]), .O(n5755) );
  INV_GATE U6110 ( .I1(n5755), .O(n5749) );
  NAND_GATE U6111 ( .I1(n5751), .I2(n5749), .O(n5746) );
  OR_GATE U6112 ( .I1(n5078), .I2(n5083), .O(n5081) );
  OR_GATE U6113 ( .I1(n5082), .I2(n5079), .O(n5080) );
  AND_GATE U6114 ( .I1(n5081), .I2(n5080), .O(n5088) );
  NAND_GATE U6115 ( .I1(n1160), .I2(n5082), .O(n5086) );
  NAND3_GATE U6116 ( .I1(n5086), .I2(n5085), .I3(n5084), .O(n5087) );
  NAND_GATE U6117 ( .I1(n5088), .I2(n5087), .O(n5732) );
  INV_GATE U6118 ( .I1(n5732), .O(n5735) );
  NAND_GATE U6119 ( .I1(B[21]), .I2(A[23]), .O(n5739) );
  INV_GATE U6120 ( .I1(n5739), .O(n5733) );
  NAND_GATE U6121 ( .I1(n5735), .I2(n5733), .O(n5730) );
  NAND_GATE U6122 ( .I1(B[21]), .I2(A[22]), .O(n5723) );
  INV_GATE U6123 ( .I1(n5723), .O(n5717) );
  OR_GATE U6124 ( .I1(n5089), .I2(n5094), .O(n5092) );
  OR_GATE U6125 ( .I1(n5093), .I2(n5090), .O(n5091) );
  AND_GATE U6126 ( .I1(n5092), .I2(n5091), .O(n5099) );
  NAND_GATE U6127 ( .I1(n1117), .I2(n5093), .O(n5097) );
  NAND3_GATE U6128 ( .I1(n5097), .I2(n5096), .I3(n5095), .O(n5098) );
  NAND_GATE U6129 ( .I1(B[21]), .I2(A[21]), .O(n5708) );
  INV_GATE U6130 ( .I1(n5708), .O(n5703) );
  NAND_GATE U6131 ( .I1(n800), .I2(n5703), .O(n5701) );
  OR_GATE U6132 ( .I1(n5100), .I2(n5105), .O(n5103) );
  OR_GATE U6133 ( .I1(n5104), .I2(n5101), .O(n5102) );
  AND_GATE U6134 ( .I1(n5103), .I2(n5102), .O(n5110) );
  NAND_GATE U6135 ( .I1(n1119), .I2(n5104), .O(n5108) );
  NAND3_GATE U6136 ( .I1(n5108), .I2(n5107), .I3(n5106), .O(n5109) );
  NAND_GATE U6137 ( .I1(B[21]), .I2(A[20]), .O(n5443) );
  INV_GATE U6138 ( .I1(n5443), .O(n5438) );
  NAND_GATE U6139 ( .I1(n798), .I2(n5438), .O(n5435) );
  OR_GATE U6140 ( .I1(n5111), .I2(n5116), .O(n5114) );
  OR_GATE U6141 ( .I1(n5115), .I2(n5112), .O(n5113) );
  AND_GATE U6142 ( .I1(n5114), .I2(n5113), .O(n5121) );
  NAND_GATE U6143 ( .I1(n1120), .I2(n5115), .O(n5119) );
  NAND3_GATE U6144 ( .I1(n5119), .I2(n5118), .I3(n5117), .O(n5120) );
  NAND_GATE U6145 ( .I1(n5121), .I2(n5120), .O(n5686) );
  NAND_GATE U6146 ( .I1(B[21]), .I2(A[19]), .O(n5692) );
  INV_GATE U6147 ( .I1(n5692), .O(n5687) );
  NAND_GATE U6148 ( .I1(n836), .I2(n5687), .O(n5684) );
  NAND_GATE U6149 ( .I1(n1095), .I2(n5128), .O(n5124) );
  NAND3_GATE U6150 ( .I1(n5124), .I2(n5123), .I3(n5122), .O(n5131) );
  OR_GATE U6151 ( .I1(n5126), .I2(n5125), .O(n5130) );
  OR_GATE U6152 ( .I1(n5128), .I2(n5127), .O(n5129) );
  NAND3_GATE U6153 ( .I1(n5131), .I2(n5130), .I3(n5129), .O(n5674) );
  NAND_GATE U6154 ( .I1(B[21]), .I2(A[18]), .O(n5677) );
  INV_GATE U6155 ( .I1(n5677), .O(n5671) );
  NAND_GATE U6156 ( .I1(n5673), .I2(n5671), .O(n5668) );
  NAND_GATE U6157 ( .I1(n937), .I2(n5137), .O(n5134) );
  NAND3_GATE U6158 ( .I1(n5134), .I2(n5133), .I3(n5132), .O(n5140) );
  OR_GATE U6159 ( .I1(n5135), .I2(n893), .O(n5139) );
  OR_GATE U6160 ( .I1(n5137), .I2(n5136), .O(n5138) );
  NAND_GATE U6161 ( .I1(B[21]), .I2(A[17]), .O(n5661) );
  INV_GATE U6162 ( .I1(n5661), .O(n5659) );
  NAND_GATE U6163 ( .I1(n935), .I2(n5659), .O(n5656) );
  NAND_GATE U6164 ( .I1(B[21]), .I2(A[16]), .O(n5646) );
  INV_GATE U6165 ( .I1(n5646), .O(n5642) );
  NAND_GATE U6166 ( .I1(n5144), .I2(n909), .O(n5142) );
  NAND3_GATE U6167 ( .I1(n5143), .I2(n5142), .I3(n5141), .O(n5150) );
  OR_GATE U6168 ( .I1(n5145), .I2(n5144), .O(n5149) );
  OR_GATE U6169 ( .I1(n5147), .I2(n5146), .O(n5148) );
  NAND3_GATE U6170 ( .I1(n5150), .I2(n5149), .I3(n5148), .O(n5643) );
  NAND_GATE U6171 ( .I1(n5642), .I2(n330), .O(n5649) );
  NAND_GATE U6172 ( .I1(n704), .I2(n5157), .O(n5152) );
  NAND3_GATE U6173 ( .I1(n5153), .I2(n5152), .I3(n5151), .O(n5160) );
  OR_GATE U6174 ( .I1(n5155), .I2(n5154), .O(n5159) );
  OR_GATE U6175 ( .I1(n5157), .I2(n5156), .O(n5158) );
  NAND3_GATE U6176 ( .I1(n5160), .I2(n5159), .I3(n5158), .O(n5629) );
  INV_GATE U6177 ( .I1(n5629), .O(n5630) );
  NAND_GATE U6178 ( .I1(B[21]), .I2(A[15]), .O(n5631) );
  NAND_GATE U6179 ( .I1(n5630), .I2(n502), .O(n5634) );
  NAND_GATE U6180 ( .I1(B[21]), .I2(A[14]), .O(n5998) );
  INV_GATE U6181 ( .I1(n5998), .O(n5620) );
  OR_GATE U6182 ( .I1(n5161), .I2(n5167), .O(n5164) );
  OR_GATE U6183 ( .I1(n5166), .I2(n5162), .O(n5163) );
  AND_GATE U6184 ( .I1(n5164), .I2(n5163), .O(n5172) );
  INV_GATE U6185 ( .I1(n5167), .O(n5165) );
  NAND_GATE U6186 ( .I1(n5165), .I2(n5166), .O(n5169) );
  NAND3_GATE U6187 ( .I1(n5170), .I2(n5169), .I3(n5168), .O(n5171) );
  NAND_GATE U6188 ( .I1(n5172), .I2(n5171), .O(n5621) );
  NAND_GATE U6189 ( .I1(n5620), .I2(n302), .O(n5356) );
  NAND_GATE U6190 ( .I1(B[21]), .I2(A[13]), .O(n6024) );
  INV_GATE U6191 ( .I1(n6024), .O(n5449) );
  NAND_GATE U6192 ( .I1(n5174), .I2(n5173), .O(n5175) );
  NAND_GATE U6193 ( .I1(n5176), .I2(n5175), .O(n5177) );
  NAND_GATE U6194 ( .I1(n5181), .I2(n5177), .O(n5179) );
  OR_GATE U6195 ( .I1(n5177), .I2(n5181), .O(n5178) );
  NAND3_GATE U6196 ( .I1(n5180), .I2(n5179), .I3(n5178), .O(n5187) );
  OR_GATE U6197 ( .I1(n5182), .I2(n5181), .O(n5186) );
  OR_GATE U6198 ( .I1(n5184), .I2(n5183), .O(n5185) );
  NAND3_GATE U6199 ( .I1(n5187), .I2(n5186), .I3(n5185), .O(n5452) );
  NAND_GATE U6200 ( .I1(n5449), .I2(n829), .O(n5354) );
  NAND_GATE U6201 ( .I1(B[21]), .I2(A[12]), .O(n6035) );
  INV_GATE U6202 ( .I1(n6035), .O(n5608) );
  NAND_GATE U6203 ( .I1(n680), .I2(n5194), .O(n5191) );
  NAND3_GATE U6204 ( .I1(n5191), .I2(n5190), .I3(n5189), .O(n5197) );
  NAND3_GATE U6205 ( .I1(n5192), .I2(n1222), .I3(n680), .O(n5196) );
  OR_GATE U6206 ( .I1(n5194), .I2(n5193), .O(n5195) );
  NAND3_GATE U6207 ( .I1(n5197), .I2(n5196), .I3(n5195), .O(n5612) );
  INV_GATE U6208 ( .I1(n5612), .O(n5610) );
  NAND_GATE U6209 ( .I1(n5608), .I2(n5610), .O(n5351) );
  NAND_GATE U6210 ( .I1(B[21]), .I2(A[11]), .O(n5471) );
  INV_GATE U6211 ( .I1(n5471), .O(n5460) );
  NAND_GATE U6212 ( .I1(B[21]), .I2(A[10]), .O(n6062) );
  INV_GATE U6213 ( .I1(n6062), .O(n5479) );
  NAND_GATE U6214 ( .I1(n356), .I2(n5210), .O(n5200) );
  NAND_GATE U6215 ( .I1(n5198), .I2(n385), .O(n5199) );
  NAND3_GATE U6216 ( .I1(n5201), .I2(n5200), .I3(n5199), .O(n5213) );
  NAND_GATE U6217 ( .I1(n5202), .I2(n5204), .O(n5207) );
  NAND3_GATE U6218 ( .I1(n5204), .I2(n1301), .I3(n1221), .O(n5206) );
  NAND3_GATE U6219 ( .I1(n5204), .I2(n5203), .I3(n387), .O(n5205) );
  NAND3_GATE U6220 ( .I1(n5207), .I2(n5206), .I3(n5205), .O(n5208) );
  NAND3_GATE U6221 ( .I1(n1223), .I2(n5208), .I3(n356), .O(n5212) );
  OR_GATE U6222 ( .I1(n5210), .I2(n5209), .O(n5211) );
  NAND3_GATE U6223 ( .I1(n5213), .I2(n5212), .I3(n5211), .O(n5477) );
  NAND_GATE U6224 ( .I1(n5479), .I2(n880), .O(n5338) );
  NAND_GATE U6225 ( .I1(B[21]), .I2(A[9]), .O(n5484) );
  INV_GATE U6226 ( .I1(n5484), .O(n5487) );
  NAND_GATE U6227 ( .I1(B[21]), .I2(A[7]), .O(n5504) );
  INV_GATE U6228 ( .I1(n5504), .O(n5294) );
  NAND_GATE U6229 ( .I1(B[21]), .I2(A[5]), .O(n5525) );
  INV_GATE U6230 ( .I1(n5525), .O(n5529) );
  NAND_GATE U6231 ( .I1(n1296), .I2(n5214), .O(n5217) );
  INV_GATE U6232 ( .I1(n5217), .O(n5219) );
  NAND_GATE U6233 ( .I1(n5220), .I2(n5219), .O(n5216) );
  INV_GATE U6234 ( .I1(n5220), .O(n5218) );
  NAND_GATE U6235 ( .I1(n5218), .I2(n5217), .O(n5215) );
  NAND_GATE U6236 ( .I1(n5216), .I2(n5215), .O(n5519) );
  NAND_GATE U6237 ( .I1(n5221), .I2(n5215), .O(n5516) );
  NAND_GATE U6238 ( .I1(n5523), .I2(n5516), .O(n5222) );
  NAND3_GATE U6239 ( .I1(n5221), .I2(n5220), .I3(n5219), .O(n5517) );
  NAND_GATE U6240 ( .I1(n5222), .I2(n5517), .O(n5531) );
  NAND_GATE U6241 ( .I1(n5529), .I2(n5531), .O(n5260) );
  INV_GATE U6242 ( .I1(n5230), .O(n5228) );
  NAND3_GATE U6243 ( .I1(n5223), .I2(n5228), .I3(n5227), .O(n5226) );
  OR_GATE U6244 ( .I1(n5227), .I2(n5224), .O(n5225) );
  AND_GATE U6245 ( .I1(n5226), .I2(n5225), .O(n5236) );
  NAND_GATE U6246 ( .I1(n5228), .I2(n5227), .O(n5234) );
  NAND3_GATE U6247 ( .I1(n5231), .I2(n5230), .I3(n5229), .O(n5233) );
  NAND3_GATE U6248 ( .I1(n5234), .I2(n5233), .I3(n5232), .O(n5235) );
  NAND_GATE U6249 ( .I1(n5236), .I2(n5235), .O(n6083) );
  INV_GATE U6250 ( .I1(n6083), .O(n6085) );
  NAND_GATE U6251 ( .I1(B[21]), .I2(A[4]), .O(n6088) );
  INV_GATE U6252 ( .I1(n6088), .O(n5578) );
  NAND_GATE U6253 ( .I1(n6085), .I2(n5578), .O(n5576) );
  INV_GATE U6254 ( .I1(n5237), .O(n5241) );
  NAND_GATE U6255 ( .I1(n5241), .I2(n5240), .O(n5239) );
  NAND_GATE U6256 ( .I1(n5237), .I2(n5244), .O(n5238) );
  NAND_GATE U6257 ( .I1(n5239), .I2(n5238), .O(n5535) );
  NAND_GATE U6258 ( .I1(n5536), .I2(n5535), .O(n5254) );
  NAND_GATE U6259 ( .I1(n5242), .I2(n5239), .O(n5537) );
  NAND_GATE U6260 ( .I1(B[21]), .I2(A[2]), .O(n5562) );
  INV_GATE U6261 ( .I1(n5562), .O(n5561) );
  NAND_GATE U6262 ( .I1(n1434), .I2(A[0]), .O(n5245) );
  NAND_GATE U6263 ( .I1(n14241), .I2(n5245), .O(n5246) );
  NAND_GATE U6264 ( .I1(B[23]), .I2(n5246), .O(n5250) );
  NAND_GATE U6265 ( .I1(n1435), .I2(A[1]), .O(n5247) );
  NAND_GATE U6266 ( .I1(n724), .I2(n5247), .O(n5248) );
  NAND_GATE U6267 ( .I1(B[22]), .I2(n5248), .O(n5249) );
  NAND_GATE U6268 ( .I1(n5250), .I2(n5249), .O(n5564) );
  NAND_GATE U6269 ( .I1(n5561), .I2(n5564), .O(n5568) );
  NAND3_GATE U6270 ( .I1(B[21]), .I2(B[22]), .I3(n1254), .O(n5569) );
  INV_GATE U6271 ( .I1(n5569), .O(n5563) );
  NAND_GATE U6272 ( .I1(n5562), .I2(n1354), .O(n5251) );
  NAND_GATE U6273 ( .I1(n5563), .I2(n5251), .O(n5252) );
  NAND_GATE U6274 ( .I1(n5568), .I2(n5252), .O(n5546) );
  NAND3_GATE U6275 ( .I1(n5254), .I2(n5253), .I3(n5546), .O(n5256) );
  NAND_GATE U6276 ( .I1(B[21]), .I2(A[3]), .O(n5549) );
  INV_GATE U6277 ( .I1(n5549), .O(n5540) );
  NAND3_GATE U6278 ( .I1(n5254), .I2(n5253), .I3(n5540), .O(n5255) );
  NAND_GATE U6279 ( .I1(n5540), .I2(n5546), .O(n5541) );
  NAND3_GATE U6280 ( .I1(n5256), .I2(n5255), .I3(n5541), .O(n6084) );
  NAND_GATE U6281 ( .I1(n6083), .I2(n6088), .O(n5257) );
  NAND_GATE U6282 ( .I1(n6084), .I2(n5257), .O(n5258) );
  NAND_GATE U6283 ( .I1(n5576), .I2(n5258), .O(n5522) );
  NAND_GATE U6284 ( .I1(n5522), .I2(n5531), .O(n5259) );
  NAND_GATE U6285 ( .I1(n5529), .I2(n5522), .O(n5530) );
  NAND3_GATE U6286 ( .I1(n5260), .I2(n5259), .I3(n5530), .O(n6168) );
  NAND_GATE U6287 ( .I1(B[21]), .I2(A[6]), .O(n5513) );
  INV_GATE U6288 ( .I1(n5277), .O(n5282) );
  NAND_GATE U6289 ( .I1(n5270), .I2(n5261), .O(n5265) );
  NAND3_GATE U6290 ( .I1(n5263), .I2(n5262), .I3(n5261), .O(n5264) );
  NAND_GATE U6291 ( .I1(n5265), .I2(n5264), .O(n5266) );
  NAND_GATE U6292 ( .I1(n5267), .I2(n5266), .O(n5275) );
  NAND_GATE U6293 ( .I1(n5269), .I2(n5268), .O(n5271) );
  NAND_GATE U6294 ( .I1(n5271), .I2(n4681), .O(n5272) );
  NAND_GATE U6295 ( .I1(n5273), .I2(n5272), .O(n5274) );
  NAND3_GATE U6296 ( .I1(n5282), .I2(n5275), .I3(n5274), .O(n5279) );
  NAND_GATE U6297 ( .I1(n5275), .I2(n5274), .O(n5276) );
  NAND_GATE U6298 ( .I1(n5277), .I2(n5276), .O(n5278) );
  NAND3_GATE U6299 ( .I1(n5280), .I2(n5279), .I3(n5278), .O(n6169) );
  NAND3_GATE U6300 ( .I1(n5284), .I2(n5282), .I3(n5281), .O(n6171) );
  NAND3_GATE U6301 ( .I1(n6169), .I2(n6171), .I3(n6170), .O(n5514) );
  NAND_GATE U6302 ( .I1(n5513), .I2(n5514), .O(n5285) );
  NAND_GATE U6303 ( .I1(n6168), .I2(n5285), .O(n5498) );
  INV_GATE U6304 ( .I1(n5513), .O(n6172) );
  NAND_GATE U6305 ( .I1(n6172), .I2(n1322), .O(n5499) );
  NAND_GATE U6306 ( .I1(n5498), .I2(n5499), .O(n5508) );
  NAND_GATE U6307 ( .I1(n5294), .I2(n5508), .O(n5494) );
  INV_GATE U6308 ( .I1(n5288), .O(n5289) );
  NAND3_GATE U6309 ( .I1(n5290), .I2(n5289), .I3(n5287), .O(n5501) );
  NAND3_GATE U6310 ( .I1(n5288), .I2(n398), .I3(n5287), .O(n5500) );
  NAND_GATE U6311 ( .I1(n5290), .I2(n5289), .O(n5292) );
  NAND_GATE U6312 ( .I1(n5293), .I2(n5292), .O(n5502) );
  NAND3_GATE U6313 ( .I1(n5501), .I2(n5500), .I3(n5502), .O(n5291) );
  NAND_GATE U6314 ( .I1(n5503), .I2(n5291), .O(n5509) );
  NAND_GATE U6315 ( .I1(n5508), .I2(n5509), .O(n5297) );
  AND_GATE U6316 ( .I1(n5500), .I2(n5501), .O(n5296) );
  NAND3_GATE U6317 ( .I1(n5293), .I2(n5292), .I3(n5503), .O(n5295) );
  NAND3_GATE U6318 ( .I1(n5296), .I2(n5295), .I3(n5294), .O(n5495) );
  NAND3_GATE U6319 ( .I1(n5494), .I2(n5297), .I3(n5495), .O(n5595) );
  NAND_GATE U6320 ( .I1(B[21]), .I2(A[8]), .O(n6207) );
  NAND3_GATE U6321 ( .I1(n1214), .I2(n5299), .I3(n5298), .O(n5300) );
  NAND4_GATE U6322 ( .I1(n5303), .I2(n5302), .I3(n5301), .I4(n5300), .O(n5304)
         );
  NAND_GATE U6323 ( .I1(n5305), .I2(n5304), .O(n5312) );
  NAND_GATE U6324 ( .I1(n764), .I2(n5312), .O(n5308) );
  NAND3_GATE U6325 ( .I1(n5308), .I2(n5307), .I3(n5306), .O(n5315) );
  NAND4_GATE U6326 ( .I1(n5310), .I2(n764), .I3(n4693), .I4(n5309), .O(n5314)
         );
  OR_GATE U6327 ( .I1(n5312), .I2(n5311), .O(n5313) );
  NAND3_GATE U6328 ( .I1(n5315), .I2(n5314), .I3(n5313), .O(n5592) );
  NAND_GATE U6329 ( .I1(n6207), .I2(n5592), .O(n5316) );
  NAND_GATE U6330 ( .I1(n5595), .I2(n5316), .O(n5318) );
  INV_GATE U6331 ( .I1(n6207), .O(n5591) );
  INV_GATE U6332 ( .I1(n5592), .O(n5594) );
  NAND_GATE U6333 ( .I1(n5591), .I2(n5594), .O(n5317) );
  NAND_GATE U6334 ( .I1(n5318), .I2(n5317), .O(n5482) );
  NAND_GATE U6335 ( .I1(n5487), .I2(n5482), .O(n5489) );
  INV_GATE U6336 ( .I1(n5323), .O(n5322) );
  NAND_GATE U6337 ( .I1(n5321), .I2(n5322), .O(n5320) );
  NAND_GATE U6338 ( .I1(n5325), .I2(n5323), .O(n5332) );
  INV_GATE U6339 ( .I1(n5332), .O(n5319) );
  NAND4_GATE U6340 ( .I1(n5327), .I2(n5326), .I3(n5319), .I4(n5329), .O(n5483)
         );
  NAND3_GATE U6341 ( .I1(n5325), .I2(n5320), .I3(n5483), .O(n5488) );
  NAND3_GATE U6342 ( .I1(n5324), .I2(n5322), .I3(n5321), .O(n5333) );
  NAND3_GATE U6343 ( .I1(n5324), .I2(n5323), .I3(n881), .O(n5331) );
  NAND3_GATE U6344 ( .I1(n5487), .I2(n5488), .I3(n1220), .O(n5335) );
  AND3_GATE U6345 ( .I1(n5327), .I2(n5326), .I3(n5325), .O(n5328) );
  NAND_GATE U6346 ( .I1(n5329), .I2(n5328), .O(n5330) );
  NAND4_GATE U6347 ( .I1(n5333), .I2(n5332), .I3(n5331), .I4(n5330), .O(n5481)
         );
  NAND_GATE U6348 ( .I1(n5483), .I2(n5481), .O(n5490) );
  NAND_GATE U6349 ( .I1(n5482), .I2(n5490), .O(n5334) );
  NAND3_GATE U6350 ( .I1(n5489), .I2(n5335), .I3(n5334), .O(n5478) );
  NAND_GATE U6351 ( .I1(n6062), .I2(n5477), .O(n5336) );
  NAND_GATE U6352 ( .I1(n5478), .I2(n5336), .O(n5337) );
  NAND_GATE U6353 ( .I1(n5338), .I2(n5337), .O(n5465) );
  NAND_GATE U6354 ( .I1(n5460), .I2(n5465), .O(n5348) );
  INV_GATE U6355 ( .I1(n5344), .O(n5339) );
  NAND_GATE U6356 ( .I1(n5340), .I2(n5339), .O(n5342) );
  NAND_GATE U6357 ( .I1(n5343), .I2(n5344), .O(n5341) );
  NAND_GATE U6358 ( .I1(n5342), .I2(n5341), .O(n5466) );
  NAND_GATE U6359 ( .I1(n5345), .I2(n5342), .O(n5457) );
  NAND3_GATE U6360 ( .I1(n5345), .I2(n5344), .I3(n5343), .O(n5456) );
  NAND3_GATE U6361 ( .I1(n5460), .I2(n5463), .I3(n5468), .O(n5347) );
  NAND3_GATE U6362 ( .I1(n5463), .I2(n5468), .I3(n5465), .O(n5346) );
  NAND3_GATE U6363 ( .I1(n5348), .I2(n5347), .I3(n5346), .O(n5609) );
  NAND_GATE U6364 ( .I1(n6035), .I2(n5612), .O(n5349) );
  NAND_GATE U6365 ( .I1(n5609), .I2(n5349), .O(n5350) );
  NAND_GATE U6366 ( .I1(n5351), .I2(n5350), .O(n5450) );
  NAND_GATE U6367 ( .I1(n6024), .I2(n5452), .O(n5352) );
  NAND_GATE U6368 ( .I1(n5450), .I2(n5352), .O(n5353) );
  NAND_GATE U6369 ( .I1(n5354), .I2(n5353), .O(n5622) );
  NAND_GATE U6370 ( .I1(n5356), .I2(n5355), .O(n5635) );
  NAND_GATE U6371 ( .I1(n5629), .I2(n5631), .O(n5357) );
  NAND_GATE U6372 ( .I1(n5635), .I2(n5357), .O(n5358) );
  NAND_GATE U6373 ( .I1(n5634), .I2(n5358), .O(n5650) );
  NAND_GATE U6374 ( .I1(n5646), .I2(n5643), .O(n5359) );
  NAND_GATE U6375 ( .I1(n5650), .I2(n5359), .O(n5360) );
  NAND_GATE U6376 ( .I1(n5649), .I2(n5360), .O(n5660) );
  NAND_GATE U6377 ( .I1(n5660), .I2(n5361), .O(n5362) );
  NAND_GATE U6378 ( .I1(n5656), .I2(n5362), .O(n5672) );
  NAND_GATE U6379 ( .I1(n5674), .I2(n5677), .O(n5363) );
  NAND_GATE U6380 ( .I1(n5672), .I2(n5363), .O(n5364) );
  NAND_GATE U6381 ( .I1(n5686), .I2(n5692), .O(n5365) );
  NAND_GATE U6382 ( .I1(n5688), .I2(n5365), .O(n5366) );
  NAND_GATE U6383 ( .I1(n5684), .I2(n5366), .O(n5439) );
  NAND_GATE U6384 ( .I1(n5437), .I2(n5443), .O(n5367) );
  NAND_GATE U6385 ( .I1(n5439), .I2(n5367), .O(n5368) );
  NAND_GATE U6386 ( .I1(n5435), .I2(n5368), .O(n5704) );
  NAND_GATE U6387 ( .I1(n367), .I2(n5708), .O(n5369) );
  NAND_GATE U6388 ( .I1(n5704), .I2(n5369), .O(n5370) );
  NAND_GATE U6389 ( .I1(n5701), .I2(n5370), .O(n5719) );
  NAND_GATE U6390 ( .I1(n5717), .I2(n5719), .O(n5715) );
  OR_GATE U6391 ( .I1(n5371), .I2(n5376), .O(n5374) );
  OR_GATE U6392 ( .I1(n5375), .I2(n5372), .O(n5373) );
  AND_GATE U6393 ( .I1(n5374), .I2(n5373), .O(n5381) );
  NAND_GATE U6394 ( .I1(n1162), .I2(n5375), .O(n5379) );
  NAND3_GATE U6395 ( .I1(n5379), .I2(n5378), .I3(n5377), .O(n5380) );
  NAND_GATE U6396 ( .I1(n5381), .I2(n5380), .O(n5716) );
  INV_GATE U6397 ( .I1(n5716), .O(n5718) );
  NAND_GATE U6398 ( .I1(n5723), .I2(n366), .O(n5382) );
  NAND_GATE U6399 ( .I1(n5718), .I2(n5382), .O(n5383) );
  NAND_GATE U6400 ( .I1(n5715), .I2(n5383), .O(n5734) );
  NAND_GATE U6401 ( .I1(n5732), .I2(n5739), .O(n5384) );
  NAND_GATE U6402 ( .I1(n5734), .I2(n5384), .O(n5385) );
  NAND_GATE U6403 ( .I1(n5730), .I2(n5385), .O(n5750) );
  NAND_GATE U6404 ( .I1(n5748), .I2(n5755), .O(n5386) );
  NAND_GATE U6405 ( .I1(n5750), .I2(n5386), .O(n5387) );
  NAND_GATE U6406 ( .I1(n5746), .I2(n5387), .O(n5766) );
  NAND_GATE U6407 ( .I1(n5764), .I2(n5771), .O(n5388) );
  NAND_GATE U6408 ( .I1(n5766), .I2(n5388), .O(n5389) );
  NAND_GATE U6409 ( .I1(n5762), .I2(n5389), .O(n5782) );
  NAND_GATE U6410 ( .I1(n5780), .I2(n5787), .O(n5390) );
  NAND_GATE U6411 ( .I1(n5782), .I2(n5390), .O(n5391) );
  NAND_GATE U6412 ( .I1(n5778), .I2(n5391), .O(n5799) );
  NAND_GATE U6413 ( .I1(n5797), .I2(n5804), .O(n5392) );
  NAND_GATE U6414 ( .I1(n5799), .I2(n5392), .O(n5393) );
  NAND_GATE U6415 ( .I1(n5794), .I2(n5393), .O(n5815) );
  NAND_GATE U6416 ( .I1(n5813), .I2(n5820), .O(n5394) );
  NAND_GATE U6417 ( .I1(n5815), .I2(n5394), .O(n5395) );
  NAND_GATE U6418 ( .I1(n5811), .I2(n5395), .O(n5425) );
  NAND_GATE U6419 ( .I1(n5423), .I2(n5430), .O(n5396) );
  NAND_GATE U6420 ( .I1(n5425), .I2(n5396), .O(n5397) );
  NAND_GATE U6421 ( .I1(n5421), .I2(n5397), .O(n5411) );
  NAND_GATE U6422 ( .I1(n5409), .I2(n5416), .O(n5398) );
  NAND_GATE U6423 ( .I1(n5411), .I2(n5398), .O(n5400) );
  NAND_GATE U6424 ( .I1(n1433), .I2(A[31]), .O(n5399) );
  NAND_GATE U6425 ( .I1(n14797), .I2(n5406), .O(n5403) );
  INV_GATE U6426 ( .I1(n5406), .O(n14796) );
  NAND_GATE U6427 ( .I1(n5401), .I2(n14796), .O(n5402) );
  NAND_GATE U6428 ( .I1(n5403), .I2(n5402), .O(\A1[51] ) );
  NAND_GATE U6429 ( .I1(n5404), .I2(n405), .O(n5405) );
  NAND_GATE U6430 ( .I1(n5406), .I2(n5405), .O(n5830) );
  INV_GATE U6431 ( .I1(n5830), .O(n14799) );
  INV_GATE U6432 ( .I1(n5407), .O(n5408) );
  NAND_GATE U6433 ( .I1(n5408), .I2(n5411), .O(n5420) );
  NAND_GATE U6434 ( .I1(n5410), .I2(n5414), .O(n5418) );
  NAND_GATE U6435 ( .I1(n5412), .I2(n5411), .O(n5413) );
  NAND_GATE U6436 ( .I1(n5414), .I2(n5413), .O(n5415) );
  NAND_GATE U6437 ( .I1(n5416), .I2(n5415), .O(n5417) );
  NAND_GATE U6438 ( .I1(n5418), .I2(n5417), .O(n5419) );
  NAND_GATE U6439 ( .I1(n5420), .I2(n5419), .O(n5833) );
  NAND_GATE U6440 ( .I1(B[20]), .I2(A[30]), .O(n5847) );
  INV_GATE U6441 ( .I1(n5847), .O(n5827) );
  INV_GATE U6442 ( .I1(n5421), .O(n5422) );
  NAND_GATE U6443 ( .I1(n5422), .I2(n5425), .O(n5434) );
  NAND_GATE U6444 ( .I1(n5424), .I2(n5428), .O(n5432) );
  NAND_GATE U6445 ( .I1(n5426), .I2(n5425), .O(n5427) );
  NAND_GATE U6446 ( .I1(n5428), .I2(n5427), .O(n5429) );
  NAND_GATE U6447 ( .I1(n5430), .I2(n5429), .O(n5431) );
  NAND_GATE U6448 ( .I1(n5432), .I2(n5431), .O(n5433) );
  NAND_GATE U6449 ( .I1(n5434), .I2(n5433), .O(n5844) );
  NAND_GATE U6450 ( .I1(n5827), .I2(n5844), .O(n5839) );
  NAND_GATE U6451 ( .I1(B[20]), .I2(A[29]), .O(n5858) );
  INV_GATE U6452 ( .I1(n5858), .O(n5825) );
  NAND_GATE U6453 ( .I1(B[20]), .I2(A[28]), .O(n5864) );
  INV_GATE U6454 ( .I1(n5864), .O(n5809) );
  NAND_GATE U6455 ( .I1(B[20]), .I2(A[27]), .O(n5880) );
  INV_GATE U6456 ( .I1(n5880), .O(n5792) );
  NAND_GATE U6457 ( .I1(B[20]), .I2(A[26]), .O(n5891) );
  INV_GATE U6458 ( .I1(n5891), .O(n5776) );
  NAND_GATE U6459 ( .I1(B[20]), .I2(A[25]), .O(n5902) );
  INV_GATE U6460 ( .I1(n5902), .O(n5760) );
  NAND_GATE U6461 ( .I1(B[20]), .I2(A[24]), .O(n5913) );
  INV_GATE U6462 ( .I1(n5913), .O(n5744) );
  NAND_GATE U6463 ( .I1(B[20]), .I2(A[23]), .O(n5924) );
  INV_GATE U6464 ( .I1(n5924), .O(n5728) );
  NAND_GATE U6465 ( .I1(B[20]), .I2(A[22]), .O(n5935) );
  INV_GATE U6466 ( .I1(n5935), .O(n5713) );
  NAND_GATE U6467 ( .I1(B[20]), .I2(A[21]), .O(n5946) );
  INV_GATE U6468 ( .I1(n5946), .O(n5699) );
  INV_GATE U6469 ( .I1(n5435), .O(n5436) );
  NAND_GATE U6470 ( .I1(n5436), .I2(n5439), .O(n5447) );
  NAND_GATE U6471 ( .I1(n5438), .I2(n5441), .O(n5445) );
  NAND_GATE U6472 ( .I1(n798), .I2(n5439), .O(n5440) );
  NAND_GATE U6473 ( .I1(n5441), .I2(n5440), .O(n5442) );
  NAND_GATE U6474 ( .I1(n5443), .I2(n5442), .O(n5444) );
  NAND_GATE U6475 ( .I1(n5445), .I2(n5444), .O(n5446) );
  NAND_GATE U6476 ( .I1(n5447), .I2(n5446), .O(n5944) );
  NAND_GATE U6477 ( .I1(n5699), .I2(n5944), .O(n5941) );
  NAND_GATE U6478 ( .I1(B[20]), .I2(A[20]), .O(n5957) );
  INV_GATE U6479 ( .I1(n5957), .O(n5697) );
  NAND_GATE U6480 ( .I1(B[20]), .I2(A[19]), .O(n6254) );
  INV_GATE U6481 ( .I1(n6254), .O(n5682) );
  NAND_GATE U6482 ( .I1(B[20]), .I2(A[18]), .O(n5968) );
  INV_GATE U6483 ( .I1(n5968), .O(n5666) );
  NAND_GATE U6484 ( .I1(B[20]), .I2(A[17]), .O(n5982) );
  INV_GATE U6485 ( .I1(n5982), .O(n5654) );
  NAND_GATE U6486 ( .I1(B[20]), .I2(A[16]), .O(n5994) );
  INV_GATE U6487 ( .I1(n5994), .O(n5985) );
  NAND_GATE U6488 ( .I1(B[20]), .I2(A[15]), .O(n6008) );
  INV_GATE U6489 ( .I1(n6008), .O(n5625) );
  NAND_GATE U6490 ( .I1(B[20]), .I2(A[14]), .O(n6030) );
  INV_GATE U6491 ( .I1(n6030), .O(n5617) );
  NAND3_GATE U6492 ( .I1(n5449), .I2(n5450), .I3(n829), .O(n6022) );
  INV_GATE U6493 ( .I1(n5450), .O(n5451) );
  NAND_GATE U6494 ( .I1(n5452), .I2(n5451), .O(n5448) );
  NAND_GATE U6495 ( .I1(n5449), .I2(n5448), .O(n6021) );
  NAND_GATE U6496 ( .I1(n829), .I2(n5450), .O(n5454) );
  NAND_GATE U6497 ( .I1(n5454), .I2(n5453), .O(n6023) );
  NAND_GATE U6498 ( .I1(n6021), .I2(n6027), .O(n5455) );
  NAND_GATE U6499 ( .I1(n6022), .I2(n5455), .O(n6017) );
  NAND_GATE U6500 ( .I1(n5617), .I2(n6017), .O(n6016) );
  NAND_GATE U6501 ( .I1(B[20]), .I2(A[13]), .O(n6038) );
  INV_GATE U6502 ( .I1(n6038), .O(n5615) );
  AND3_GATE U6503 ( .I1(n5456), .I2(n5465), .I3(n5460), .O(n5459) );
  NAND_GATE U6504 ( .I1(n5457), .I2(n5463), .O(n5458) );
  NAND_GATE U6505 ( .I1(n5459), .I2(n5458), .O(n5462) );
  NAND4_GATE U6506 ( .I1(n5468), .I2(n5463), .I3(n5460), .I4(n361), .O(n5461)
         );
  AND_GATE U6507 ( .I1(n5462), .I2(n5461), .O(n5473) );
  NAND_GATE U6508 ( .I1(n5467), .I2(n5466), .O(n5463) );
  NAND_GATE U6509 ( .I1(n5468), .I2(n5463), .O(n5464) );
  NAND_GATE U6510 ( .I1(n5465), .I2(n5464), .O(n5470) );
  NAND3_GATE U6511 ( .I1(n5468), .I2(n5463), .I3(n361), .O(n5469) );
  NAND3_GATE U6512 ( .I1(n5471), .I2(n5470), .I3(n5469), .O(n5472) );
  NAND_GATE U6513 ( .I1(n5473), .I2(n5472), .O(n6057) );
  NAND_GATE U6514 ( .I1(B[20]), .I2(A[12]), .O(n6056) );
  INV_GATE U6515 ( .I1(n6056), .O(n6054) );
  NAND_GATE U6516 ( .I1(n355), .I2(n6054), .O(n6052) );
  NAND_GATE U6517 ( .I1(B[20]), .I2(A[11]), .O(n6069) );
  INV_GATE U6518 ( .I1(n6069), .O(n5604) );
  NAND_GATE U6519 ( .I1(n880), .I2(n5478), .O(n5475) );
  INV_GATE U6520 ( .I1(n5478), .O(n5476) );
  NAND_GATE U6521 ( .I1(n5477), .I2(n5476), .O(n5474) );
  NAND_GATE U6522 ( .I1(n5475), .I2(n5474), .O(n6061) );
  NAND_GATE U6523 ( .I1(n5479), .I2(n5474), .O(n6063) );
  NAND_GATE U6524 ( .I1(n6066), .I2(n6063), .O(n5480) );
  NAND3_GATE U6525 ( .I1(n5479), .I2(n5478), .I3(n880), .O(n6064) );
  NAND_GATE U6526 ( .I1(n5480), .I2(n6064), .O(n6072) );
  NAND_GATE U6527 ( .I1(n5604), .I2(n6072), .O(n6074) );
  NAND_GATE U6528 ( .I1(B[20]), .I2(A[10]), .O(n6369) );
  INV_GATE U6529 ( .I1(n6369), .O(n6220) );
  NAND_GATE U6530 ( .I1(n299), .I2(n5490), .O(n5486) );
  NAND3_GATE U6531 ( .I1(n5483), .I2(n5482), .I3(n5481), .O(n5485) );
  NAND3_GATE U6532 ( .I1(n5486), .I2(n5485), .I3(n5484), .O(n5493) );
  NAND4_GATE U6533 ( .I1(n5488), .I2(n299), .I3(n5487), .I4(n1220), .O(n5492)
         );
  OR_GATE U6534 ( .I1(n5490), .I2(n5489), .O(n5491) );
  NAND3_GATE U6535 ( .I1(n5493), .I2(n5492), .I3(n5491), .O(n6221) );
  INV_GATE U6536 ( .I1(n6221), .O(n6222) );
  NAND_GATE U6537 ( .I1(n6220), .I2(n6222), .O(n5603) );
  NAND_GATE U6538 ( .I1(B[20]), .I2(A[9]), .O(n6214) );
  INV_GATE U6539 ( .I1(n6214), .O(n5598) );
  OR_GATE U6540 ( .I1(n5509), .I2(n5494), .O(n5497) );
  OR_GATE U6541 ( .I1(n5495), .I2(n5508), .O(n5496) );
  NAND_GATE U6542 ( .I1(n5497), .I2(n5496), .O(n6193) );
  NAND3_GATE U6543 ( .I1(n5499), .I2(n5498), .I3(n5504), .O(n5507) );
  NAND4_GATE U6544 ( .I1(n5502), .I2(n5504), .I3(n5501), .I4(n5500), .O(n5506)
         );
  NAND3_GATE U6545 ( .I1(n5507), .I2(n5506), .I3(n5505), .O(n5512) );
  INV_GATE U6546 ( .I1(n5508), .O(n5510) );
  NAND_GATE U6547 ( .I1(n5510), .I2(n5509), .O(n5511) );
  INV_GATE U6548 ( .I1(n6197), .O(n6200) );
  NAND_GATE U6549 ( .I1(B[20]), .I2(A[8]), .O(n6198) );
  INV_GATE U6550 ( .I1(n6198), .O(n6196) );
  NAND_GATE U6551 ( .I1(n6200), .I2(n6196), .O(n6192) );
  NAND3_GATE U6552 ( .I1(n6168), .I2(n5513), .I3(n1322), .O(n6173) );
  NAND_GATE U6553 ( .I1(B[20]), .I2(A[7]), .O(n6182) );
  INV_GATE U6554 ( .I1(n6182), .O(n5586) );
  NAND3_GATE U6555 ( .I1(n6168), .I2(n6172), .I3(n1322), .O(n6178) );
  NAND3_GATE U6556 ( .I1(n5515), .I2(n6178), .I3(n6172), .O(n5585) );
  NAND_GATE U6557 ( .I1(n1209), .I2(n1258), .O(n5588) );
  INV_GATE U6558 ( .I1(n5516), .O(n5518) );
  NAND_GATE U6559 ( .I1(n5518), .I2(n5517), .O(n5524) );
  NAND_GATE U6560 ( .I1(n5520), .I2(n5519), .O(n5523) );
  NAND_GATE U6561 ( .I1(n5524), .I2(n5523), .O(n5521) );
  NAND_GATE U6562 ( .I1(n5522), .I2(n5521), .O(n5527) );
  INV_GATE U6563 ( .I1(n5522), .O(n5528) );
  NAND3_GATE U6564 ( .I1(n5524), .I2(n5523), .I3(n5528), .O(n5526) );
  NAND3_GATE U6565 ( .I1(n5527), .I2(n5526), .I3(n5525), .O(n5534) );
  NAND3_GATE U6566 ( .I1(n5529), .I2(n5528), .I3(n5531), .O(n5533) );
  OR_GATE U6567 ( .I1(n5531), .I2(n5530), .O(n5532) );
  NAND3_GATE U6568 ( .I1(n5534), .I2(n5533), .I3(n5532), .O(n6158) );
  INV_GATE U6569 ( .I1(n6158), .O(n6154) );
  NAND_GATE U6570 ( .I1(B[20]), .I2(A[6]), .O(n6156) );
  INV_GATE U6571 ( .I1(n6156), .O(n6163) );
  NAND_GATE U6572 ( .I1(n6154), .I2(n6163), .O(n6153) );
  INV_GATE U6573 ( .I1(n5546), .O(n5544) );
  NAND_GATE U6574 ( .I1(n5537), .I2(n5254), .O(n5538) );
  NAND_GATE U6575 ( .I1(n5539), .I2(n5538), .O(n5545) );
  OR_GATE U6576 ( .I1(n5545), .I2(n5541), .O(n5542) );
  AND_GATE U6577 ( .I1(n5543), .I2(n5542), .O(n5551) );
  NAND_GATE U6578 ( .I1(n5544), .I2(n5545), .O(n5548) );
  NAND3_GATE U6579 ( .I1(n5549), .I2(n5548), .I3(n5547), .O(n5550) );
  NAND_GATE U6580 ( .I1(n5551), .I2(n5550), .O(n6142) );
  NAND_GATE U6581 ( .I1(B[20]), .I2(A[4]), .O(n6141) );
  INV_GATE U6582 ( .I1(n6141), .O(n6144) );
  NAND_GATE U6583 ( .I1(B[20]), .I2(A[3]), .O(n6104) );
  INV_GATE U6584 ( .I1(n6104), .O(n5572) );
  NAND_GATE U6585 ( .I1(B[20]), .I2(A[2]), .O(n6126) );
  INV_GATE U6586 ( .I1(n6126), .O(n6122) );
  NAND_GATE U6587 ( .I1(n1433), .I2(A[0]), .O(n5552) );
  NAND_GATE U6588 ( .I1(n14241), .I2(n5552), .O(n5553) );
  NAND_GATE U6589 ( .I1(B[22]), .I2(n5553), .O(n5557) );
  NAND_GATE U6590 ( .I1(n1434), .I2(A[1]), .O(n5554) );
  NAND_GATE U6591 ( .I1(n724), .I2(n5554), .O(n5555) );
  NAND_GATE U6592 ( .I1(B[21]), .I2(n5555), .O(n5556) );
  NAND_GATE U6593 ( .I1(n5557), .I2(n5556), .O(n6124) );
  NAND_GATE U6594 ( .I1(n6122), .I2(n6124), .O(n6120) );
  NAND3_GATE U6595 ( .I1(B[20]), .I2(B[21]), .I3(n1254), .O(n6125) );
  INV_GATE U6596 ( .I1(n6125), .O(n6123) );
  NAND_GATE U6597 ( .I1(n6126), .I2(n1370), .O(n5558) );
  NAND_GATE U6598 ( .I1(n6123), .I2(n5558), .O(n5559) );
  NAND_GATE U6599 ( .I1(n6120), .I2(n5559), .O(n6105) );
  NAND_GATE U6600 ( .I1(n5572), .I2(n6105), .O(n6107) );
  NAND_GATE U6601 ( .I1(n1354), .I2(n5569), .O(n5560) );
  NAND_GATE U6602 ( .I1(n5561), .I2(n5560), .O(n5567) );
  NAND3_GATE U6603 ( .I1(n1354), .I2(n5562), .I3(n5569), .O(n5566) );
  NAND_GATE U6604 ( .I1(n5564), .I2(n5563), .O(n5565) );
  NAND3_GATE U6605 ( .I1(n5567), .I2(n5566), .I3(n5565), .O(n5571) );
  OR_GATE U6606 ( .I1(n5569), .I2(n5568), .O(n5570) );
  NAND_GATE U6607 ( .I1(n5571), .I2(n5570), .O(n6108) );
  NAND_GATE U6608 ( .I1(n6105), .I2(n6108), .O(n5573) );
  NAND_GATE U6609 ( .I1(n5572), .I2(n6108), .O(n6106) );
  NAND3_GATE U6610 ( .I1(n6107), .I2(n5573), .I3(n6106), .O(n6138) );
  NAND_GATE U6611 ( .I1(n6142), .I2(n6141), .O(n5574) );
  NAND_GATE U6612 ( .I1(n6138), .I2(n5574), .O(n5575) );
  NAND_GATE U6613 ( .I1(n6136), .I2(n5575), .O(n6092) );
  INV_GATE U6614 ( .I1(n6084), .O(n6082) );
  NAND3_GATE U6615 ( .I1(n6088), .I2(n6082), .I3(n6083), .O(n5579) );
  NAND_GATE U6616 ( .I1(n6083), .I2(n6082), .O(n5577) );
  NAND_GATE U6617 ( .I1(n5578), .I2(n5577), .O(n6079) );
  NAND3_GATE U6618 ( .I1(n5579), .I2(n6086), .I3(n6079), .O(n5580) );
  NAND_GATE U6619 ( .I1(n6081), .I2(n5580), .O(n6098) );
  NAND_GATE U6620 ( .I1(n6092), .I2(n6098), .O(n5582) );
  NAND_GATE U6621 ( .I1(B[20]), .I2(A[5]), .O(n6093) );
  INV_GATE U6622 ( .I1(n6093), .O(n6096) );
  NAND_GATE U6623 ( .I1(n6096), .I2(n6098), .O(n5581) );
  NAND_GATE U6624 ( .I1(n6096), .I2(n6092), .O(n6097) );
  NAND3_GATE U6625 ( .I1(n5582), .I2(n5581), .I3(n6097), .O(n6155) );
  NAND_GATE U6626 ( .I1(n6158), .I2(n6156), .O(n5583) );
  NAND_GATE U6627 ( .I1(n6155), .I2(n5583), .O(n5584) );
  NAND_GATE U6628 ( .I1(n6153), .I2(n5584), .O(n6179) );
  NAND3_GATE U6629 ( .I1(n5585), .I2(n1209), .I3(n6179), .O(n5587) );
  NAND_GATE U6630 ( .I1(n5586), .I2(n6179), .O(n6184) );
  NAND_GATE U6631 ( .I1(n6197), .I2(n6198), .O(n5589) );
  NAND_GATE U6632 ( .I1(n6199), .I2(n5589), .O(n5590) );
  NAND_GATE U6633 ( .I1(n5598), .I2(n6211), .O(n6204) );
  INV_GATE U6634 ( .I1(n5595), .O(n5593) );
  NAND_GATE U6635 ( .I1(n5591), .I2(n5597), .O(n6203) );
  NAND_GATE U6636 ( .I1(n5593), .I2(n5592), .O(n5597) );
  NAND_GATE U6637 ( .I1(n5595), .I2(n5594), .O(n5596) );
  NAND_GATE U6638 ( .I1(n5597), .I2(n5596), .O(n6206) );
  NAND_GATE U6639 ( .I1(n6207), .I2(n6206), .O(n6205) );
  NAND3_GATE U6640 ( .I1(n6211), .I2(n6209), .I3(n6205), .O(n5600) );
  NAND_GATE U6641 ( .I1(n6205), .I2(n1384), .O(n5599) );
  NAND_GATE U6642 ( .I1(n6369), .I2(n6221), .O(n5601) );
  NAND_GATE U6643 ( .I1(n5), .I2(n5601), .O(n5602) );
  NAND_GATE U6644 ( .I1(n5603), .I2(n5602), .O(n6075) );
  NAND_GATE U6645 ( .I1(n6072), .I2(n6075), .O(n5605) );
  NAND_GATE U6646 ( .I1(n5604), .I2(n6075), .O(n6073) );
  NAND_GATE U6647 ( .I1(n6057), .I2(n6056), .O(n5606) );
  NAND_GATE U6648 ( .I1(n6055), .I2(n5606), .O(n5607) );
  NAND_GATE U6649 ( .I1(n6052), .I2(n5607), .O(n6041) );
  NAND_GATE U6650 ( .I1(n5615), .I2(n6041), .O(n6045) );
  INV_GATE U6651 ( .I1(n5609), .O(n5611) );
  NAND_GATE U6652 ( .I1(n5608), .I2(n5613), .O(n6044) );
  NAND3_GATE U6653 ( .I1(n5608), .I2(n5609), .I3(n5610), .O(n6046) );
  NAND_GATE U6654 ( .I1(n5610), .I2(n5609), .O(n5614) );
  NAND_GATE U6655 ( .I1(n5612), .I2(n5611), .O(n5613) );
  NAND_GATE U6656 ( .I1(n5614), .I2(n5613), .O(n6034) );
  NAND_GATE U6657 ( .I1(n6035), .I2(n6034), .O(n6043) );
  NAND3_GATE U6658 ( .I1(n5615), .I2(n6036), .I3(n6043), .O(n6042) );
  NAND3_GATE U6659 ( .I1(n6041), .I2(n6036), .I3(n6043), .O(n5616) );
  NAND3_GATE U6660 ( .I1(n6045), .I2(n6042), .I3(n5616), .O(n6029) );
  NAND_GATE U6661 ( .I1(n6017), .I2(n6029), .O(n5618) );
  NAND_GATE U6662 ( .I1(n5617), .I2(n6029), .O(n6018) );
  NAND3_GATE U6663 ( .I1(n6016), .I2(n5618), .I3(n6018), .O(n6009) );
  NAND_GATE U6664 ( .I1(n5625), .I2(n6009), .O(n6011) );
  NAND3_GATE U6665 ( .I1(n5622), .I2(n302), .I3(n5620), .O(n6001) );
  NAND_GATE U6666 ( .I1(n5621), .I2(n782), .O(n5619) );
  NAND_GATE U6667 ( .I1(n5620), .I2(n5619), .O(n5999) );
  NAND_GATE U6668 ( .I1(n5619), .I2(n5623), .O(n5997) );
  NAND_GATE U6669 ( .I1(n5999), .I2(n6005), .O(n5624) );
  NAND_GATE U6670 ( .I1(n6001), .I2(n5624), .O(n6012) );
  NAND_GATE U6671 ( .I1(n5625), .I2(n6012), .O(n6010) );
  NAND_GATE U6672 ( .I1(n6009), .I2(n6012), .O(n5626) );
  NAND3_GATE U6673 ( .I1(n6011), .I2(n6010), .I3(n5626), .O(n5991) );
  NAND_GATE U6674 ( .I1(n5985), .I2(n5991), .O(n5986) );
  INV_GATE U6675 ( .I1(n5635), .O(n5628) );
  NAND_GATE U6676 ( .I1(n5629), .I2(n5628), .O(n5627) );
  NAND_GATE U6677 ( .I1(n502), .I2(n5627), .O(n5633) );
  NAND_GATE U6678 ( .I1(n5633), .I2(n5632), .O(n5638) );
  INV_GATE U6679 ( .I1(n5634), .O(n5636) );
  NAND_GATE U6680 ( .I1(n5636), .I2(n5635), .O(n5637) );
  NAND_GATE U6681 ( .I1(n5638), .I2(n5637), .O(n5990) );
  NAND_GATE U6682 ( .I1(n5985), .I2(n5990), .O(n5640) );
  NAND_GATE U6683 ( .I1(n5991), .I2(n5990), .O(n5639) );
  NAND3_GATE U6684 ( .I1(n5986), .I2(n5640), .I3(n5639), .O(n5979) );
  NAND_GATE U6685 ( .I1(n5654), .I2(n5979), .O(n5974) );
  NAND_GATE U6686 ( .I1(n5642), .I2(n5641), .O(n5648) );
  NAND_GATE U6687 ( .I1(n330), .I2(n5650), .O(n5644) );
  NAND_GATE U6688 ( .I1(n5644), .I2(n5641), .O(n5645) );
  NAND_GATE U6689 ( .I1(n5646), .I2(n5645), .O(n5647) );
  NAND_GATE U6690 ( .I1(n5648), .I2(n5647), .O(n5653) );
  INV_GATE U6691 ( .I1(n5649), .O(n5651) );
  NAND_GATE U6692 ( .I1(n5651), .I2(n5650), .O(n5652) );
  NAND_GATE U6693 ( .I1(n5653), .I2(n5652), .O(n5978) );
  NAND_GATE U6694 ( .I1(n5979), .I2(n5978), .O(n5655) );
  NAND3_GATE U6695 ( .I1(n5974), .I2(n5973), .I3(n5655), .O(n5967) );
  NAND_GATE U6696 ( .I1(n5666), .I2(n5967), .O(n5963) );
  INV_GATE U6697 ( .I1(n5656), .O(n5657) );
  NAND_GATE U6698 ( .I1(n5657), .I2(n5660), .O(n5665) );
  NAND_GATE U6699 ( .I1(n5659), .I2(n5658), .O(n5663) );
  NAND_GATE U6700 ( .I1(n5663), .I2(n5662), .O(n5664) );
  NAND_GATE U6701 ( .I1(n5665), .I2(n5664), .O(n5966) );
  NAND_GATE U6702 ( .I1(n5967), .I2(n5966), .O(n5667) );
  NAND3_GATE U6703 ( .I1(n5963), .I2(n5962), .I3(n5667), .O(n6253) );
  NAND_GATE U6704 ( .I1(n5682), .I2(n6253), .O(n6249) );
  INV_GATE U6705 ( .I1(n5668), .O(n5669) );
  NAND_GATE U6706 ( .I1(n5669), .I2(n5672), .O(n5681) );
  NAND_GATE U6707 ( .I1(n5671), .I2(n5670), .O(n5679) );
  NAND_GATE U6708 ( .I1(n5673), .I2(n5672), .O(n5675) );
  NAND_GATE U6709 ( .I1(n5675), .I2(n5670), .O(n5676) );
  NAND_GATE U6710 ( .I1(n5677), .I2(n5676), .O(n5678) );
  NAND_GATE U6711 ( .I1(n5679), .I2(n5678), .O(n5680) );
  NAND_GATE U6712 ( .I1(n5681), .I2(n5680), .O(n6252) );
  NAND_GATE U6713 ( .I1(n5682), .I2(n6252), .O(n6248) );
  NAND_GATE U6714 ( .I1(n6253), .I2(n6252), .O(n5683) );
  NAND3_GATE U6715 ( .I1(n6249), .I2(n6248), .I3(n5683), .O(n5956) );
  NAND_GATE U6716 ( .I1(n5697), .I2(n5956), .O(n5952) );
  INV_GATE U6717 ( .I1(n5684), .O(n5685) );
  NAND_GATE U6718 ( .I1(n5685), .I2(n5688), .O(n5696) );
  NAND_GATE U6719 ( .I1(n5687), .I2(n5690), .O(n5694) );
  NAND_GATE U6720 ( .I1(n5690), .I2(n5689), .O(n5691) );
  NAND_GATE U6721 ( .I1(n5692), .I2(n5691), .O(n5693) );
  NAND_GATE U6722 ( .I1(n5694), .I2(n5693), .O(n5695) );
  NAND_GATE U6723 ( .I1(n5696), .I2(n5695), .O(n5955) );
  NAND_GATE U6724 ( .I1(n5956), .I2(n5955), .O(n5698) );
  NAND3_GATE U6725 ( .I1(n5952), .I2(n5951), .I3(n5698), .O(n5945) );
  NAND_GATE U6726 ( .I1(n5699), .I2(n5945), .O(n5940) );
  NAND_GATE U6727 ( .I1(n5944), .I2(n5945), .O(n5700) );
  NAND3_GATE U6728 ( .I1(n5941), .I2(n5940), .I3(n5700), .O(n5934) );
  NAND_GATE U6729 ( .I1(n5713), .I2(n5934), .O(n5929) );
  INV_GATE U6730 ( .I1(n5701), .O(n5702) );
  NAND_GATE U6731 ( .I1(n5702), .I2(n5704), .O(n5712) );
  NAND_GATE U6732 ( .I1(n5703), .I2(n5706), .O(n5710) );
  NAND_GATE U6733 ( .I1(n800), .I2(n5704), .O(n5705) );
  NAND_GATE U6734 ( .I1(n5706), .I2(n5705), .O(n5707) );
  NAND_GATE U6735 ( .I1(n5708), .I2(n5707), .O(n5709) );
  NAND_GATE U6736 ( .I1(n5710), .I2(n5709), .O(n5711) );
  NAND_GATE U6737 ( .I1(n5712), .I2(n5711), .O(n5933) );
  NAND_GATE U6738 ( .I1(n5713), .I2(n5933), .O(n5928) );
  NAND_GATE U6739 ( .I1(n5934), .I2(n5933), .O(n5714) );
  NAND3_GATE U6740 ( .I1(n5929), .I2(n5928), .I3(n5714), .O(n5923) );
  NAND_GATE U6741 ( .I1(n5728), .I2(n5923), .O(n5919) );
  OR_GATE U6742 ( .I1(n5716), .I2(n5715), .O(n5727) );
  NAND_GATE U6743 ( .I1(n366), .I2(n5716), .O(n5721) );
  NAND_GATE U6744 ( .I1(n5717), .I2(n5721), .O(n5725) );
  NAND_GATE U6745 ( .I1(n5719), .I2(n5718), .O(n5720) );
  NAND_GATE U6746 ( .I1(n5721), .I2(n5720), .O(n5722) );
  NAND_GATE U6747 ( .I1(n5723), .I2(n5722), .O(n5724) );
  NAND_GATE U6748 ( .I1(n5725), .I2(n5724), .O(n5726) );
  NAND_GATE U6749 ( .I1(n5727), .I2(n5726), .O(n5922) );
  NAND_GATE U6750 ( .I1(n5728), .I2(n5922), .O(n5918) );
  NAND_GATE U6751 ( .I1(n5923), .I2(n5922), .O(n5729) );
  NAND3_GATE U6752 ( .I1(n5919), .I2(n5918), .I3(n5729), .O(n5912) );
  NAND_GATE U6753 ( .I1(n5744), .I2(n5912), .O(n5908) );
  INV_GATE U6754 ( .I1(n5730), .O(n5731) );
  NAND_GATE U6755 ( .I1(n5731), .I2(n5734), .O(n5743) );
  NAND_GATE U6756 ( .I1(n5733), .I2(n5737), .O(n5741) );
  NAND_GATE U6757 ( .I1(n5735), .I2(n5734), .O(n5736) );
  NAND_GATE U6758 ( .I1(n5737), .I2(n5736), .O(n5738) );
  NAND_GATE U6759 ( .I1(n5739), .I2(n5738), .O(n5740) );
  NAND_GATE U6760 ( .I1(n5741), .I2(n5740), .O(n5742) );
  NAND_GATE U6761 ( .I1(n5743), .I2(n5742), .O(n5911) );
  NAND_GATE U6762 ( .I1(n5912), .I2(n5911), .O(n5745) );
  NAND3_GATE U6763 ( .I1(n5908), .I2(n5907), .I3(n5745), .O(n5901) );
  NAND_GATE U6764 ( .I1(n5760), .I2(n5901), .O(n5897) );
  INV_GATE U6765 ( .I1(n5746), .O(n5747) );
  NAND_GATE U6766 ( .I1(n5747), .I2(n5750), .O(n5759) );
  NAND_GATE U6767 ( .I1(n5749), .I2(n5753), .O(n5757) );
  NAND_GATE U6768 ( .I1(n5751), .I2(n5750), .O(n5752) );
  NAND_GATE U6769 ( .I1(n5753), .I2(n5752), .O(n5754) );
  NAND_GATE U6770 ( .I1(n5755), .I2(n5754), .O(n5756) );
  NAND_GATE U6771 ( .I1(n5757), .I2(n5756), .O(n5758) );
  NAND_GATE U6772 ( .I1(n5759), .I2(n5758), .O(n5900) );
  NAND_GATE U6773 ( .I1(n5760), .I2(n5900), .O(n5896) );
  NAND_GATE U6774 ( .I1(n5901), .I2(n5900), .O(n5761) );
  NAND3_GATE U6775 ( .I1(n5897), .I2(n5896), .I3(n5761), .O(n5890) );
  NAND_GATE U6776 ( .I1(n5776), .I2(n5890), .O(n5886) );
  INV_GATE U6777 ( .I1(n5762), .O(n5763) );
  NAND_GATE U6778 ( .I1(n5763), .I2(n5766), .O(n5775) );
  NAND_GATE U6779 ( .I1(n5765), .I2(n5769), .O(n5773) );
  NAND_GATE U6780 ( .I1(n5767), .I2(n5766), .O(n5768) );
  NAND_GATE U6781 ( .I1(n5769), .I2(n5768), .O(n5770) );
  NAND_GATE U6782 ( .I1(n5771), .I2(n5770), .O(n5772) );
  NAND_GATE U6783 ( .I1(n5773), .I2(n5772), .O(n5774) );
  NAND_GATE U6784 ( .I1(n5775), .I2(n5774), .O(n5889) );
  NAND_GATE U6785 ( .I1(n5776), .I2(n5889), .O(n5885) );
  NAND_GATE U6786 ( .I1(n5890), .I2(n5889), .O(n5777) );
  NAND3_GATE U6787 ( .I1(n5886), .I2(n5885), .I3(n5777), .O(n5879) );
  NAND_GATE U6788 ( .I1(n5792), .I2(n5879), .O(n5875) );
  INV_GATE U6789 ( .I1(n5778), .O(n5779) );
  NAND_GATE U6790 ( .I1(n5779), .I2(n5782), .O(n5791) );
  NAND_GATE U6791 ( .I1(n5781), .I2(n5785), .O(n5789) );
  NAND_GATE U6792 ( .I1(n5783), .I2(n5782), .O(n5784) );
  NAND_GATE U6793 ( .I1(n5785), .I2(n5784), .O(n5786) );
  NAND_GATE U6794 ( .I1(n5787), .I2(n5786), .O(n5788) );
  NAND_GATE U6795 ( .I1(n5789), .I2(n5788), .O(n5790) );
  NAND_GATE U6796 ( .I1(n5791), .I2(n5790), .O(n5878) );
  NAND_GATE U6797 ( .I1(n5792), .I2(n5878), .O(n5874) );
  NAND_GATE U6798 ( .I1(n5879), .I2(n5878), .O(n5793) );
  NAND3_GATE U6799 ( .I1(n5875), .I2(n5874), .I3(n5793), .O(n5863) );
  NAND_GATE U6800 ( .I1(n5809), .I2(n5863), .O(n5867) );
  INV_GATE U6801 ( .I1(n5794), .O(n5795) );
  NAND_GATE U6802 ( .I1(n5795), .I2(n5799), .O(n5808) );
  INV_GATE U6803 ( .I1(n5799), .O(n5796) );
  NAND_GATE U6804 ( .I1(n5797), .I2(n5796), .O(n5802) );
  NAND_GATE U6805 ( .I1(n5798), .I2(n5802), .O(n5806) );
  NAND_GATE U6806 ( .I1(n5800), .I2(n5799), .O(n5801) );
  NAND_GATE U6807 ( .I1(n5802), .I2(n5801), .O(n5803) );
  NAND_GATE U6808 ( .I1(n5804), .I2(n5803), .O(n5805) );
  NAND_GATE U6809 ( .I1(n5806), .I2(n5805), .O(n5807) );
  NAND_GATE U6810 ( .I1(n5808), .I2(n5807), .O(n5868) );
  NAND_GATE U6811 ( .I1(n5809), .I2(n5868), .O(n5871) );
  NAND_GATE U6812 ( .I1(n5863), .I2(n5868), .O(n5810) );
  NAND3_GATE U6813 ( .I1(n5867), .I2(n5871), .I3(n5810), .O(n5857) );
  NAND_GATE U6814 ( .I1(n5825), .I2(n5857), .O(n5853) );
  INV_GATE U6815 ( .I1(n5811), .O(n5812) );
  NAND_GATE U6816 ( .I1(n5812), .I2(n5815), .O(n5824) );
  NAND_GATE U6817 ( .I1(n5814), .I2(n5818), .O(n5822) );
  NAND_GATE U6818 ( .I1(n5816), .I2(n5815), .O(n5817) );
  NAND_GATE U6819 ( .I1(n5818), .I2(n5817), .O(n5819) );
  NAND_GATE U6820 ( .I1(n5820), .I2(n5819), .O(n5821) );
  NAND_GATE U6821 ( .I1(n5822), .I2(n5821), .O(n5823) );
  NAND_GATE U6822 ( .I1(n5824), .I2(n5823), .O(n5856) );
  NAND_GATE U6823 ( .I1(n5825), .I2(n5856), .O(n5852) );
  NAND_GATE U6824 ( .I1(n5857), .I2(n5856), .O(n5826) );
  NAND3_GATE U6825 ( .I1(n5853), .I2(n5852), .I3(n5826), .O(n5846) );
  NAND_GATE U6826 ( .I1(n5846), .I2(n5844), .O(n5828) );
  NAND_GATE U6827 ( .I1(n5827), .I2(n5846), .O(n5840) );
  AND3_GATE U6828 ( .I1(n5839), .I2(n5828), .I3(n5840), .O(n5835) );
  NAND_GATE U6829 ( .I1(n1432), .I2(A[31]), .O(n5834) );
  NAND_GATE U6830 ( .I1(n5835), .I2(n5834), .O(n5829) );
  NAND_GATE U6831 ( .I1(n5833), .I2(n5829), .O(n5838) );
  NAND_GATE U6832 ( .I1(n14799), .I2(n5838), .O(n5832) );
  INV_GATE U6833 ( .I1(n5838), .O(n14798) );
  NAND_GATE U6834 ( .I1(n5830), .I2(n14798), .O(n5831) );
  NAND_GATE U6835 ( .I1(n5832), .I2(n5831), .O(\A1[50] ) );
  INV_GATE U6836 ( .I1(n5833), .O(n5836) );
  NAND3_GATE U6837 ( .I1(n5836), .I2(n5835), .I3(n5834), .O(n5837) );
  NAND_GATE U6838 ( .I1(n5838), .I2(n5837), .O(n6283) );
  INV_GATE U6839 ( .I1(n6283), .O(n14801) );
  OR_GATE U6840 ( .I1(n5839), .I2(n5846), .O(n5842) );
  OR_GATE U6841 ( .I1(n5844), .I2(n5840), .O(n5841) );
  AND_GATE U6842 ( .I1(n5842), .I2(n5841), .O(n5851) );
  INV_GATE U6843 ( .I1(n5846), .O(n5843) );
  NAND_GATE U6844 ( .I1(n5843), .I2(n5844), .O(n5849) );
  INV_GATE U6845 ( .I1(n5844), .O(n5845) );
  NAND_GATE U6846 ( .I1(n5846), .I2(n5845), .O(n5848) );
  NAND3_GATE U6847 ( .I1(n5849), .I2(n5848), .I3(n5847), .O(n5850) );
  OR_GATE U6848 ( .I1(n5852), .I2(n5857), .O(n5855) );
  OR_GATE U6849 ( .I1(n5856), .I2(n5853), .O(n5854) );
  AND_GATE U6850 ( .I1(n5855), .I2(n5854), .O(n5862) );
  NAND_GATE U6851 ( .I1(n1163), .I2(n5856), .O(n5860) );
  NAND3_GATE U6852 ( .I1(n5860), .I2(n5859), .I3(n5858), .O(n5861) );
  NAND_GATE U6853 ( .I1(n5862), .I2(n5861), .O(n6290) );
  INV_GATE U6854 ( .I1(n6290), .O(n6293) );
  NAND_GATE U6855 ( .I1(B[19]), .I2(A[30]), .O(n6714) );
  INV_GATE U6856 ( .I1(n6714), .O(n6291) );
  NAND_GATE U6857 ( .I1(n6293), .I2(n6291), .O(n6289) );
  INV_GATE U6858 ( .I1(n5863), .O(n5872) );
  NAND_GATE U6859 ( .I1(n5872), .I2(n5868), .O(n5866) );
  NAND3_GATE U6860 ( .I1(n5866), .I2(n5865), .I3(n5864), .O(n5870) );
  OR_GATE U6861 ( .I1(n5868), .I2(n5867), .O(n5869) );
  NAND_GATE U6862 ( .I1(n5870), .I2(n5869), .O(n5873) );
  INV_GATE U6863 ( .I1(n6688), .O(n6691) );
  NAND_GATE U6864 ( .I1(B[19]), .I2(A[29]), .O(n6697) );
  INV_GATE U6865 ( .I1(n6697), .O(n6689) );
  NAND_GATE U6866 ( .I1(n6691), .I2(n6689), .O(n6686) );
  NAND_GATE U6867 ( .I1(n5873), .I2(n6697), .O(n6278) );
  NAND_GATE U6868 ( .I1(n402), .I2(n6697), .O(n6277) );
  OR_GATE U6869 ( .I1(n5874), .I2(n5879), .O(n5877) );
  OR_GATE U6870 ( .I1(n5878), .I2(n5875), .O(n5876) );
  AND_GATE U6871 ( .I1(n5877), .I2(n5876), .O(n5884) );
  NAND_GATE U6872 ( .I1(n5879), .I2(n1159), .O(n5881) );
  NAND3_GATE U6873 ( .I1(n5882), .I2(n5881), .I3(n5880), .O(n5883) );
  NAND_GATE U6874 ( .I1(n5884), .I2(n5883), .O(n6300) );
  INV_GATE U6875 ( .I1(n6300), .O(n6303) );
  NAND_GATE U6876 ( .I1(B[19]), .I2(A[28]), .O(n6307) );
  INV_GATE U6877 ( .I1(n6307), .O(n6301) );
  NAND_GATE U6878 ( .I1(n6303), .I2(n6301), .O(n6298) );
  OR_GATE U6879 ( .I1(n5885), .I2(n5890), .O(n5888) );
  OR_GATE U6880 ( .I1(n5889), .I2(n5886), .O(n5887) );
  AND_GATE U6881 ( .I1(n5888), .I2(n5887), .O(n5895) );
  NAND_GATE U6882 ( .I1(n5890), .I2(n1139), .O(n5892) );
  NAND3_GATE U6883 ( .I1(n5893), .I2(n5892), .I3(n5891), .O(n5894) );
  NAND_GATE U6884 ( .I1(n5895), .I2(n5894), .O(n6671) );
  INV_GATE U6885 ( .I1(n6671), .O(n6674) );
  NAND_GATE U6886 ( .I1(B[19]), .I2(A[27]), .O(n6678) );
  INV_GATE U6887 ( .I1(n6678), .O(n6672) );
  NAND_GATE U6888 ( .I1(n6674), .I2(n6672), .O(n6669) );
  OR_GATE U6889 ( .I1(n5896), .I2(n5901), .O(n5899) );
  OR_GATE U6890 ( .I1(n5900), .I2(n5897), .O(n5898) );
  AND_GATE U6891 ( .I1(n5899), .I2(n5898), .O(n5906) );
  NAND_GATE U6892 ( .I1(n5901), .I2(n1140), .O(n5903) );
  NAND3_GATE U6893 ( .I1(n5904), .I2(n5903), .I3(n5902), .O(n5905) );
  NAND_GATE U6894 ( .I1(n5906), .I2(n5905), .O(n6655) );
  INV_GATE U6895 ( .I1(n6655), .O(n6658) );
  NAND_GATE U6896 ( .I1(B[19]), .I2(A[26]), .O(n6662) );
  INV_GATE U6897 ( .I1(n6662), .O(n6656) );
  NAND_GATE U6898 ( .I1(n6658), .I2(n6656), .O(n6653) );
  OR_GATE U6899 ( .I1(n5907), .I2(n5912), .O(n5910) );
  OR_GATE U6900 ( .I1(n5911), .I2(n5908), .O(n5909) );
  AND_GATE U6901 ( .I1(n5910), .I2(n5909), .O(n5917) );
  NAND_GATE U6902 ( .I1(n1141), .I2(n5911), .O(n5915) );
  NAND3_GATE U6903 ( .I1(n5915), .I2(n5914), .I3(n5913), .O(n5916) );
  NAND_GATE U6904 ( .I1(B[19]), .I2(A[25]), .O(n6646) );
  INV_GATE U6905 ( .I1(n6646), .O(n6641) );
  NAND_GATE U6906 ( .I1(n713), .I2(n6641), .O(n6638) );
  OR_GATE U6907 ( .I1(n5918), .I2(n5923), .O(n5921) );
  OR_GATE U6908 ( .I1(n5922), .I2(n5919), .O(n5920) );
  NAND_GATE U6909 ( .I1(n1142), .I2(n5922), .O(n5926) );
  NAND3_GATE U6910 ( .I1(n5926), .I2(n5925), .I3(n5924), .O(n5927) );
  NAND_GATE U6911 ( .I1(B[19]), .I2(A[24]), .O(n6632) );
  INV_GATE U6912 ( .I1(n6632), .O(n6627) );
  NAND_GATE U6913 ( .I1(n750), .I2(n6627), .O(n6624) );
  OR_GATE U6914 ( .I1(n5928), .I2(n5934), .O(n5931) );
  OR_GATE U6915 ( .I1(n5933), .I2(n5929), .O(n5930) );
  AND_GATE U6916 ( .I1(n5931), .I2(n5930), .O(n5939) );
  INV_GATE U6917 ( .I1(n5934), .O(n5932) );
  NAND_GATE U6918 ( .I1(n5932), .I2(n5933), .O(n5937) );
  NAND3_GATE U6919 ( .I1(n5937), .I2(n5936), .I3(n5935), .O(n5938) );
  NAND_GATE U6920 ( .I1(B[19]), .I2(A[23]), .O(n6617) );
  INV_GATE U6921 ( .I1(n6617), .O(n6612) );
  NAND_GATE U6922 ( .I1(n797), .I2(n6612), .O(n6609) );
  OR_GATE U6923 ( .I1(n5940), .I2(n5944), .O(n5943) );
  OR_GATE U6924 ( .I1(n5945), .I2(n5941), .O(n5942) );
  AND_GATE U6925 ( .I1(n5943), .I2(n5942), .O(n5950) );
  NAND_GATE U6926 ( .I1(n5944), .I2(n1118), .O(n5948) );
  NAND3_GATE U6927 ( .I1(n5948), .I2(n5947), .I3(n5946), .O(n5949) );
  NAND_GATE U6928 ( .I1(B[19]), .I2(A[22]), .O(n6602) );
  INV_GATE U6929 ( .I1(n6602), .O(n6597) );
  NAND_GATE U6930 ( .I1(n939), .I2(n6597), .O(n6594) );
  OR_GATE U6931 ( .I1(n5951), .I2(n5956), .O(n5954) );
  OR_GATE U6932 ( .I1(n5955), .I2(n5952), .O(n5953) );
  AND_GATE U6933 ( .I1(n5954), .I2(n5953), .O(n5961) );
  NAND_GATE U6934 ( .I1(n700), .I2(n5955), .O(n5959) );
  NAND3_GATE U6935 ( .I1(n5959), .I2(n5958), .I3(n5957), .O(n5960) );
  NAND_GATE U6936 ( .I1(n5961), .I2(n5960), .O(n6583) );
  NAND_GATE U6937 ( .I1(B[19]), .I2(A[21]), .O(n6589) );
  INV_GATE U6938 ( .I1(n6589), .O(n6584) );
  NAND_GATE U6939 ( .I1(n834), .I2(n6584), .O(n6580) );
  NAND_GATE U6940 ( .I1(B[19]), .I2(A[20]), .O(n6573) );
  INV_GATE U6941 ( .I1(n6573), .O(n6567) );
  OR_GATE U6942 ( .I1(n5962), .I2(n5967), .O(n5965) );
  OR_GATE U6943 ( .I1(n5966), .I2(n5963), .O(n5964) );
  AND_GATE U6944 ( .I1(n5965), .I2(n5964), .O(n5972) );
  NAND_GATE U6945 ( .I1(n1100), .I2(n5966), .O(n5970) );
  NAND3_GATE U6946 ( .I1(n5970), .I2(n5969), .I3(n5968), .O(n5971) );
  NAND_GATE U6947 ( .I1(n5972), .I2(n5971), .O(n6558) );
  NAND_GATE U6948 ( .I1(B[19]), .I2(A[19]), .O(n6559) );
  INV_GATE U6949 ( .I1(n6559), .O(n6556) );
  NAND_GATE U6950 ( .I1(n347), .I2(n6556), .O(n6553) );
  NAND_GATE U6951 ( .I1(B[19]), .I2(A[18]), .O(n6315) );
  OR_GATE U6952 ( .I1(n5973), .I2(n5979), .O(n5976) );
  OR_GATE U6953 ( .I1(n5978), .I2(n5974), .O(n5975) );
  AND_GATE U6954 ( .I1(n5976), .I2(n5975), .O(n5984) );
  INV_GATE U6955 ( .I1(n5979), .O(n5977) );
  NAND_GATE U6956 ( .I1(n5977), .I2(n5978), .O(n5981) );
  NAND_GATE U6957 ( .I1(n5979), .I2(n332), .O(n5980) );
  NAND3_GATE U6958 ( .I1(n5982), .I2(n5981), .I3(n5980), .O(n5983) );
  NAND_GATE U6959 ( .I1(n5984), .I2(n5983), .O(n6314) );
  NAND_GATE U6960 ( .I1(n510), .I2(n1382), .O(n6318) );
  NAND_GATE U6961 ( .I1(B[19]), .I2(A[17]), .O(n6328) );
  INV_GATE U6962 ( .I1(n6328), .O(n6324) );
  INV_GATE U6963 ( .I1(n5991), .O(n5989) );
  NAND3_GATE U6964 ( .I1(n5989), .I2(n5985), .I3(n5990), .O(n5988) );
  OR_GATE U6965 ( .I1(n5990), .I2(n5986), .O(n5987) );
  AND_GATE U6966 ( .I1(n5988), .I2(n5987), .O(n5996) );
  NAND_GATE U6967 ( .I1(n5989), .I2(n5990), .O(n5993) );
  NAND3_GATE U6968 ( .I1(n5994), .I2(n5993), .I3(n5992), .O(n5995) );
  NAND_GATE U6969 ( .I1(n5996), .I2(n5995), .O(n6325) );
  NAND_GATE U6970 ( .I1(B[19]), .I2(A[16]), .O(n7108) );
  INV_GATE U6971 ( .I1(n7108), .O(n6541) );
  NAND_GATE U6972 ( .I1(n5998), .I2(n5997), .O(n6005) );
  INV_GATE U6973 ( .I1(n5999), .O(n6000) );
  NAND_GATE U6974 ( .I1(n6001), .I2(n6000), .O(n6004) );
  NAND_GATE U6975 ( .I1(n6005), .I2(n6004), .O(n6002) );
  NAND_GATE U6976 ( .I1(n6009), .I2(n6002), .O(n6007) );
  INV_GATE U6977 ( .I1(n6009), .O(n6003) );
  NAND3_GATE U6978 ( .I1(n6005), .I2(n6004), .I3(n6003), .O(n6006) );
  NAND3_GATE U6979 ( .I1(n6008), .I2(n6007), .I3(n6006), .O(n6015) );
  OR_GATE U6980 ( .I1(n6010), .I2(n6009), .O(n6014) );
  OR_GATE U6981 ( .I1(n6012), .I2(n6011), .O(n6013) );
  NAND3_GATE U6982 ( .I1(n6015), .I2(n6014), .I3(n6013), .O(n6543) );
  NAND_GATE U6983 ( .I1(n6541), .I2(n310), .O(n6540) );
  NAND_GATE U6984 ( .I1(B[19]), .I2(A[15]), .O(n6876) );
  INV_GATE U6985 ( .I1(n6876), .O(n6340) );
  OR_GATE U6986 ( .I1(n6018), .I2(n6017), .O(n6019) );
  INV_GATE U6987 ( .I1(n6029), .O(n6025) );
  NAND_GATE U6988 ( .I1(n6024), .I2(n6023), .O(n6027) );
  NAND3_GATE U6989 ( .I1(n6026), .I2(n6025), .I3(n6027), .O(n6032) );
  NAND_GATE U6990 ( .I1(n6027), .I2(n6026), .O(n6028) );
  NAND_GATE U6991 ( .I1(n6029), .I2(n6028), .O(n6031) );
  NAND3_GATE U6992 ( .I1(n6032), .I2(n6031), .I3(n6030), .O(n6033) );
  INV_GATE U6993 ( .I1(n6339), .O(n6341) );
  NAND_GATE U6994 ( .I1(n6340), .I2(n6341), .O(n6239) );
  NAND_GATE U6995 ( .I1(B[19]), .I2(A[14]), .O(n6533) );
  INV_GATE U6996 ( .I1(n6533), .O(n6525) );
  NAND3_GATE U6997 ( .I1(n6036), .I2(n6043), .I3(n706), .O(n6040) );
  NAND_GATE U6998 ( .I1(n6036), .I2(n6043), .O(n6037) );
  NAND_GATE U6999 ( .I1(n6041), .I2(n6037), .O(n6039) );
  NAND3_GATE U7000 ( .I1(n6040), .I2(n6039), .I3(n6038), .O(n6051) );
  OR_GATE U7001 ( .I1(n6042), .I2(n6041), .O(n6050) );
  NAND_GATE U7002 ( .I1(n6044), .I2(n6043), .O(n6048) );
  INV_GATE U7003 ( .I1(n6045), .O(n6047) );
  NAND3_GATE U7004 ( .I1(n6048), .I2(n6047), .I3(n6046), .O(n6049) );
  NAND3_GATE U7005 ( .I1(n6051), .I2(n6050), .I3(n6049), .O(n6529) );
  NAND_GATE U7006 ( .I1(n6525), .I2(n6527), .O(n6236) );
  NAND_GATE U7007 ( .I1(B[19]), .I2(A[13]), .O(n6346) );
  INV_GATE U7008 ( .I1(n6346), .O(n6351) );
  NAND_GATE U7009 ( .I1(n6057), .I2(n1285), .O(n6053) );
  NAND_GATE U7010 ( .I1(n6054), .I2(n6053), .O(n6060) );
  NAND_GATE U7011 ( .I1(n355), .I2(n6055), .O(n6059) );
  NAND3_GATE U7012 ( .I1(n6057), .I2(n1285), .I3(n6056), .O(n6058) );
  NAND3_GATE U7013 ( .I1(n6060), .I2(n6059), .I3(n6058), .O(n6345) );
  NAND_GATE U7014 ( .I1(n6344), .I2(n6345), .O(n6350) );
  NAND_GATE U7015 ( .I1(n6351), .I2(n6350), .O(n6233) );
  NAND_GATE U7016 ( .I1(B[19]), .I2(A[12]), .O(n6913) );
  INV_GATE U7017 ( .I1(n6913), .O(n6356) );
  NAND_GATE U7018 ( .I1(n6062), .I2(n6061), .O(n6066) );
  INV_GATE U7019 ( .I1(n6075), .O(n6065) );
  NAND3_GATE U7020 ( .I1(n6066), .I2(n6065), .I3(n6067), .O(n6071) );
  NAND_GATE U7021 ( .I1(n6067), .I2(n6066), .O(n6068) );
  NAND_GATE U7022 ( .I1(n6075), .I2(n6068), .O(n6070) );
  NAND3_GATE U7023 ( .I1(n6071), .I2(n6070), .I3(n6069), .O(n6078) );
  OR_GATE U7024 ( .I1(n6073), .I2(n6072), .O(n6077) );
  OR_GATE U7025 ( .I1(n6075), .I2(n6074), .O(n6076) );
  NAND3_GATE U7026 ( .I1(n6078), .I2(n6077), .I3(n6076), .O(n6359) );
  NAND_GATE U7027 ( .I1(n6356), .I2(n878), .O(n6231) );
  NAND_GATE U7028 ( .I1(B[19]), .I2(A[11]), .O(n6373) );
  INV_GATE U7029 ( .I1(n6373), .O(n6227) );
  NAND_GATE U7030 ( .I1(B[19]), .I2(A[10]), .O(n6925) );
  INV_GATE U7031 ( .I1(n6925), .O(n6509) );
  NAND_GATE U7032 ( .I1(B[19]), .I2(A[9]), .O(n6381) );
  INV_GATE U7033 ( .I1(n6381), .O(n6384) );
  NAND_GATE U7034 ( .I1(B[19]), .I2(A[7]), .O(n6400) );
  INV_GATE U7035 ( .I1(n6400), .O(n6164) );
  INV_GATE U7036 ( .I1(n6079), .O(n6080) );
  NAND_GATE U7037 ( .I1(n6081), .I2(n6080), .O(n6090) );
  NAND_GATE U7038 ( .I1(n6085), .I2(n6084), .O(n6086) );
  NAND_GATE U7039 ( .I1(n5577), .I2(n6086), .O(n6087) );
  NAND_GATE U7040 ( .I1(n6088), .I2(n6087), .O(n6089) );
  NAND3_GATE U7041 ( .I1(n6090), .I2(n6089), .I3(n867), .O(n6095) );
  NAND_GATE U7042 ( .I1(n6090), .I2(n6089), .O(n6091) );
  NAND_GATE U7043 ( .I1(n6092), .I2(n6091), .O(n6094) );
  NAND3_GATE U7044 ( .I1(n6095), .I2(n6094), .I3(n6093), .O(n6101) );
  NAND3_GATE U7045 ( .I1(n867), .I2(n6096), .I3(n6098), .O(n6100) );
  OR_GATE U7046 ( .I1(n6098), .I2(n6097), .O(n6099) );
  NAND_GATE U7047 ( .I1(B[19]), .I2(A[6]), .O(n6481) );
  INV_GATE U7048 ( .I1(n6481), .O(n6486) );
  NAND_GATE U7049 ( .I1(n1291), .I2(n6486), .O(n6479) );
  NAND_GATE U7050 ( .I1(B[19]), .I2(A[4]), .O(n6468) );
  INV_GATE U7051 ( .I1(n6468), .O(n6461) );
  NAND_GATE U7052 ( .I1(n1232), .I2(n6108), .O(n6102) );
  NAND3_GATE U7053 ( .I1(n6104), .I2(n6103), .I3(n6102), .O(n6111) );
  OR_GATE U7054 ( .I1(n6106), .I2(n6105), .O(n6110) );
  OR_GATE U7055 ( .I1(n6108), .I2(n6107), .O(n6109) );
  NAND3_GATE U7056 ( .I1(n6111), .I2(n6110), .I3(n6109), .O(n6464) );
  INV_GATE U7057 ( .I1(n6464), .O(n6462) );
  NAND_GATE U7058 ( .I1(n6461), .I2(n6462), .O(n6471) );
  NAND_GATE U7059 ( .I1(B[19]), .I2(A[3]), .O(n6430) );
  INV_GATE U7060 ( .I1(n6430), .O(n6132) );
  NAND_GATE U7061 ( .I1(B[19]), .I2(A[2]), .O(n6452) );
  INV_GATE U7062 ( .I1(n6452), .O(n6446) );
  NAND_GATE U7063 ( .I1(n1432), .I2(A[0]), .O(n6112) );
  NAND_GATE U7064 ( .I1(n14241), .I2(n6112), .O(n6113) );
  NAND_GATE U7065 ( .I1(B[21]), .I2(n6113), .O(n6117) );
  NAND_GATE U7066 ( .I1(n1433), .I2(A[1]), .O(n6114) );
  NAND_GATE U7067 ( .I1(n724), .I2(n6114), .O(n6115) );
  NAND_GATE U7068 ( .I1(B[20]), .I2(n6115), .O(n6116) );
  NAND_GATE U7069 ( .I1(n6117), .I2(n6116), .O(n6448) );
  NAND_GATE U7070 ( .I1(n6446), .I2(n6448), .O(n6443) );
  NAND3_GATE U7071 ( .I1(B[19]), .I2(B[20]), .I3(n1254), .O(n6444) );
  INV_GATE U7072 ( .I1(n6444), .O(n6447) );
  INV_GATE U7073 ( .I1(n6448), .O(n6445) );
  NAND_GATE U7074 ( .I1(n6452), .I2(n6445), .O(n6118) );
  NAND_GATE U7075 ( .I1(n6447), .I2(n6118), .O(n6119) );
  NAND_GATE U7076 ( .I1(n6443), .I2(n6119), .O(n6429) );
  NAND_GATE U7077 ( .I1(n6132), .I2(n6429), .O(n6425) );
  OR_GATE U7078 ( .I1(n6125), .I2(n6120), .O(n6131) );
  NAND_GATE U7079 ( .I1(n1370), .I2(n6125), .O(n6121) );
  NAND_GATE U7080 ( .I1(n6122), .I2(n6121), .O(n6129) );
  NAND_GATE U7081 ( .I1(n6124), .I2(n6123), .O(n6128) );
  NAND3_GATE U7082 ( .I1(n1370), .I2(n6126), .I3(n6125), .O(n6127) );
  NAND3_GATE U7083 ( .I1(n6129), .I2(n6128), .I3(n6127), .O(n6130) );
  NAND_GATE U7084 ( .I1(n6131), .I2(n6130), .O(n6428) );
  NAND_GATE U7085 ( .I1(n6429), .I2(n6428), .O(n6133) );
  NAND_GATE U7086 ( .I1(n6132), .I2(n6428), .O(n6424) );
  NAND3_GATE U7087 ( .I1(n6425), .I2(n6133), .I3(n6424), .O(n6472) );
  NAND_GATE U7088 ( .I1(n6468), .I2(n6464), .O(n6134) );
  NAND_GATE U7089 ( .I1(n6472), .I2(n6134), .O(n6135) );
  NAND_GATE U7090 ( .I1(n6471), .I2(n6135), .O(n6418) );
  INV_GATE U7091 ( .I1(n6148), .O(n6137) );
  NAND_GATE U7092 ( .I1(n6418), .I2(n6137), .O(n6151) );
  NAND_GATE U7093 ( .I1(n6139), .I2(n6143), .O(n6140) );
  NAND_GATE U7094 ( .I1(n6141), .I2(n6140), .O(n6146) );
  NAND_GATE U7095 ( .I1(n6142), .I2(n1304), .O(n6143) );
  NAND_GATE U7096 ( .I1(n6144), .I2(n6143), .O(n6145) );
  NAND3_GATE U7097 ( .I1(n6146), .I2(n6418), .I3(n6145), .O(n6150) );
  NAND_GATE U7098 ( .I1(B[19]), .I2(A[5]), .O(n6421) );
  INV_GATE U7099 ( .I1(n6421), .O(n6415) );
  NAND_GATE U7100 ( .I1(n6415), .I2(n6418), .O(n6414) );
  NAND_GATE U7101 ( .I1(n6146), .I2(n6145), .O(n6147) );
  NAND_GATE U7102 ( .I1(n6148), .I2(n6147), .O(n6419) );
  NAND_GATE U7103 ( .I1(n6415), .I2(n6419), .O(n6149) );
  NAND4_GATE U7104 ( .I1(n6151), .I2(n6150), .I3(n6414), .I4(n6149), .O(n6482)
         );
  NAND_GATE U7105 ( .I1(n6484), .I2(n6481), .O(n6152) );
  NAND_GATE U7106 ( .I1(n6482), .I2(n6152), .O(n6398) );
  NAND_GATE U7107 ( .I1(n6479), .I2(n6398), .O(n6407) );
  NAND_GATE U7108 ( .I1(n6164), .I2(n6407), .O(n6409) );
  INV_GATE U7109 ( .I1(n6155), .O(n6157) );
  NAND3_GATE U7110 ( .I1(n6156), .I2(n6157), .I3(n6158), .O(n6161) );
  NAND3_GATE U7111 ( .I1(n6156), .I2(n6155), .I3(n6154), .O(n6160) );
  NAND_GATE U7112 ( .I1(n6158), .I2(n6157), .O(n6162) );
  NAND_GATE U7113 ( .I1(n6163), .I2(n6162), .O(n6399) );
  NAND_GATE U7114 ( .I1(n6166), .I2(n6399), .O(n6159) );
  NAND_GATE U7115 ( .I1(n6396), .I2(n6159), .O(n6410) );
  NAND_GATE U7116 ( .I1(n6407), .I2(n6410), .O(n6167) );
  AND_GATE U7117 ( .I1(n6161), .I2(n6160), .O(n6166) );
  NAND3_GATE U7118 ( .I1(n6163), .I2(n6162), .I3(n6396), .O(n6165) );
  NAND3_GATE U7119 ( .I1(n6166), .I2(n6165), .I3(n6164), .O(n6408) );
  NAND3_GATE U7120 ( .I1(n6409), .I2(n6167), .I3(n6408), .O(n6944) );
  NAND_GATE U7121 ( .I1(B[19]), .I2(A[8]), .O(n6949) );
  NAND_GATE U7122 ( .I1(n6168), .I2(n6172), .O(n6176) );
  NAND4_GATE U7123 ( .I1(n6172), .I2(n6171), .I3(n6170), .I4(n6169), .O(n6175)
         );
  NAND4_GATE U7124 ( .I1(n6176), .I2(n6175), .I3(n6174), .I4(n6173), .O(n6177)
         );
  NAND_GATE U7125 ( .I1(n6178), .I2(n6177), .O(n6185) );
  INV_GATE U7126 ( .I1(n6179), .O(n6183) );
  NAND_GATE U7127 ( .I1(n6183), .I2(n6185), .O(n6180) );
  NAND3_GATE U7128 ( .I1(n6182), .I2(n6181), .I3(n6180), .O(n6188) );
  NAND3_GATE U7129 ( .I1(n1209), .I2(n6183), .I3(n1258), .O(n6187) );
  OR_GATE U7130 ( .I1(n6185), .I2(n6184), .O(n6186) );
  NAND3_GATE U7131 ( .I1(n6188), .I2(n6187), .I3(n6186), .O(n6945) );
  NAND_GATE U7132 ( .I1(n6949), .I2(n6945), .O(n6189) );
  NAND_GATE U7133 ( .I1(n6944), .I2(n6189), .O(n6191) );
  INV_GATE U7134 ( .I1(n6949), .O(n6497) );
  INV_GATE U7135 ( .I1(n6945), .O(n6943) );
  NAND_GATE U7136 ( .I1(n6497), .I2(n6943), .O(n6190) );
  NAND_GATE U7137 ( .I1(n6191), .I2(n6190), .O(n6378) );
  NAND_GATE U7138 ( .I1(n6384), .I2(n6378), .O(n6391) );
  NAND_GATE U7139 ( .I1(n6193), .I2(n7), .O(n6194) );
  NAND3_GATE U7140 ( .I1(n6196), .I2(n6195), .I3(n6194), .O(n6386) );
  NAND3_GATE U7141 ( .I1(n6198), .I2(n7), .I3(n6197), .O(n6385) );
  NAND_GATE U7142 ( .I1(n6200), .I2(n6199), .O(n6383) );
  NAND3_GATE U7143 ( .I1(n6386), .I2(n6385), .I3(n6383), .O(n6377) );
  NAND_GATE U7144 ( .I1(n6382), .I2(n6377), .O(n6392) );
  NAND_GATE U7145 ( .I1(n6378), .I2(n6392), .O(n6202) );
  NAND_GATE U7146 ( .I1(n6384), .I2(n6392), .O(n6201) );
  NAND3_GATE U7147 ( .I1(n6391), .I2(n6202), .I3(n6201), .O(n6513) );
  NAND_GATE U7148 ( .I1(n6509), .I2(n6513), .O(n6506) );
  NAND3_GATE U7149 ( .I1(n765), .I2(n6205), .I3(n1384), .O(n6215) );
  NAND3_GATE U7150 ( .I1(n765), .I2(n6209), .I3(n6208), .O(n6213) );
  NAND_GATE U7151 ( .I1(n6209), .I2(n6208), .O(n6210) );
  NAND_GATE U7152 ( .I1(n6211), .I2(n6210), .O(n6212) );
  NAND3_GATE U7153 ( .I1(n6214), .I2(n6213), .I3(n6212), .O(n6216) );
  NAND3_GATE U7154 ( .I1(n6217), .I2(n6215), .I3(n6216), .O(n6510) );
  INV_GATE U7155 ( .I1(n6510), .O(n6512) );
  NAND_GATE U7156 ( .I1(n6509), .I2(n6512), .O(n6219) );
  NAND4_GATE U7157 ( .I1(n6217), .I2(n6216), .I3(n6513), .I4(n6215), .O(n6218)
         );
  NAND3_GATE U7158 ( .I1(n6506), .I2(n6219), .I3(n6218), .O(n6372) );
  NAND_GATE U7159 ( .I1(n6227), .I2(n6372), .O(n6362) );
  NAND3_GATE U7160 ( .I1(n6220), .I2(n5), .I3(n6222), .O(n6367) );
  NAND_GATE U7161 ( .I1(n6220), .I2(n6224), .O(n6366) );
  NAND_GATE U7162 ( .I1(n6221), .I2(n796), .O(n6224) );
  NAND_GATE U7163 ( .I1(n6224), .I2(n6223), .O(n6368) );
  NAND_GATE U7164 ( .I1(n6369), .I2(n6368), .O(n6225) );
  NAND_GATE U7165 ( .I1(n6366), .I2(n6225), .O(n6226) );
  NAND_GATE U7166 ( .I1(n6367), .I2(n6226), .O(n6363) );
  NAND_GATE U7167 ( .I1(n6227), .I2(n6363), .O(n6361) );
  NAND_GATE U7168 ( .I1(n6372), .I2(n6363), .O(n6228) );
  NAND3_GATE U7169 ( .I1(n6362), .I2(n6361), .I3(n6228), .O(n6357) );
  NAND_GATE U7170 ( .I1(n6913), .I2(n6359), .O(n6229) );
  NAND_GATE U7171 ( .I1(n6357), .I2(n6229), .O(n6230) );
  NAND_GATE U7172 ( .I1(n6231), .I2(n6230), .O(n6343) );
  NAND_GATE U7173 ( .I1(n6350), .I2(n6343), .O(n6232) );
  NAND_GATE U7174 ( .I1(n6351), .I2(n6343), .O(n6349) );
  NAND3_GATE U7175 ( .I1(n6233), .I2(n6232), .I3(n6349), .O(n6526) );
  NAND_GATE U7176 ( .I1(n6533), .I2(n6529), .O(n6234) );
  NAND_GATE U7177 ( .I1(n6526), .I2(n6234), .O(n6235) );
  NAND_GATE U7178 ( .I1(n6236), .I2(n6235), .O(n6342) );
  NAND_GATE U7179 ( .I1(n6876), .I2(n6339), .O(n6237) );
  NAND_GATE U7180 ( .I1(n6342), .I2(n6237), .O(n6238) );
  NAND_GATE U7181 ( .I1(n7108), .I2(n6543), .O(n6240) );
  NAND_GATE U7182 ( .I1(n6542), .I2(n6240), .O(n6241) );
  NAND_GATE U7183 ( .I1(n6328), .I2(n6325), .O(n6242) );
  NAND_GATE U7184 ( .I1(n6332), .I2(n6242), .O(n6243) );
  NAND_GATE U7185 ( .I1(n6331), .I2(n6243), .O(n6319) );
  NAND_GATE U7186 ( .I1(n6315), .I2(n6314), .O(n6244) );
  NAND_GATE U7187 ( .I1(n6319), .I2(n6244), .O(n6245) );
  NAND_GATE U7188 ( .I1(n6318), .I2(n6245), .O(n6557) );
  NAND_GATE U7189 ( .I1(n6558), .I2(n6559), .O(n6246) );
  NAND_GATE U7190 ( .I1(n6557), .I2(n6246), .O(n6247) );
  NAND_GATE U7191 ( .I1(n6567), .I2(n327), .O(n6566) );
  OR_GATE U7192 ( .I1(n6252), .I2(n6249), .O(n6250) );
  AND_GATE U7193 ( .I1(n6251), .I2(n6250), .O(n6258) );
  NAND_GATE U7194 ( .I1(n180), .I2(n6252), .O(n6256) );
  NAND3_GATE U7195 ( .I1(n6256), .I2(n6255), .I3(n6254), .O(n6257) );
  NAND_GATE U7196 ( .I1(n6258), .I2(n6257), .O(n6569) );
  INV_GATE U7197 ( .I1(n6569), .O(n6568) );
  NAND_GATE U7198 ( .I1(n6573), .I2(n827), .O(n6259) );
  NAND_GATE U7199 ( .I1(n6568), .I2(n6259), .O(n6260) );
  NAND_GATE U7200 ( .I1(n6566), .I2(n6260), .O(n6585) );
  NAND_GATE U7201 ( .I1(n6583), .I2(n6589), .O(n6261) );
  NAND_GATE U7202 ( .I1(n6585), .I2(n6261), .O(n6262) );
  NAND_GATE U7203 ( .I1(n6580), .I2(n6262), .O(n6598) );
  NAND_GATE U7204 ( .I1(n6596), .I2(n6602), .O(n6263) );
  NAND_GATE U7205 ( .I1(n6598), .I2(n6263), .O(n6264) );
  NAND_GATE U7206 ( .I1(n6594), .I2(n6264), .O(n6613) );
  NAND_GATE U7207 ( .I1(n6611), .I2(n6617), .O(n6265) );
  NAND_GATE U7208 ( .I1(n6613), .I2(n6265), .O(n6266) );
  NAND_GATE U7209 ( .I1(n6609), .I2(n6266), .O(n6628) );
  NAND_GATE U7210 ( .I1(n6626), .I2(n6632), .O(n6267) );
  NAND_GATE U7211 ( .I1(n6628), .I2(n6267), .O(n6268) );
  NAND_GATE U7212 ( .I1(n6624), .I2(n6268), .O(n6642) );
  NAND_GATE U7213 ( .I1(n6640), .I2(n6646), .O(n6269) );
  NAND_GATE U7214 ( .I1(n6642), .I2(n6269), .O(n6270) );
  NAND_GATE U7215 ( .I1(n6638), .I2(n6270), .O(n6657) );
  NAND_GATE U7216 ( .I1(n6655), .I2(n6662), .O(n6271) );
  NAND_GATE U7217 ( .I1(n6657), .I2(n6271), .O(n6272) );
  NAND_GATE U7218 ( .I1(n6653), .I2(n6272), .O(n6673) );
  NAND_GATE U7219 ( .I1(n6671), .I2(n6678), .O(n6273) );
  NAND_GATE U7220 ( .I1(n6673), .I2(n6273), .O(n6274) );
  NAND_GATE U7221 ( .I1(n6669), .I2(n6274), .O(n6302) );
  NAND_GATE U7222 ( .I1(n6300), .I2(n6307), .O(n6275) );
  NAND_GATE U7223 ( .I1(n6302), .I2(n6275), .O(n6276) );
  NAND_GATE U7224 ( .I1(n6298), .I2(n6276), .O(n6690) );
  NAND3_GATE U7225 ( .I1(n6278), .I2(n6277), .I3(n6690), .O(n6279) );
  NAND_GATE U7226 ( .I1(n6686), .I2(n6279), .O(n6292) );
  NAND_GATE U7227 ( .I1(n6290), .I2(n6714), .O(n6280) );
  NAND_GATE U7228 ( .I1(n6292), .I2(n6280), .O(n6282) );
  NAND_GATE U7229 ( .I1(n1431), .I2(A[31]), .O(n6281) );
  NAND3_GATE U7230 ( .I1(n6289), .I2(n6282), .I3(n6281), .O(n6286) );
  NAND_GATE U7231 ( .I1(n403), .I2(n6286), .O(n6288) );
  NAND_GATE U7232 ( .I1(n14801), .I2(n6288), .O(n6285) );
  INV_GATE U7233 ( .I1(n6288), .O(n14800) );
  NAND_GATE U7234 ( .I1(n6283), .I2(n14800), .O(n6284) );
  NAND_GATE U7235 ( .I1(n6285), .I2(n6284), .O(\A1[49] ) );
  NAND_GATE U7236 ( .I1(n6288), .I2(n6287), .O(n6708) );
  INV_GATE U7237 ( .I1(n6708), .O(n14803) );
  NAND_GATE U7238 ( .I1(n6291), .I2(n6295), .O(n6711) );
  NAND_GATE U7239 ( .I1(n6293), .I2(n6292), .O(n6294) );
  NAND_GATE U7240 ( .I1(n6295), .I2(n6294), .O(n6713) );
  NAND_GATE U7241 ( .I1(n6714), .I2(n6713), .O(n6296) );
  NAND_GATE U7242 ( .I1(n6711), .I2(n6296), .O(n6297) );
  NAND_GATE U7243 ( .I1(n6712), .I2(n6297), .O(n6707) );
  NAND_GATE U7244 ( .I1(n1430), .I2(A[31]), .O(n6719) );
  INV_GATE U7245 ( .I1(n6298), .O(n6299) );
  NAND_GATE U7246 ( .I1(n6299), .I2(n6302), .O(n6311) );
  NAND_GATE U7247 ( .I1(n6301), .I2(n6305), .O(n6309) );
  NAND_GATE U7248 ( .I1(n6303), .I2(n6302), .O(n6304) );
  NAND_GATE U7249 ( .I1(n6305), .I2(n6304), .O(n6306) );
  NAND_GATE U7250 ( .I1(n6307), .I2(n6306), .O(n6308) );
  NAND_GATE U7251 ( .I1(n6309), .I2(n6308), .O(n6310) );
  NAND_GATE U7252 ( .I1(n6311), .I2(n6310), .O(n6740) );
  NAND_GATE U7253 ( .I1(B[18]), .I2(A[28]), .O(n6756) );
  INV_GATE U7254 ( .I1(n6756), .O(n6683) );
  NAND_GATE U7255 ( .I1(B[18]), .I2(A[27]), .O(n6767) );
  INV_GATE U7256 ( .I1(n6767), .O(n6667) );
  NAND_GATE U7257 ( .I1(B[18]), .I2(A[26]), .O(n6778) );
  INV_GATE U7258 ( .I1(n6778), .O(n6651) );
  NAND_GATE U7259 ( .I1(B[18]), .I2(A[25]), .O(n6789) );
  INV_GATE U7260 ( .I1(n6789), .O(n6636) );
  NAND_GATE U7261 ( .I1(B[18]), .I2(A[24]), .O(n6800) );
  INV_GATE U7262 ( .I1(n6800), .O(n6622) );
  NAND_GATE U7263 ( .I1(B[18]), .I2(A[23]), .O(n6810) );
  INV_GATE U7264 ( .I1(n6810), .O(n6607) );
  NAND_GATE U7265 ( .I1(B[18]), .I2(A[22]), .O(n6821) );
  INV_GATE U7266 ( .I1(n6821), .O(n6592) );
  NAND_GATE U7267 ( .I1(B[18]), .I2(A[21]), .O(n6832) );
  INV_GATE U7268 ( .I1(n6832), .O(n6578) );
  NAND_GATE U7269 ( .I1(B[18]), .I2(A[20]), .O(n6843) );
  INV_GATE U7270 ( .I1(n6843), .O(n6564) );
  NAND_GATE U7271 ( .I1(B[18]), .I2(A[19]), .O(n6852) );
  INV_GATE U7272 ( .I1(n6852), .O(n6551) );
  NAND_GATE U7273 ( .I1(n6314), .I2(n6313), .O(n6312) );
  NAND_GATE U7274 ( .I1(n510), .I2(n6312), .O(n6317) );
  NAND_GATE U7275 ( .I1(n6317), .I2(n6316), .O(n6322) );
  INV_GATE U7276 ( .I1(n6318), .O(n6320) );
  NAND_GATE U7277 ( .I1(n6320), .I2(n6319), .O(n6321) );
  NAND_GATE U7278 ( .I1(n6322), .I2(n6321), .O(n6849) );
  NAND_GATE U7279 ( .I1(n6551), .I2(n6849), .O(n6853) );
  NAND_GATE U7280 ( .I1(B[18]), .I2(A[18]), .O(n6860) );
  INV_GATE U7281 ( .I1(n6860), .O(n6549) );
  NAND_GATE U7282 ( .I1(n6325), .I2(n666), .O(n6323) );
  NAND_GATE U7283 ( .I1(n6324), .I2(n6323), .O(n6330) );
  NAND_GATE U7284 ( .I1(n6326), .I2(n6323), .O(n6327) );
  NAND_GATE U7285 ( .I1(n6328), .I2(n6327), .O(n6329) );
  NAND_GATE U7286 ( .I1(n6330), .I2(n6329), .O(n6335) );
  INV_GATE U7287 ( .I1(n6331), .O(n6333) );
  NAND_GATE U7288 ( .I1(n6333), .I2(n6332), .O(n6334) );
  NAND_GATE U7289 ( .I1(n6335), .I2(n6334), .O(n6861) );
  NAND_GATE U7290 ( .I1(n6549), .I2(n6861), .O(n6863) );
  NAND_GATE U7291 ( .I1(B[18]), .I2(A[17]), .O(n7115) );
  INV_GATE U7292 ( .I1(n7115), .O(n6547) );
  NAND_GATE U7293 ( .I1(n6341), .I2(n6342), .O(n6337) );
  INV_GATE U7294 ( .I1(n6342), .O(n6338) );
  NAND_GATE U7295 ( .I1(n6339), .I2(n6338), .O(n6336) );
  NAND_GATE U7296 ( .I1(n6337), .I2(n6336), .O(n6875) );
  NAND_GATE U7297 ( .I1(n6340), .I2(n6336), .O(n6870) );
  NAND3_GATE U7298 ( .I1(n6342), .I2(n6341), .I3(n6340), .O(n6872) );
  NAND_GATE U7299 ( .I1(B[18]), .I2(A[16]), .O(n6881) );
  INV_GATE U7300 ( .I1(n6881), .O(n6538) );
  NAND3_GATE U7301 ( .I1(n6869), .I2(n6879), .I3(n6538), .O(n6868) );
  NAND_GATE U7302 ( .I1(B[18]), .I2(A[15]), .O(n6892) );
  INV_GATE U7303 ( .I1(n6892), .O(n6889) );
  NAND_GATE U7304 ( .I1(B[18]), .I2(A[14]), .O(n7205) );
  INV_GATE U7305 ( .I1(n7205), .O(n6904) );
  NAND_GATE U7306 ( .I1(n6350), .I2(n879), .O(n6348) );
  NAND3_GATE U7307 ( .I1(n6345), .I2(n6344), .I3(n6343), .O(n6347) );
  NAND3_GATE U7308 ( .I1(n6348), .I2(n6347), .I3(n6346), .O(n6354) );
  OR_GATE U7309 ( .I1(n6349), .I2(n6350), .O(n6353) );
  NAND3_GATE U7310 ( .I1(n879), .I2(n6351), .I3(n6350), .O(n6352) );
  NAND3_GATE U7311 ( .I1(n6354), .I2(n6353), .I3(n6352), .O(n6899) );
  NAND_GATE U7312 ( .I1(n6904), .I2(n6902), .O(n6524) );
  NAND_GATE U7313 ( .I1(B[18]), .I2(A[13]), .O(n6917) );
  INV_GATE U7314 ( .I1(n6917), .O(n6521) );
  INV_GATE U7315 ( .I1(n6357), .O(n6358) );
  NAND_GATE U7316 ( .I1(n6359), .I2(n6358), .O(n6355) );
  NAND_GATE U7317 ( .I1(n6356), .I2(n6355), .O(n6906) );
  NAND3_GATE U7318 ( .I1(n6356), .I2(n6357), .I3(n878), .O(n6907) );
  NAND_GATE U7319 ( .I1(n878), .I2(n6357), .O(n6360) );
  NAND_GATE U7320 ( .I1(n6360), .I2(n6355), .O(n6912) );
  NAND_GATE U7321 ( .I1(n6913), .I2(n6912), .O(n6520) );
  NAND3_GATE U7322 ( .I1(n6521), .I2(n6914), .I3(n6520), .O(n6909) );
  NAND_GATE U7323 ( .I1(B[18]), .I2(A[12]), .O(n7081) );
  INV_GATE U7324 ( .I1(n7081), .O(n7088) );
  OR_GATE U7325 ( .I1(n6361), .I2(n6372), .O(n6365) );
  OR_GATE U7326 ( .I1(n6363), .I2(n6362), .O(n6364) );
  NAND_GATE U7327 ( .I1(n6370), .I2(n6225), .O(n6371) );
  NAND_GATE U7328 ( .I1(n6372), .I2(n6371), .O(n6374) );
  NAND3_GATE U7329 ( .I1(n6375), .I2(n6374), .I3(n6373), .O(n6376) );
  INV_GATE U7330 ( .I1(n7083), .O(n7080) );
  NAND_GATE U7331 ( .I1(n7088), .I2(n7080), .O(n6519) );
  NAND_GATE U7332 ( .I1(B[18]), .I2(A[11]), .O(n6933) );
  INV_GATE U7333 ( .I1(n6933), .O(n6515) );
  NAND_GATE U7334 ( .I1(B[18]), .I2(A[10]), .O(n7245) );
  INV_GATE U7335 ( .I1(n7245), .O(n7066) );
  INV_GATE U7336 ( .I1(n6378), .O(n6390) );
  NAND_GATE U7337 ( .I1(n6390), .I2(n6392), .O(n6380) );
  NAND3_GATE U7338 ( .I1(n6382), .I2(n6378), .I3(n6377), .O(n6379) );
  NAND3_GATE U7339 ( .I1(n6380), .I2(n6379), .I3(n6381), .O(n6395) );
  OR_GATE U7340 ( .I1(n6382), .I2(n6381), .O(n6388) );
  NAND4_GATE U7341 ( .I1(n6386), .I2(n6385), .I3(n6384), .I4(n6383), .O(n6387)
         );
  NAND_GATE U7342 ( .I1(n6388), .I2(n6387), .O(n6389) );
  NAND_GATE U7343 ( .I1(n6390), .I2(n6389), .O(n6394) );
  OR_GATE U7344 ( .I1(n6392), .I2(n6391), .O(n6393) );
  NAND3_GATE U7345 ( .I1(n6395), .I2(n6394), .I3(n6393), .O(n7068) );
  NAND_GATE U7346 ( .I1(n7066), .I2(n7070), .O(n6505) );
  NAND_GATE U7347 ( .I1(B[18]), .I2(A[9]), .O(n7061) );
  INV_GATE U7348 ( .I1(n7061), .O(n6939) );
  NAND_GATE U7349 ( .I1(B[18]), .I2(A[8]), .O(n7261) );
  INV_GATE U7350 ( .I1(n7261), .O(n7047) );
  INV_GATE U7351 ( .I1(n6396), .O(n6397) );
  NAND_GATE U7352 ( .I1(n6400), .I2(n6397), .O(n6403) );
  NAND3_GATE U7353 ( .I1(n6479), .I2(n6400), .I3(n6398), .O(n6402) );
  NAND3_GATE U7354 ( .I1(n6166), .I2(n6400), .I3(n6399), .O(n6401) );
  NAND3_GATE U7355 ( .I1(n6403), .I2(n6402), .I3(n6401), .O(n6406) );
  INV_GATE U7356 ( .I1(n6407), .O(n6404) );
  NAND_GATE U7357 ( .I1(n6404), .I2(n6410), .O(n6405) );
  NAND_GATE U7358 ( .I1(n6406), .I2(n6405), .O(n6413) );
  OR_GATE U7359 ( .I1(n6408), .I2(n6407), .O(n6412) );
  OR_GATE U7360 ( .I1(n6410), .I2(n6409), .O(n6411) );
  NAND3_GATE U7361 ( .I1(n6413), .I2(n6412), .I3(n6411), .O(n7049) );
  INV_GATE U7362 ( .I1(n7049), .O(n7051) );
  NAND_GATE U7363 ( .I1(n7047), .I2(n7051), .O(n6496) );
  OR_GATE U7364 ( .I1(n6419), .I2(n6414), .O(n6417) );
  INV_GATE U7365 ( .I1(n6418), .O(n6420) );
  NAND3_GATE U7366 ( .I1(n6420), .I2(n6415), .I3(n6419), .O(n6416) );
  AND_GATE U7367 ( .I1(n6417), .I2(n6416), .O(n7033) );
  NAND_GATE U7368 ( .I1(n6420), .I2(n6419), .O(n6422) );
  NAND3_GATE U7369 ( .I1(n6423), .I2(n6422), .I3(n6421), .O(n7032) );
  NAND_GATE U7370 ( .I1(n7033), .I2(n7032), .O(n7030) );
  NAND_GATE U7371 ( .I1(B[18]), .I2(A[6]), .O(n7031) );
  INV_GATE U7372 ( .I1(n7031), .O(n7034) );
  NAND_GATE U7373 ( .I1(B[18]), .I2(A[5]), .O(n6968) );
  INV_GATE U7374 ( .I1(n6968), .O(n6476) );
  OR_GATE U7375 ( .I1(n6424), .I2(n6429), .O(n6427) );
  OR_GATE U7376 ( .I1(n6428), .I2(n6425), .O(n6426) );
  AND_GATE U7377 ( .I1(n6427), .I2(n6426), .O(n6434) );
  NAND_GATE U7378 ( .I1(n1227), .I2(n6428), .O(n6432) );
  NAND3_GATE U7379 ( .I1(n6432), .I2(n6431), .I3(n6430), .O(n6433) );
  NAND_GATE U7380 ( .I1(n6434), .I2(n6433), .O(n7014) );
  INV_GATE U7381 ( .I1(n7014), .O(n7017) );
  NAND_GATE U7382 ( .I1(B[18]), .I2(A[4]), .O(n7021) );
  INV_GATE U7383 ( .I1(n7021), .O(n7015) );
  NAND_GATE U7384 ( .I1(n7017), .I2(n7015), .O(n7012) );
  NAND_GATE U7385 ( .I1(B[18]), .I2(A[3]), .O(n6983) );
  INV_GATE U7386 ( .I1(n6983), .O(n6457) );
  NAND_GATE U7387 ( .I1(B[18]), .I2(A[2]), .O(n7003) );
  INV_GATE U7388 ( .I1(n7003), .O(n6999) );
  NAND_GATE U7389 ( .I1(n1431), .I2(A[0]), .O(n6435) );
  NAND_GATE U7390 ( .I1(n14241), .I2(n6435), .O(n6436) );
  NAND_GATE U7391 ( .I1(B[20]), .I2(n6436), .O(n6440) );
  NAND_GATE U7392 ( .I1(n1432), .I2(A[1]), .O(n6437) );
  NAND_GATE U7393 ( .I1(n724), .I2(n6437), .O(n6438) );
  NAND_GATE U7394 ( .I1(B[19]), .I2(n6438), .O(n6439) );
  NAND_GATE U7395 ( .I1(n6440), .I2(n6439), .O(n7001) );
  NAND_GATE U7396 ( .I1(n6999), .I2(n7001), .O(n6996) );
  NAND3_GATE U7397 ( .I1(B[18]), .I2(B[19]), .I3(n1254), .O(n6997) );
  INV_GATE U7398 ( .I1(n6997), .O(n7000) );
  INV_GATE U7399 ( .I1(n7001), .O(n6998) );
  NAND_GATE U7400 ( .I1(n7003), .I2(n6998), .O(n6441) );
  NAND_GATE U7401 ( .I1(n7000), .I2(n6441), .O(n6442) );
  NAND_GATE U7402 ( .I1(n6996), .I2(n6442), .O(n6982) );
  NAND_GATE U7403 ( .I1(n6457), .I2(n6982), .O(n6977) );
  OR_GATE U7404 ( .I1(n6444), .I2(n6443), .O(n6456) );
  NAND_GATE U7405 ( .I1(n6446), .I2(n6450), .O(n6454) );
  NAND_GATE U7406 ( .I1(n6448), .I2(n6447), .O(n6449) );
  NAND_GATE U7407 ( .I1(n6450), .I2(n6449), .O(n6451) );
  NAND_GATE U7408 ( .I1(n6452), .I2(n6451), .O(n6453) );
  NAND_GATE U7409 ( .I1(n6454), .I2(n6453), .O(n6455) );
  NAND_GATE U7410 ( .I1(n6456), .I2(n6455), .O(n6981) );
  NAND_GATE U7411 ( .I1(n6982), .I2(n6981), .O(n6458) );
  NAND_GATE U7412 ( .I1(n6457), .I2(n6981), .O(n6976) );
  NAND_GATE U7413 ( .I1(n7014), .I2(n7021), .O(n6459) );
  NAND_GATE U7414 ( .I1(n7016), .I2(n6459), .O(n6460) );
  NAND_GATE U7415 ( .I1(n7012), .I2(n6460), .O(n6969) );
  NAND_GATE U7416 ( .I1(n6476), .I2(n6969), .O(n6971) );
  INV_GATE U7417 ( .I1(n6472), .O(n6463) );
  NAND_GATE U7418 ( .I1(n6461), .I2(n6465), .O(n6470) );
  NAND_GATE U7419 ( .I1(n6462), .I2(n6472), .O(n6466) );
  NAND_GATE U7420 ( .I1(n6464), .I2(n6463), .O(n6465) );
  NAND_GATE U7421 ( .I1(n6466), .I2(n6465), .O(n6467) );
  NAND_GATE U7422 ( .I1(n6468), .I2(n6467), .O(n6469) );
  NAND_GATE U7423 ( .I1(n6470), .I2(n6469), .O(n6475) );
  INV_GATE U7424 ( .I1(n6471), .O(n6473) );
  NAND_GATE U7425 ( .I1(n6473), .I2(n6472), .O(n6474) );
  NAND_GATE U7426 ( .I1(n6475), .I2(n6474), .O(n6972) );
  NAND_GATE U7427 ( .I1(n6969), .I2(n6972), .O(n6477) );
  NAND_GATE U7428 ( .I1(n6476), .I2(n6972), .O(n6970) );
  NAND3_GATE U7429 ( .I1(n6971), .I2(n6477), .I3(n6970), .O(n7039) );
  NAND_GATE U7430 ( .I1(n7030), .I2(n7031), .O(n6478) );
  INV_GATE U7431 ( .I1(n6479), .O(n6480) );
  NAND_GATE U7432 ( .I1(n6480), .I2(n6482), .O(n6491) );
  INV_GATE U7433 ( .I1(n6482), .O(n6483) );
  NAND3_GATE U7434 ( .I1(n6481), .I2(n6483), .I3(n6484), .O(n6489) );
  NAND_GATE U7435 ( .I1(n1291), .I2(n6482), .O(n6488) );
  NAND_GATE U7436 ( .I1(n6486), .I2(n6485), .O(n6487) );
  NAND3_GATE U7437 ( .I1(n6489), .I2(n6488), .I3(n6487), .O(n6490) );
  NAND_GATE U7438 ( .I1(n6491), .I2(n6490), .O(n6962) );
  NAND_GATE U7439 ( .I1(n6956), .I2(n6962), .O(n6493) );
  NAND_GATE U7440 ( .I1(B[18]), .I2(A[7]), .O(n6959) );
  INV_GATE U7441 ( .I1(n6959), .O(n6960) );
  NAND_GATE U7442 ( .I1(n6960), .I2(n6962), .O(n6492) );
  NAND_GATE U7443 ( .I1(n6960), .I2(n6956), .O(n6961) );
  NAND3_GATE U7444 ( .I1(n6493), .I2(n6492), .I3(n6961), .O(n7050) );
  NAND_GATE U7445 ( .I1(n7261), .I2(n7049), .O(n6494) );
  NAND_GATE U7446 ( .I1(n7050), .I2(n6494), .O(n6495) );
  NAND_GATE U7447 ( .I1(n6496), .I2(n6495), .O(n6951) );
  NAND_GATE U7448 ( .I1(n6939), .I2(n6951), .O(n6938) );
  NAND3_GATE U7449 ( .I1(n6944), .I2(n6497), .I3(n6943), .O(n6942) );
  NAND3_GATE U7450 ( .I1(n6949), .I2(n6945), .I3(n6946), .O(n6499) );
  NAND_GATE U7451 ( .I1(n6944), .I2(n6943), .O(n6498) );
  NAND_GATE U7452 ( .I1(n6497), .I2(n6947), .O(n6941) );
  NAND3_GATE U7453 ( .I1(n6499), .I2(n6498), .I3(n6941), .O(n6500) );
  NAND_GATE U7454 ( .I1(n6942), .I2(n6500), .O(n6940) );
  NAND_GATE U7455 ( .I1(n6951), .I2(n6940), .O(n6502) );
  NAND_GATE U7456 ( .I1(n6939), .I2(n6940), .O(n6501) );
  NAND3_GATE U7457 ( .I1(n6938), .I2(n6502), .I3(n6501), .O(n7069) );
  NAND_GATE U7458 ( .I1(n7245), .I2(n7068), .O(n6503) );
  NAND_GATE U7459 ( .I1(n7069), .I2(n6503), .O(n6504) );
  NAND_GATE U7460 ( .I1(n6505), .I2(n6504), .O(n6932) );
  NAND_GATE U7461 ( .I1(n6515), .I2(n6932), .O(n6921) );
  INV_GATE U7462 ( .I1(n6506), .O(n6507) );
  NAND_GATE U7463 ( .I1(n6507), .I2(n6512), .O(n6927) );
  INV_GATE U7464 ( .I1(n6513), .O(n6511) );
  NAND_GATE U7465 ( .I1(n6511), .I2(n6510), .O(n6508) );
  NAND_GATE U7466 ( .I1(n6509), .I2(n6508), .O(n6926) );
  NAND_GATE U7467 ( .I1(n6926), .I2(n6929), .O(n6514) );
  NAND_GATE U7468 ( .I1(n6927), .I2(n6514), .O(n6922) );
  NAND_GATE U7469 ( .I1(n6932), .I2(n6922), .O(n6516) );
  NAND_GATE U7470 ( .I1(n6515), .I2(n6922), .O(n6920) );
  NAND3_GATE U7471 ( .I1(n6921), .I2(n6516), .I3(n6920), .O(n7079) );
  NAND_GATE U7472 ( .I1(n7081), .I2(n7083), .O(n6517) );
  NAND_GATE U7473 ( .I1(n7079), .I2(n6517), .O(n6518) );
  NAND_GATE U7474 ( .I1(n6519), .I2(n6518), .O(n6916) );
  NAND_GATE U7475 ( .I1(n7205), .I2(n6899), .O(n6522) );
  NAND_GATE U7476 ( .I1(n6903), .I2(n6522), .O(n6523) );
  NAND_GATE U7477 ( .I1(n6524), .I2(n6523), .O(n6890) );
  NAND_GATE U7478 ( .I1(n6889), .I2(n6890), .O(n6887) );
  INV_GATE U7479 ( .I1(n6526), .O(n6528) );
  NAND3_GATE U7480 ( .I1(n6525), .I2(n6530), .I3(n6531), .O(n6535) );
  NAND_GATE U7481 ( .I1(n6527), .I2(n6526), .O(n6531) );
  NAND_GATE U7482 ( .I1(n6529), .I2(n6528), .O(n6530) );
  NAND_GATE U7483 ( .I1(n6531), .I2(n6530), .O(n6532) );
  NAND_GATE U7484 ( .I1(n6533), .I2(n6532), .O(n6534) );
  NAND_GATE U7485 ( .I1(n6889), .I2(n783), .O(n6537) );
  NAND_GATE U7486 ( .I1(n6890), .I2(n783), .O(n6536) );
  NAND3_GATE U7487 ( .I1(n6887), .I2(n6537), .I3(n6536), .O(n6878) );
  NAND3_GATE U7488 ( .I1(n6869), .I2(n6878), .I3(n6879), .O(n6539) );
  NAND_GATE U7489 ( .I1(n6538), .I2(n6878), .O(n6871) );
  NAND3_GATE U7490 ( .I1(n6868), .I2(n6539), .I3(n6871), .O(n7116) );
  NAND_GATE U7491 ( .I1(n6547), .I2(n7116), .O(n7118) );
  NAND_GATE U7492 ( .I1(n6541), .I2(n6544), .O(n7105) );
  NAND_GATE U7493 ( .I1(n310), .I2(n6542), .O(n6545) );
  NAND_GATE U7494 ( .I1(n6543), .I2(n747), .O(n6544) );
  NAND_GATE U7495 ( .I1(n6545), .I2(n6544), .O(n7107) );
  NAND_GATE U7496 ( .I1(n7105), .I2(n7112), .O(n6546) );
  NAND_GATE U7497 ( .I1(n7106), .I2(n6546), .O(n7119) );
  NAND_GATE U7498 ( .I1(n7116), .I2(n7119), .O(n6548) );
  NAND_GATE U7499 ( .I1(n6549), .I2(n6864), .O(n6862) );
  NAND_GATE U7500 ( .I1(n6861), .I2(n6864), .O(n6550) );
  NAND3_GATE U7501 ( .I1(n6863), .I2(n6862), .I3(n6550), .O(n6854) );
  NAND_GATE U7502 ( .I1(n6849), .I2(n6854), .O(n6552) );
  NAND_GATE U7503 ( .I1(n6551), .I2(n6854), .O(n6848) );
  NAND3_GATE U7504 ( .I1(n6853), .I2(n6552), .I3(n6848), .O(n6842) );
  NAND_GATE U7505 ( .I1(n6564), .I2(n6842), .O(n6838) );
  INV_GATE U7506 ( .I1(n6553), .O(n6554) );
  NAND_GATE U7507 ( .I1(n6554), .I2(n6557), .O(n6563) );
  NAND_GATE U7508 ( .I1(n6556), .I2(n6555), .O(n6561) );
  NAND_GATE U7509 ( .I1(n6561), .I2(n6560), .O(n6562) );
  NAND_GATE U7510 ( .I1(n6563), .I2(n6562), .O(n6841) );
  NAND_GATE U7511 ( .I1(n6564), .I2(n6841), .O(n6837) );
  NAND_GATE U7512 ( .I1(n6842), .I2(n6841), .O(n6565) );
  NAND3_GATE U7513 ( .I1(n6838), .I2(n6837), .I3(n6565), .O(n6831) );
  NAND_GATE U7514 ( .I1(n6578), .I2(n6831), .O(n6827) );
  OR_GATE U7515 ( .I1(n6569), .I2(n6566), .O(n6577) );
  NAND_GATE U7516 ( .I1(n6567), .I2(n6570), .O(n6575) );
  NAND_GATE U7517 ( .I1(n327), .I2(n6568), .O(n6571) );
  NAND_GATE U7518 ( .I1(n827), .I2(n6569), .O(n6570) );
  NAND_GATE U7519 ( .I1(n6571), .I2(n6570), .O(n6572) );
  NAND_GATE U7520 ( .I1(n6573), .I2(n6572), .O(n6574) );
  NAND_GATE U7521 ( .I1(n6575), .I2(n6574), .O(n6576) );
  NAND_GATE U7522 ( .I1(n6577), .I2(n6576), .O(n6830) );
  NAND_GATE U7523 ( .I1(n6578), .I2(n6830), .O(n6826) );
  NAND_GATE U7524 ( .I1(n6831), .I2(n6830), .O(n6579) );
  NAND3_GATE U7525 ( .I1(n6827), .I2(n6826), .I3(n6579), .O(n6820) );
  NAND_GATE U7526 ( .I1(n6592), .I2(n6820), .O(n6816) );
  INV_GATE U7527 ( .I1(n6580), .O(n6581) );
  NAND_GATE U7528 ( .I1(n6581), .I2(n6585), .O(n6591) );
  INV_GATE U7529 ( .I1(n6585), .O(n6582) );
  NAND_GATE U7530 ( .I1(n6583), .I2(n6582), .O(n6587) );
  NAND_GATE U7531 ( .I1(n6584), .I2(n6587), .O(n6590) );
  NAND_GATE U7532 ( .I1(n834), .I2(n6585), .O(n6586) );
  NAND_GATE U7533 ( .I1(n6587), .I2(n6586), .O(n6588) );
  NAND_GATE U7534 ( .I1(n6820), .I2(n6819), .O(n6593) );
  NAND3_GATE U7535 ( .I1(n6816), .I2(n6815), .I3(n6593), .O(n6809) );
  NAND_GATE U7536 ( .I1(n6607), .I2(n6809), .O(n6805) );
  INV_GATE U7537 ( .I1(n6594), .O(n6595) );
  NAND_GATE U7538 ( .I1(n6595), .I2(n6598), .O(n6606) );
  NAND_GATE U7539 ( .I1(n6597), .I2(n6600), .O(n6604) );
  NAND_GATE U7540 ( .I1(n939), .I2(n6598), .O(n6599) );
  NAND_GATE U7541 ( .I1(n6600), .I2(n6599), .O(n6601) );
  NAND_GATE U7542 ( .I1(n6602), .I2(n6601), .O(n6603) );
  NAND_GATE U7543 ( .I1(n6604), .I2(n6603), .O(n6605) );
  NAND_GATE U7544 ( .I1(n6606), .I2(n6605), .O(n6808) );
  NAND_GATE U7545 ( .I1(n6607), .I2(n6808), .O(n6804) );
  NAND_GATE U7546 ( .I1(n6809), .I2(n6808), .O(n6608) );
  NAND3_GATE U7547 ( .I1(n6805), .I2(n6804), .I3(n6608), .O(n6799) );
  NAND_GATE U7548 ( .I1(n6622), .I2(n6799), .O(n6795) );
  INV_GATE U7549 ( .I1(n6609), .O(n6610) );
  NAND_GATE U7550 ( .I1(n6610), .I2(n6613), .O(n6621) );
  NAND_GATE U7551 ( .I1(n6612), .I2(n6615), .O(n6619) );
  NAND_GATE U7552 ( .I1(n797), .I2(n6613), .O(n6614) );
  NAND_GATE U7553 ( .I1(n6615), .I2(n6614), .O(n6616) );
  NAND_GATE U7554 ( .I1(n6617), .I2(n6616), .O(n6618) );
  NAND_GATE U7555 ( .I1(n6619), .I2(n6618), .O(n6620) );
  NAND_GATE U7556 ( .I1(n6621), .I2(n6620), .O(n6798) );
  NAND_GATE U7557 ( .I1(n6622), .I2(n6798), .O(n6794) );
  NAND_GATE U7558 ( .I1(n6799), .I2(n6798), .O(n6623) );
  NAND3_GATE U7559 ( .I1(n6795), .I2(n6794), .I3(n6623), .O(n6788) );
  NAND_GATE U7560 ( .I1(n6636), .I2(n6788), .O(n6784) );
  INV_GATE U7561 ( .I1(n6624), .O(n6625) );
  NAND_GATE U7562 ( .I1(n6625), .I2(n6628), .O(n6635) );
  NAND_GATE U7563 ( .I1(n6627), .I2(n6630), .O(n6634) );
  NAND_GATE U7564 ( .I1(n750), .I2(n6628), .O(n6629) );
  NAND_GATE U7565 ( .I1(n6630), .I2(n6629), .O(n6631) );
  NAND_GATE U7566 ( .I1(n6632), .I2(n6631), .O(n6633) );
  NAND_GATE U7567 ( .I1(n6788), .I2(n6787), .O(n6637) );
  NAND3_GATE U7568 ( .I1(n6784), .I2(n6783), .I3(n6637), .O(n6777) );
  NAND_GATE U7569 ( .I1(n6651), .I2(n6777), .O(n6773) );
  INV_GATE U7570 ( .I1(n6638), .O(n6639) );
  NAND_GATE U7571 ( .I1(n6639), .I2(n6642), .O(n6650) );
  NAND_GATE U7572 ( .I1(n6641), .I2(n6644), .O(n6648) );
  NAND_GATE U7573 ( .I1(n713), .I2(n6642), .O(n6643) );
  NAND_GATE U7574 ( .I1(n6644), .I2(n6643), .O(n6645) );
  NAND_GATE U7575 ( .I1(n6646), .I2(n6645), .O(n6647) );
  NAND_GATE U7576 ( .I1(n6648), .I2(n6647), .O(n6649) );
  NAND_GATE U7577 ( .I1(n6650), .I2(n6649), .O(n6776) );
  NAND_GATE U7578 ( .I1(n6651), .I2(n6776), .O(n6772) );
  NAND_GATE U7579 ( .I1(n6777), .I2(n6776), .O(n6652) );
  NAND3_GATE U7580 ( .I1(n6773), .I2(n6772), .I3(n6652), .O(n6766) );
  NAND_GATE U7581 ( .I1(n6667), .I2(n6766), .O(n6762) );
  INV_GATE U7582 ( .I1(n6653), .O(n6654) );
  NAND_GATE U7583 ( .I1(n6654), .I2(n6657), .O(n6666) );
  NAND_GATE U7584 ( .I1(n6656), .I2(n6660), .O(n6664) );
  NAND_GATE U7585 ( .I1(n6658), .I2(n6657), .O(n6659) );
  NAND_GATE U7586 ( .I1(n6660), .I2(n6659), .O(n6661) );
  NAND_GATE U7587 ( .I1(n6662), .I2(n6661), .O(n6663) );
  NAND_GATE U7588 ( .I1(n6664), .I2(n6663), .O(n6665) );
  NAND_GATE U7589 ( .I1(n6666), .I2(n6665), .O(n6765) );
  NAND_GATE U7590 ( .I1(n6766), .I2(n6765), .O(n6668) );
  NAND3_GATE U7591 ( .I1(n6762), .I2(n6761), .I3(n6668), .O(n6755) );
  NAND_GATE U7592 ( .I1(n6683), .I2(n6755), .O(n6749) );
  INV_GATE U7593 ( .I1(n6669), .O(n6670) );
  NAND_GATE U7594 ( .I1(n6670), .I2(n6673), .O(n6682) );
  NAND_GATE U7595 ( .I1(n6672), .I2(n6676), .O(n6680) );
  NAND_GATE U7596 ( .I1(n6674), .I2(n6673), .O(n6675) );
  NAND_GATE U7597 ( .I1(n6676), .I2(n6675), .O(n6677) );
  NAND_GATE U7598 ( .I1(n6678), .I2(n6677), .O(n6679) );
  NAND_GATE U7599 ( .I1(n6680), .I2(n6679), .O(n6681) );
  NAND_GATE U7600 ( .I1(n6682), .I2(n6681), .O(n6753) );
  NAND_GATE U7601 ( .I1(n6683), .I2(n6753), .O(n6748) );
  NAND_GATE U7602 ( .I1(n6755), .I2(n6753), .O(n6684) );
  NAND3_GATE U7603 ( .I1(n6749), .I2(n6748), .I3(n6684), .O(n6735) );
  NAND_GATE U7604 ( .I1(n6740), .I2(n6735), .O(n6702) );
  NAND_GATE U7605 ( .I1(B[18]), .I2(A[29]), .O(n6737) );
  INV_GATE U7606 ( .I1(n6737), .O(n6685) );
  NAND_GATE U7607 ( .I1(n6740), .I2(n6685), .O(n6744) );
  NAND_GATE U7608 ( .I1(n6735), .I2(n6685), .O(n6741) );
  NAND_GATE U7609 ( .I1(n6744), .I2(n6741), .O(n6703) );
  INV_GATE U7610 ( .I1(n6690), .O(n6687) );
  NAND_GATE U7611 ( .I1(n6688), .I2(n6687), .O(n6693) );
  NAND_GATE U7612 ( .I1(n6689), .I2(n6693), .O(n6698) );
  NAND_GATE U7613 ( .I1(n6691), .I2(n6690), .O(n6692) );
  NAND_GATE U7614 ( .I1(n6693), .I2(n6692), .O(n6696) );
  NAND_GATE U7615 ( .I1(n6697), .I2(n6696), .O(n6694) );
  NAND_GATE U7616 ( .I1(n6698), .I2(n6694), .O(n6695) );
  NAND_GATE U7617 ( .I1(n6699), .I2(n6695), .O(n6722) );
  NAND_GATE U7618 ( .I1(n6727), .I2(n6722), .O(n6718) );
  INV_GATE U7619 ( .I1(n6698), .O(n6700) );
  NAND_GATE U7620 ( .I1(n6700), .I2(n6699), .O(n6701) );
  NAND_GATE U7621 ( .I1(B[18]), .I2(A[30]), .O(n6725) );
  INV_GATE U7622 ( .I1(n6725), .O(n6728) );
  NAND3_GATE U7623 ( .I1(n6694), .I2(n6701), .I3(n6728), .O(n6729) );
  OR_GATE U7624 ( .I1(n6702), .I2(n6725), .O(n6705) );
  NAND_GATE U7625 ( .I1(n6728), .I2(n6703), .O(n6704) );
  AND3_GATE U7626 ( .I1(n6729), .I2(n6705), .I3(n6704), .O(n6717) );
  NAND3_GATE U7627 ( .I1(n6719), .I2(n6718), .I3(n6717), .O(n6706) );
  NAND_GATE U7628 ( .I1(n6707), .I2(n6706), .O(n6721) );
  NAND_GATE U7629 ( .I1(n14803), .I2(n6721), .O(n6710) );
  NAND_GATE U7630 ( .I1(n6708), .I2(n14802), .O(n6709) );
  NAND_GATE U7631 ( .I1(n6710), .I2(n6709), .O(\A1[48] ) );
  NAND_GATE U7632 ( .I1(n6715), .I2(n6296), .O(n6716) );
  NAND4_GATE U7633 ( .I1(n6719), .I2(n6718), .I3(n6717), .I4(n6716), .O(n6720)
         );
  INV_GATE U7634 ( .I1(n6722), .O(n6726) );
  NAND_GATE U7635 ( .I1(n6727), .I2(n6726), .O(n6724) );
  INV_GATE U7636 ( .I1(n6727), .O(n6730) );
  NAND_GATE U7637 ( .I1(n6730), .I2(n6722), .O(n6723) );
  NAND3_GATE U7638 ( .I1(n6725), .I2(n6724), .I3(n6723), .O(n6734) );
  NAND3_GATE U7639 ( .I1(n6728), .I2(n6727), .I3(n6726), .O(n6733) );
  INV_GATE U7640 ( .I1(n6729), .O(n6731) );
  NAND_GATE U7641 ( .I1(n6731), .I2(n6730), .O(n6732) );
  NAND_GATE U7642 ( .I1(n6740), .I2(n369), .O(n6739) );
  INV_GATE U7643 ( .I1(n6740), .O(n6736) );
  NAND_GATE U7644 ( .I1(n6736), .I2(n6735), .O(n6738) );
  NAND3_GATE U7645 ( .I1(n6739), .I2(n6738), .I3(n6737), .O(n6743) );
  OR_GATE U7646 ( .I1(n6741), .I2(n6740), .O(n6742) );
  NAND_GATE U7647 ( .I1(n6743), .I2(n6742), .O(n6745) );
  INV_GATE U7648 ( .I1(n7158), .O(n7161) );
  NAND_GATE U7649 ( .I1(B[17]), .I2(A[30]), .O(n7165) );
  INV_GATE U7650 ( .I1(n7165), .O(n7159) );
  NAND_GATE U7651 ( .I1(n1429), .I2(A[31]), .O(n7150) );
  NAND_GATE U7652 ( .I1(n6745), .I2(n7165), .O(n7148) );
  INV_GATE U7653 ( .I1(n6746), .O(n6747) );
  NAND_GATE U7654 ( .I1(n6747), .I2(n7165), .O(n7147) );
  OR_GATE U7655 ( .I1(n6748), .I2(n6755), .O(n6751) );
  OR_GATE U7656 ( .I1(n6753), .I2(n6749), .O(n6750) );
  AND_GATE U7657 ( .I1(n6751), .I2(n6750), .O(n6760) );
  INV_GATE U7658 ( .I1(n6755), .O(n6752) );
  NAND_GATE U7659 ( .I1(n6752), .I2(n6753), .O(n6758) );
  INV_GATE U7660 ( .I1(n6753), .O(n6754) );
  NAND_GATE U7661 ( .I1(n6755), .I2(n6754), .O(n6757) );
  NAND3_GATE U7662 ( .I1(n6758), .I2(n6757), .I3(n6756), .O(n6759) );
  NAND_GATE U7663 ( .I1(n6760), .I2(n6759), .O(n7172) );
  INV_GATE U7664 ( .I1(n7172), .O(n7175) );
  NAND_GATE U7665 ( .I1(B[17]), .I2(A[29]), .O(n7179) );
  INV_GATE U7666 ( .I1(n7179), .O(n7173) );
  NAND_GATE U7667 ( .I1(n7175), .I2(n7173), .O(n7170) );
  OR_GATE U7668 ( .I1(n6761), .I2(n6766), .O(n6764) );
  OR_GATE U7669 ( .I1(n6765), .I2(n6762), .O(n6763) );
  AND_GATE U7670 ( .I1(n6764), .I2(n6763), .O(n6771) );
  NAND_GATE U7671 ( .I1(n986), .I2(n6765), .O(n6769) );
  NAND3_GATE U7672 ( .I1(n6769), .I2(n6768), .I3(n6767), .O(n6770) );
  NAND_GATE U7673 ( .I1(n6771), .I2(n6770), .O(n7569) );
  INV_GATE U7674 ( .I1(n7569), .O(n7572) );
  NAND_GATE U7675 ( .I1(B[17]), .I2(A[28]), .O(n7576) );
  INV_GATE U7676 ( .I1(n7576), .O(n7570) );
  NAND_GATE U7677 ( .I1(n7572), .I2(n7570), .O(n7566) );
  OR_GATE U7678 ( .I1(n6772), .I2(n6777), .O(n6775) );
  OR_GATE U7679 ( .I1(n6776), .I2(n6773), .O(n6774) );
  AND_GATE U7680 ( .I1(n6775), .I2(n6774), .O(n6782) );
  NAND_GATE U7681 ( .I1(n987), .I2(n6776), .O(n6780) );
  NAND3_GATE U7682 ( .I1(n6780), .I2(n6779), .I3(n6778), .O(n6781) );
  NAND_GATE U7683 ( .I1(n6782), .I2(n6781), .O(n7552) );
  INV_GATE U7684 ( .I1(n7552), .O(n7555) );
  NAND_GATE U7685 ( .I1(B[17]), .I2(A[27]), .O(n7559) );
  INV_GATE U7686 ( .I1(n7559), .O(n7553) );
  NAND_GATE U7687 ( .I1(n7555), .I2(n7553), .O(n7549) );
  OR_GATE U7688 ( .I1(n6783), .I2(n6788), .O(n6786) );
  OR_GATE U7689 ( .I1(n6787), .I2(n6784), .O(n6785) );
  AND_GATE U7690 ( .I1(n6786), .I2(n6785), .O(n6793) );
  NAND_GATE U7691 ( .I1(n982), .I2(n6787), .O(n6791) );
  NAND3_GATE U7692 ( .I1(n6791), .I2(n6790), .I3(n6789), .O(n6792) );
  NAND_GATE U7693 ( .I1(n6793), .I2(n6792), .O(n7536) );
  NAND_GATE U7694 ( .I1(B[17]), .I2(A[26]), .O(n7542) );
  INV_GATE U7695 ( .I1(n7542), .O(n7537) );
  NAND_GATE U7696 ( .I1(n318), .I2(n7537), .O(n7534) );
  OR_GATE U7697 ( .I1(n6794), .I2(n6799), .O(n6797) );
  OR_GATE U7698 ( .I1(n6798), .I2(n6795), .O(n6796) );
  NAND_GATE U7699 ( .I1(n973), .I2(n6798), .O(n6802) );
  NAND3_GATE U7700 ( .I1(n6802), .I2(n6801), .I3(n6800), .O(n6803) );
  NAND_GATE U7701 ( .I1(B[17]), .I2(A[25]), .O(n7527) );
  INV_GATE U7702 ( .I1(n7527), .O(n7522) );
  NAND_GATE U7703 ( .I1(n938), .I2(n7522), .O(n7519) );
  OR_GATE U7704 ( .I1(n6804), .I2(n6809), .O(n6807) );
  OR_GATE U7705 ( .I1(n6808), .I2(n6805), .O(n6806) );
  AND_GATE U7706 ( .I1(n6807), .I2(n6806), .O(n6814) );
  NAND_GATE U7707 ( .I1(n960), .I2(n6808), .O(n6812) );
  NAND3_GATE U7708 ( .I1(n6812), .I2(n6811), .I3(n6810), .O(n6813) );
  NAND_GATE U7709 ( .I1(B[17]), .I2(A[24]), .O(n7512) );
  INV_GATE U7710 ( .I1(n7512), .O(n7507) );
  NAND_GATE U7711 ( .I1(n910), .I2(n7507), .O(n7504) );
  OR_GATE U7712 ( .I1(n6815), .I2(n6820), .O(n6818) );
  OR_GATE U7713 ( .I1(n6819), .I2(n6816), .O(n6817) );
  AND_GATE U7714 ( .I1(n6818), .I2(n6817), .O(n6825) );
  NAND_GATE U7715 ( .I1(n962), .I2(n6819), .O(n6823) );
  NAND3_GATE U7716 ( .I1(n6823), .I2(n6822), .I3(n6821), .O(n6824) );
  NAND_GATE U7717 ( .I1(n6825), .I2(n6824), .O(n7491) );
  NAND_GATE U7718 ( .I1(B[17]), .I2(A[23]), .O(n7497) );
  INV_GATE U7719 ( .I1(n7497), .O(n7492) );
  NAND_GATE U7720 ( .I1(n833), .I2(n7492), .O(n7489) );
  OR_GATE U7721 ( .I1(n6830), .I2(n6827), .O(n6828) );
  AND_GATE U7722 ( .I1(n6829), .I2(n6828), .O(n6836) );
  NAND_GATE U7723 ( .I1(n949), .I2(n6830), .O(n6834) );
  NAND3_GATE U7724 ( .I1(n6834), .I2(n6833), .I3(n6832), .O(n6835) );
  NAND_GATE U7725 ( .I1(n6836), .I2(n6835), .O(n7481) );
  INV_GATE U7726 ( .I1(n7481), .O(n7480) );
  NAND_GATE U7727 ( .I1(B[17]), .I2(A[22]), .O(n7482) );
  INV_GATE U7728 ( .I1(n7482), .O(n7478) );
  NAND_GATE U7729 ( .I1(n7480), .I2(n7478), .O(n7475) );
  OR_GATE U7730 ( .I1(n6841), .I2(n6838), .O(n6839) );
  AND_GATE U7731 ( .I1(n6840), .I2(n6839), .O(n6847) );
  NAND_GATE U7732 ( .I1(n953), .I2(n6841), .O(n6845) );
  NAND3_GATE U7733 ( .I1(n6845), .I2(n6844), .I3(n6843), .O(n6846) );
  NAND_GATE U7734 ( .I1(B[17]), .I2(A[21]), .O(n7468) );
  INV_GATE U7735 ( .I1(n7468), .O(n7466) );
  NAND_GATE U7736 ( .I1(n825), .I2(n7466), .O(n7463) );
  OR_GATE U7737 ( .I1(n6848), .I2(n6849), .O(n6857) );
  NAND_GATE U7738 ( .I1(n6849), .I2(n505), .O(n6851) );
  NAND3_GATE U7739 ( .I1(n6852), .I2(n6851), .I3(n6850), .O(n6856) );
  OR_GATE U7740 ( .I1(n6854), .I2(n6853), .O(n6855) );
  NAND3_GATE U7741 ( .I1(n6857), .I2(n6856), .I3(n6855), .O(n7187) );
  NAND_GATE U7742 ( .I1(B[17]), .I2(A[20]), .O(n7188) );
  INV_GATE U7743 ( .I1(n7188), .O(n7185) );
  NAND_GATE U7744 ( .I1(n703), .I2(n7185), .O(n7191) );
  NAND_GATE U7745 ( .I1(B[17]), .I2(A[19]), .O(n7712) );
  INV_GATE U7746 ( .I1(n7712), .O(n7197) );
  NAND_GATE U7747 ( .I1(n6861), .I2(n665), .O(n6859) );
  NAND3_GATE U7748 ( .I1(n6860), .I2(n6859), .I3(n6858), .O(n6867) );
  OR_GATE U7749 ( .I1(n6862), .I2(n6861), .O(n6866) );
  OR_GATE U7750 ( .I1(n6864), .I2(n6863), .O(n6865) );
  NAND3_GATE U7751 ( .I1(n6867), .I2(n6866), .I3(n6865), .O(n7198) );
  INV_GATE U7752 ( .I1(n7198), .O(n7200) );
  NAND_GATE U7753 ( .I1(n7197), .I2(n7200), .O(n7196) );
  NAND_GATE U7754 ( .I1(B[17]), .I2(A[18]), .O(n7445) );
  INV_GATE U7755 ( .I1(n7445), .O(n7448) );
  NAND_GATE U7756 ( .I1(B[17]), .I2(A[17]), .O(n7440) );
  INV_GATE U7757 ( .I1(n7440), .O(n7433) );
  OR_GATE U7758 ( .I1(n6878), .I2(n6868), .O(n6886) );
  NAND_GATE U7759 ( .I1(n6876), .I2(n6875), .O(n6869) );
  NAND_GATE U7760 ( .I1(n6870), .I2(n6869), .O(n6874) );
  INV_GATE U7761 ( .I1(n6871), .O(n6873) );
  NAND3_GATE U7762 ( .I1(n6874), .I2(n6873), .I3(n6872), .O(n6885) );
  NAND_GATE U7763 ( .I1(n6879), .I2(n6869), .O(n6877) );
  NAND_GATE U7764 ( .I1(n6878), .I2(n6877), .O(n6883) );
  INV_GATE U7765 ( .I1(n6878), .O(n6880) );
  NAND3_GATE U7766 ( .I1(n6880), .I2(n6869), .I3(n6879), .O(n6882) );
  NAND3_GATE U7767 ( .I1(n6883), .I2(n6882), .I3(n6881), .O(n6884) );
  NAND3_GATE U7768 ( .I1(n6886), .I2(n6885), .I3(n6884), .O(n7435) );
  INV_GATE U7769 ( .I1(n7435), .O(n7437) );
  INV_GATE U7770 ( .I1(n6887), .O(n6888) );
  NAND_GATE U7771 ( .I1(n6888), .I2(n360), .O(n6897) );
  INV_GATE U7772 ( .I1(n6890), .O(n6891) );
  NAND3_GATE U7773 ( .I1(n783), .I2(n6891), .I3(n6889), .O(n6896) );
  NAND_GATE U7774 ( .I1(n6890), .I2(n360), .O(n6894) );
  NAND_GATE U7775 ( .I1(n6891), .I2(n783), .O(n6893) );
  NAND3_GATE U7776 ( .I1(n6894), .I2(n6893), .I3(n6892), .O(n6895) );
  NAND3_GATE U7777 ( .I1(n6897), .I2(n6896), .I3(n6895), .O(n7418) );
  NAND_GATE U7778 ( .I1(B[17]), .I2(A[16]), .O(n7419) );
  INV_GATE U7779 ( .I1(n7419), .O(n7417) );
  NAND_GATE U7780 ( .I1(n353), .I2(n7417), .O(n7423) );
  INV_GATE U7781 ( .I1(n6903), .O(n6898) );
  NAND_GATE U7782 ( .I1(n6904), .I2(n6900), .O(n7206) );
  NAND_GATE U7783 ( .I1(n6902), .I2(n6903), .O(n6901) );
  NAND_GATE U7784 ( .I1(n6899), .I2(n6898), .O(n6900) );
  NAND_GATE U7785 ( .I1(n6901), .I2(n6900), .O(n7204) );
  NAND_GATE U7786 ( .I1(n7206), .I2(n7209), .O(n6905) );
  NAND3_GATE U7787 ( .I1(n6904), .I2(n6903), .I3(n6902), .O(n7207) );
  NAND_GATE U7788 ( .I1(n6905), .I2(n7207), .O(n7215) );
  NAND_GATE U7789 ( .I1(B[17]), .I2(A[14]), .O(n7224) );
  INV_GATE U7790 ( .I1(n7224), .O(n7223) );
  NAND_GATE U7791 ( .I1(n6906), .I2(n6520), .O(n6908) );
  NAND3_GATE U7792 ( .I1(n6908), .I2(n1396), .I3(n6907), .O(n6911) );
  OR_GATE U7793 ( .I1(n6916), .I2(n6909), .O(n6910) );
  AND_GATE U7794 ( .I1(n6911), .I2(n6910), .O(n7095) );
  NAND_GATE U7795 ( .I1(n6914), .I2(n6520), .O(n6915) );
  OR_GATE U7796 ( .I1(n6915), .I2(n6916), .O(n6919) );
  NAND_GATE U7797 ( .I1(n6916), .I2(n6915), .O(n6918) );
  NAND3_GATE U7798 ( .I1(n6919), .I2(n6918), .I3(n6917), .O(n7096) );
  NAND_GATE U7799 ( .I1(n7095), .I2(n7096), .O(n7225) );
  INV_GATE U7800 ( .I1(n7225), .O(n7221) );
  NAND_GATE U7801 ( .I1(n7223), .I2(n7221), .O(n7229) );
  NAND_GATE U7802 ( .I1(B[17]), .I2(A[13]), .O(n7233) );
  INV_GATE U7803 ( .I1(n7233), .O(n7086) );
  OR_GATE U7804 ( .I1(n6920), .I2(n6932), .O(n6924) );
  OR_GATE U7805 ( .I1(n6922), .I2(n6921), .O(n6923) );
  AND_GATE U7806 ( .I1(n6924), .I2(n6923), .O(n6937) );
  INV_GATE U7807 ( .I1(n6932), .O(n6928) );
  NAND3_GATE U7808 ( .I1(n6929), .I2(n6928), .I3(n6930), .O(n6935) );
  NAND_GATE U7809 ( .I1(n6930), .I2(n6929), .O(n6931) );
  NAND_GATE U7810 ( .I1(n6932), .I2(n6931), .O(n6934) );
  NAND3_GATE U7811 ( .I1(n6935), .I2(n6934), .I3(n6933), .O(n6936) );
  NAND_GATE U7812 ( .I1(n6937), .I2(n6936), .O(n7397) );
  NAND_GATE U7813 ( .I1(B[17]), .I2(A[12]), .O(n7398) );
  INV_GATE U7814 ( .I1(n7398), .O(n7405) );
  NAND_GATE U7815 ( .I1(n757), .I2(n7405), .O(n7395) );
  NAND_GATE U7816 ( .I1(B[17]), .I2(A[11]), .O(n7249) );
  INV_GATE U7817 ( .I1(n7249), .O(n7074) );
  NAND_GATE U7818 ( .I1(B[17]), .I2(A[10]), .O(n7381) );
  INV_GATE U7819 ( .I1(n6951), .O(n6952) );
  NAND3_GATE U7820 ( .I1(n6940), .I2(n6952), .I3(n6939), .O(n7056) );
  NAND_GATE U7821 ( .I1(n6946), .I2(n6945), .O(n6947) );
  NAND_GATE U7822 ( .I1(n6498), .I2(n6947), .O(n6948) );
  NAND_GATE U7823 ( .I1(n6949), .I2(n6948), .O(n6953) );
  NAND_GATE U7824 ( .I1(n6954), .I2(n6953), .O(n6950) );
  NAND_GATE U7825 ( .I1(n6951), .I2(n6950), .O(n7060) );
  NAND3_GATE U7826 ( .I1(n6954), .I2(n6953), .I3(n6952), .O(n7059) );
  NAND3_GATE U7827 ( .I1(n7061), .I2(n7060), .I3(n7059), .O(n6955) );
  NAND3_GATE U7828 ( .I1(n7057), .I2(n7056), .I3(n6955), .O(n7382) );
  NAND_GATE U7829 ( .I1(B[17]), .I2(A[9]), .O(n7265) );
  INV_GATE U7830 ( .I1(n7265), .O(n7268) );
  NAND_GATE U7831 ( .I1(B[17]), .I2(A[8]), .O(n7900) );
  INV_GATE U7832 ( .I1(n7900), .O(n7368) );
  NAND_GATE U7833 ( .I1(n1272), .I2(n6962), .O(n6958) );
  NAND_GATE U7834 ( .I1(n6956), .I2(n694), .O(n6957) );
  NAND3_GATE U7835 ( .I1(n6959), .I2(n6958), .I3(n6957), .O(n6965) );
  NAND3_GATE U7836 ( .I1(n1272), .I2(n6960), .I3(n6962), .O(n6964) );
  OR_GATE U7837 ( .I1(n6962), .I2(n6961), .O(n6963) );
  NAND3_GATE U7838 ( .I1(n6965), .I2(n6964), .I3(n6963), .O(n7370) );
  INV_GATE U7839 ( .I1(n7370), .O(n7372) );
  NAND_GATE U7840 ( .I1(n7368), .I2(n7372), .O(n7367) );
  NAND_GATE U7841 ( .I1(B[17]), .I2(A[6]), .O(n7354) );
  INV_GATE U7842 ( .I1(n7354), .O(n7349) );
  NAND_GATE U7843 ( .I1(n1364), .I2(n6972), .O(n6967) );
  NAND3_GATE U7844 ( .I1(n6968), .I2(n6967), .I3(n6966), .O(n6975) );
  OR_GATE U7845 ( .I1(n6970), .I2(n6969), .O(n6974) );
  OR_GATE U7846 ( .I1(n6972), .I2(n6971), .O(n6973) );
  NAND3_GATE U7847 ( .I1(n6975), .I2(n6974), .I3(n6973), .O(n7352) );
  INV_GATE U7848 ( .I1(n7352), .O(n7350) );
  NAND_GATE U7849 ( .I1(n7349), .I2(n7350), .O(n7357) );
  NAND_GATE U7850 ( .I1(B[17]), .I2(A[5]), .O(n7284) );
  INV_GATE U7851 ( .I1(n7284), .O(n7026) );
  OR_GATE U7852 ( .I1(n6981), .I2(n6977), .O(n6978) );
  AND_GATE U7853 ( .I1(n6979), .I2(n6978), .O(n6987) );
  INV_GATE U7854 ( .I1(n6982), .O(n6980) );
  NAND_GATE U7855 ( .I1(n6980), .I2(n6981), .O(n6985) );
  NAND_GATE U7856 ( .I1(n6982), .I2(n1316), .O(n6984) );
  NAND3_GATE U7857 ( .I1(n6985), .I2(n6984), .I3(n6983), .O(n6986) );
  NAND_GATE U7858 ( .I1(n6987), .I2(n6986), .O(n7333) );
  INV_GATE U7859 ( .I1(n7333), .O(n7336) );
  NAND_GATE U7860 ( .I1(B[17]), .I2(A[4]), .O(n7340) );
  INV_GATE U7861 ( .I1(n7340), .O(n7334) );
  NAND_GATE U7862 ( .I1(n7336), .I2(n7334), .O(n7331) );
  NAND_GATE U7863 ( .I1(B[17]), .I2(A[3]), .O(n7300) );
  INV_GATE U7864 ( .I1(n7300), .O(n7008) );
  NAND_GATE U7865 ( .I1(B[17]), .I2(A[2]), .O(n7322) );
  INV_GATE U7866 ( .I1(n7322), .O(n7316) );
  NAND_GATE U7867 ( .I1(n14241), .I2(n6988), .O(n6989) );
  NAND_GATE U7868 ( .I1(B[19]), .I2(n6989), .O(n6993) );
  NAND_GATE U7869 ( .I1(n1431), .I2(A[1]), .O(n6990) );
  NAND_GATE U7870 ( .I1(n724), .I2(n6990), .O(n6991) );
  NAND_GATE U7871 ( .I1(B[18]), .I2(n6991), .O(n6992) );
  NAND_GATE U7872 ( .I1(n6993), .I2(n6992), .O(n7318) );
  NAND_GATE U7873 ( .I1(n7316), .I2(n7318), .O(n7313) );
  NAND3_GATE U7874 ( .I1(B[17]), .I2(B[18]), .I3(n1254), .O(n7314) );
  INV_GATE U7875 ( .I1(n7314), .O(n7317) );
  INV_GATE U7876 ( .I1(n7318), .O(n7315) );
  NAND_GATE U7877 ( .I1(n7322), .I2(n7315), .O(n6994) );
  NAND_GATE U7878 ( .I1(n7317), .I2(n6994), .O(n6995) );
  NAND_GATE U7879 ( .I1(n7313), .I2(n6995), .O(n7299) );
  NAND_GATE U7880 ( .I1(n7008), .I2(n7299), .O(n7295) );
  OR_GATE U7881 ( .I1(n6997), .I2(n6996), .O(n7007) );
  NAND_GATE U7882 ( .I1(n6998), .I2(n6997), .O(n7002) );
  NAND_GATE U7883 ( .I1(n6999), .I2(n7002), .O(n7005) );
  NAND_GATE U7884 ( .I1(n7005), .I2(n7004), .O(n7006) );
  NAND_GATE U7885 ( .I1(n7007), .I2(n7006), .O(n7298) );
  NAND_GATE U7886 ( .I1(n7299), .I2(n7298), .O(n7009) );
  NAND_GATE U7887 ( .I1(n7008), .I2(n7298), .O(n7294) );
  NAND3_GATE U7888 ( .I1(n7295), .I2(n7009), .I3(n7294), .O(n7335) );
  NAND_GATE U7889 ( .I1(n7333), .I2(n7340), .O(n7010) );
  NAND_GATE U7890 ( .I1(n7335), .I2(n7010), .O(n7011) );
  NAND_GATE U7891 ( .I1(n7331), .I2(n7011), .O(n7287) );
  NAND_GATE U7892 ( .I1(n7026), .I2(n7287), .O(n7289) );
  INV_GATE U7893 ( .I1(n7012), .O(n7013) );
  NAND_GATE U7894 ( .I1(n7013), .I2(n7016), .O(n7025) );
  NAND_GATE U7895 ( .I1(n7014), .I2(n792), .O(n7019) );
  NAND_GATE U7896 ( .I1(n7015), .I2(n7019), .O(n7023) );
  NAND_GATE U7897 ( .I1(n7019), .I2(n7018), .O(n7020) );
  NAND_GATE U7898 ( .I1(n7021), .I2(n7020), .O(n7022) );
  NAND_GATE U7899 ( .I1(n7023), .I2(n7022), .O(n7024) );
  NAND_GATE U7900 ( .I1(n7025), .I2(n7024), .O(n7290) );
  NAND_GATE U7901 ( .I1(n7287), .I2(n7290), .O(n7027) );
  NAND_GATE U7902 ( .I1(n7026), .I2(n7290), .O(n7288) );
  NAND3_GATE U7903 ( .I1(n7289), .I2(n7027), .I3(n7288), .O(n7358) );
  NAND_GATE U7904 ( .I1(n7354), .I2(n7352), .O(n7028) );
  NAND_GATE U7905 ( .I1(n7358), .I2(n7028), .O(n7029) );
  NAND_GATE U7906 ( .I1(n7357), .I2(n7029), .O(n7277) );
  NAND3_GATE U7907 ( .I1(n7031), .I2(n1044), .I3(n7030), .O(n7037) );
  NAND_GATE U7908 ( .I1(n7034), .I2(n7039), .O(n7036) );
  NAND3_GATE U7909 ( .I1(n7034), .I2(n7033), .I3(n7032), .O(n7035) );
  NAND4_GATE U7910 ( .I1(n7038), .I2(n7037), .I3(n7036), .I4(n7035), .O(n7041)
         );
  NAND_GATE U7911 ( .I1(n1365), .I2(n7039), .O(n7040) );
  NAND_GATE U7912 ( .I1(n7041), .I2(n7040), .O(n7280) );
  NAND_GATE U7913 ( .I1(n7277), .I2(n7280), .O(n7043) );
  NAND_GATE U7914 ( .I1(B[17]), .I2(A[7]), .O(n7276) );
  INV_GATE U7915 ( .I1(n7276), .O(n7042) );
  NAND_GATE U7916 ( .I1(n7042), .I2(n7280), .O(n7278) );
  NAND_GATE U7917 ( .I1(n7042), .I2(n7277), .O(n7279) );
  NAND3_GATE U7918 ( .I1(n7043), .I2(n7278), .I3(n7279), .O(n7371) );
  NAND_GATE U7919 ( .I1(n7900), .I2(n7370), .O(n7044) );
  NAND_GATE U7920 ( .I1(n7371), .I2(n7044), .O(n7045) );
  NAND_GATE U7921 ( .I1(n7367), .I2(n7045), .O(n7264) );
  NAND_GATE U7922 ( .I1(n7268), .I2(n7264), .O(n7269) );
  NAND3_GATE U7923 ( .I1(n7047), .I2(n7050), .I3(n7051), .O(n7259) );
  INV_GATE U7924 ( .I1(n7050), .O(n7048) );
  NAND_GATE U7925 ( .I1(n7049), .I2(n7048), .O(n7046) );
  NAND_GATE U7926 ( .I1(n7051), .I2(n7050), .O(n7052) );
  NAND_GATE U7927 ( .I1(n7046), .I2(n7052), .O(n7260) );
  NAND_GATE U7928 ( .I1(n7259), .I2(n7053), .O(n7270) );
  NAND_GATE U7929 ( .I1(n7264), .I2(n7270), .O(n7055) );
  NAND_GATE U7930 ( .I1(n7268), .I2(n7270), .O(n7054) );
  NAND3_GATE U7931 ( .I1(n7269), .I2(n7055), .I3(n7054), .O(n7387) );
  NAND_GATE U7932 ( .I1(n7057), .I2(n7056), .O(n7058) );
  NAND_GATE U7933 ( .I1(n7381), .I2(n7058), .O(n7063) );
  NAND4_GATE U7934 ( .I1(n7061), .I2(n7060), .I3(n7381), .I4(n7059), .O(n7062)
         );
  NAND3_GATE U7935 ( .I1(n7387), .I2(n7063), .I3(n7062), .O(n7064) );
  NAND_GATE U7936 ( .I1(n7386), .I2(n7064), .O(n7252) );
  NAND_GATE U7937 ( .I1(n7074), .I2(n7252), .O(n7254) );
  NAND3_GATE U7938 ( .I1(n7066), .I2(n7069), .I3(n7070), .O(n7243) );
  INV_GATE U7939 ( .I1(n7069), .O(n7067) );
  NAND_GATE U7940 ( .I1(n7068), .I2(n7067), .O(n7065) );
  NAND_GATE U7941 ( .I1(n7070), .I2(n7069), .O(n7071) );
  NAND_GATE U7942 ( .I1(n7065), .I2(n7071), .O(n7244) );
  NAND_GATE U7943 ( .I1(n7073), .I2(n7248), .O(n7072) );
  NAND_GATE U7944 ( .I1(n7243), .I2(n7072), .O(n7255) );
  NAND_GATE U7945 ( .I1(n7252), .I2(n7255), .O(n7076) );
  NAND_GATE U7946 ( .I1(n7243), .I2(n1347), .O(n7075) );
  NAND3_GATE U7947 ( .I1(n7248), .I2(n7075), .I3(n7074), .O(n7253) );
  NAND3_GATE U7948 ( .I1(n7254), .I2(n7076), .I3(n7253), .O(n7399) );
  NAND_GATE U7949 ( .I1(n7397), .I2(n7398), .O(n7077) );
  NAND_GATE U7950 ( .I1(n7399), .I2(n7077), .O(n7078) );
  NAND_GATE U7951 ( .I1(n7395), .I2(n7078), .O(n7236) );
  NAND_GATE U7952 ( .I1(n7086), .I2(n7236), .O(n7238) );
  INV_GATE U7953 ( .I1(n7079), .O(n7082) );
  NAND_GATE U7954 ( .I1(n7083), .I2(n7082), .O(n7087) );
  NAND3_GATE U7955 ( .I1(n7088), .I2(n7079), .I3(n7080), .O(n7093) );
  NAND3_GATE U7956 ( .I1(n7088), .I2(n7087), .I3(n7093), .O(n7085) );
  NAND3_GATE U7957 ( .I1(n7080), .I2(n7079), .I3(n7081), .O(n7089) );
  NAND3_GATE U7958 ( .I1(n7083), .I2(n7082), .I3(n7081), .O(n7091) );
  AND_GATE U7959 ( .I1(n7089), .I2(n7091), .O(n7084) );
  NAND3_GATE U7960 ( .I1(n7086), .I2(n7085), .I3(n7084), .O(n7237) );
  NAND_GATE U7961 ( .I1(n7088), .I2(n7087), .O(n7090) );
  NAND3_GATE U7962 ( .I1(n7091), .I2(n7090), .I3(n7089), .O(n7092) );
  NAND_GATE U7963 ( .I1(n7093), .I2(n7092), .O(n7239) );
  NAND_GATE U7964 ( .I1(n7236), .I2(n7239), .O(n7094) );
  NAND3_GATE U7965 ( .I1(n7238), .I2(n7237), .I3(n7094), .O(n7230) );
  NAND3_GATE U7966 ( .I1(n7096), .I2(n7230), .I3(n7095), .O(n7098) );
  NAND_GATE U7967 ( .I1(n7223), .I2(n7230), .O(n7097) );
  NAND3_GATE U7968 ( .I1(n7229), .I2(n7098), .I3(n7097), .O(n7218) );
  NAND_GATE U7969 ( .I1(n7215), .I2(n7218), .O(n7100) );
  NAND_GATE U7970 ( .I1(B[17]), .I2(A[15]), .O(n7212) );
  INV_GATE U7971 ( .I1(n7212), .O(n7099) );
  NAND_GATE U7972 ( .I1(n7099), .I2(n7218), .O(n7216) );
  NAND_GATE U7973 ( .I1(n7099), .I2(n7215), .O(n7217) );
  NAND_GATE U7974 ( .I1(n7418), .I2(n7419), .O(n7101) );
  NAND_GATE U7975 ( .I1(n7424), .I2(n7101), .O(n7102) );
  NAND_GATE U7976 ( .I1(n7423), .I2(n7102), .O(n7436) );
  NAND_GATE U7977 ( .I1(n7440), .I2(n7435), .O(n7103) );
  NAND_GATE U7978 ( .I1(n7436), .I2(n7103), .O(n7104) );
  NAND_GATE U7979 ( .I1(n7430), .I2(n7104), .O(n7449) );
  NAND_GATE U7980 ( .I1(n7448), .I2(n7449), .O(n7453) );
  NAND_GATE U7981 ( .I1(n7108), .I2(n7107), .O(n7112) );
  NAND_GATE U7982 ( .I1(n7110), .I2(n7112), .O(n7109) );
  NAND_GATE U7983 ( .I1(n7116), .I2(n7109), .O(n7114) );
  INV_GATE U7984 ( .I1(n7116), .O(n7111) );
  NAND3_GATE U7985 ( .I1(n7112), .I2(n7111), .I3(n7110), .O(n7113) );
  NAND3_GATE U7986 ( .I1(n7115), .I2(n7114), .I3(n7113), .O(n7122) );
  OR_GATE U7987 ( .I1(n7117), .I2(n7116), .O(n7121) );
  OR_GATE U7988 ( .I1(n7119), .I2(n7118), .O(n7120) );
  NAND3_GATE U7989 ( .I1(n7122), .I2(n7121), .I3(n7120), .O(n7454) );
  NAND_GATE U7990 ( .I1(n7445), .I2(n7446), .O(n7123) );
  NAND_GATE U7991 ( .I1(n307), .I2(n7123), .O(n7124) );
  NAND_GATE U7992 ( .I1(n7712), .I2(n7198), .O(n7125) );
  NAND_GATE U7993 ( .I1(n7199), .I2(n7125), .O(n7126) );
  NAND_GATE U7994 ( .I1(n7196), .I2(n7126), .O(n7192) );
  NAND_GATE U7995 ( .I1(n7187), .I2(n7188), .O(n7127) );
  NAND_GATE U7996 ( .I1(n7192), .I2(n7127), .O(n7128) );
  NAND_GATE U7997 ( .I1(n7191), .I2(n7128), .O(n7467) );
  NAND_GATE U7998 ( .I1(n808), .I2(n7468), .O(n7129) );
  NAND_GATE U7999 ( .I1(n7467), .I2(n7129), .O(n7130) );
  NAND_GATE U8000 ( .I1(n7463), .I2(n7130), .O(n7479) );
  NAND_GATE U8001 ( .I1(n7481), .I2(n7482), .O(n7131) );
  NAND_GATE U8002 ( .I1(n7479), .I2(n7131), .O(n7132) );
  NAND_GATE U8003 ( .I1(n7475), .I2(n7132), .O(n7493) );
  NAND_GATE U8004 ( .I1(n7491), .I2(n7497), .O(n7133) );
  NAND_GATE U8005 ( .I1(n7493), .I2(n7133), .O(n7134) );
  NAND_GATE U8006 ( .I1(n7489), .I2(n7134), .O(n7508) );
  NAND_GATE U8007 ( .I1(n7506), .I2(n7512), .O(n7135) );
  NAND_GATE U8008 ( .I1(n7508), .I2(n7135), .O(n7136) );
  NAND_GATE U8009 ( .I1(n7504), .I2(n7136), .O(n7523) );
  NAND_GATE U8010 ( .I1(n7521), .I2(n7527), .O(n7137) );
  NAND_GATE U8011 ( .I1(n7523), .I2(n7137), .O(n7138) );
  NAND_GATE U8012 ( .I1(n7519), .I2(n7138), .O(n7538) );
  NAND_GATE U8013 ( .I1(n7536), .I2(n7542), .O(n7139) );
  NAND_GATE U8014 ( .I1(n7538), .I2(n7139), .O(n7140) );
  NAND_GATE U8015 ( .I1(n7534), .I2(n7140), .O(n7554) );
  NAND_GATE U8016 ( .I1(n7552), .I2(n7559), .O(n7141) );
  NAND_GATE U8017 ( .I1(n7554), .I2(n7141), .O(n7142) );
  NAND_GATE U8018 ( .I1(n7549), .I2(n7142), .O(n7571) );
  NAND_GATE U8019 ( .I1(n7569), .I2(n7576), .O(n7143) );
  NAND_GATE U8020 ( .I1(n7571), .I2(n7143), .O(n7144) );
  NAND_GATE U8021 ( .I1(n7566), .I2(n7144), .O(n7174) );
  NAND_GATE U8022 ( .I1(n7172), .I2(n7179), .O(n7145) );
  NAND_GATE U8023 ( .I1(n7174), .I2(n7145), .O(n7146) );
  NAND_GATE U8024 ( .I1(n7170), .I2(n7146), .O(n7160) );
  NAND3_GATE U8025 ( .I1(n7148), .I2(n7147), .I3(n7160), .O(n7149) );
  NAND3_GATE U8026 ( .I1(n7155), .I2(n7150), .I3(n7149), .O(n14806) );
  NAND_GATE U8027 ( .I1(n14805), .I2(n14806), .O(n7154) );
  NAND_GATE U8028 ( .I1(n14804), .I2(n7154), .O(n7152) );
  NAND_GATE U8029 ( .I1(n7152), .I2(n7151), .O(\A1[47] ) );
  NAND_GATE U8030 ( .I1(n7154), .I2(n7153), .O(n7586) );
  INV_GATE U8031 ( .I1(n7586), .O(n14808) );
  INV_GATE U8032 ( .I1(n7155), .O(n7156) );
  NAND_GATE U8033 ( .I1(n7156), .I2(n7160), .O(n7169) );
  INV_GATE U8034 ( .I1(n7160), .O(n7157) );
  NAND_GATE U8035 ( .I1(n7158), .I2(n7157), .O(n7163) );
  NAND_GATE U8036 ( .I1(n7159), .I2(n7163), .O(n7167) );
  NAND_GATE U8037 ( .I1(n7161), .I2(n7160), .O(n7162) );
  NAND_GATE U8038 ( .I1(n7163), .I2(n7162), .O(n7164) );
  NAND_GATE U8039 ( .I1(n7165), .I2(n7164), .O(n7166) );
  NAND_GATE U8040 ( .I1(n7167), .I2(n7166), .O(n7168) );
  NAND_GATE U8041 ( .I1(n7169), .I2(n7168), .O(n7589) );
  NAND_GATE U8042 ( .I1(B[16]), .I2(A[30]), .O(n7602) );
  INV_GATE U8043 ( .I1(n7602), .O(n7583) );
  INV_GATE U8044 ( .I1(n7170), .O(n7171) );
  NAND_GATE U8045 ( .I1(n7171), .I2(n7174), .O(n7183) );
  NAND_GATE U8046 ( .I1(n7173), .I2(n7177), .O(n7181) );
  NAND_GATE U8047 ( .I1(n7175), .I2(n7174), .O(n7176) );
  NAND_GATE U8048 ( .I1(n7177), .I2(n7176), .O(n7178) );
  NAND_GATE U8049 ( .I1(n7179), .I2(n7178), .O(n7180) );
  NAND_GATE U8050 ( .I1(n7181), .I2(n7180), .O(n7182) );
  NAND_GATE U8051 ( .I1(n7183), .I2(n7182), .O(n7600) );
  NAND_GATE U8052 ( .I1(n7583), .I2(n7600), .O(n7595) );
  NAND_GATE U8053 ( .I1(B[16]), .I2(A[29]), .O(n7613) );
  INV_GATE U8054 ( .I1(n7613), .O(n7581) );
  NAND_GATE U8055 ( .I1(B[16]), .I2(A[28]), .O(n7624) );
  INV_GATE U8056 ( .I1(n7624), .O(n7564) );
  NAND_GATE U8057 ( .I1(B[16]), .I2(A[27]), .O(n7635) );
  INV_GATE U8058 ( .I1(n7635), .O(n7547) );
  NAND_GATE U8059 ( .I1(B[16]), .I2(A[26]), .O(n7645) );
  INV_GATE U8060 ( .I1(n7645), .O(n7532) );
  NAND_GATE U8061 ( .I1(B[16]), .I2(A[25]), .O(n7655) );
  INV_GATE U8062 ( .I1(n7655), .O(n7517) );
  NAND_GATE U8063 ( .I1(B[16]), .I2(A[24]), .O(n7665) );
  INV_GATE U8064 ( .I1(n7665), .O(n7502) );
  NAND_GATE U8065 ( .I1(B[16]), .I2(A[23]), .O(n7676) );
  INV_GATE U8066 ( .I1(n7676), .O(n7487) );
  NAND_GATE U8067 ( .I1(B[16]), .I2(A[22]), .O(n7687) );
  INV_GATE U8068 ( .I1(n7687), .O(n7473) );
  NAND_GATE U8069 ( .I1(B[16]), .I2(A[21]), .O(n7700) );
  INV_GATE U8070 ( .I1(n7700), .O(n7461) );
  INV_GATE U8071 ( .I1(n7192), .O(n7186) );
  NAND_GATE U8072 ( .I1(n7187), .I2(n7186), .O(n7184) );
  NAND_GATE U8073 ( .I1(n7185), .I2(n7184), .O(n7190) );
  NAND_GATE U8074 ( .I1(n7190), .I2(n7189), .O(n7195) );
  INV_GATE U8075 ( .I1(n7191), .O(n7193) );
  NAND_GATE U8076 ( .I1(n7193), .I2(n7192), .O(n7194) );
  NAND_GATE U8077 ( .I1(n7195), .I2(n7194), .O(n7696) );
  NAND_GATE U8078 ( .I1(n7461), .I2(n7696), .O(n7693) );
  NAND_GATE U8079 ( .I1(B[16]), .I2(A[20]), .O(n7717) );
  INV_GATE U8080 ( .I1(n7717), .O(n7459) );
  NAND_GATE U8081 ( .I1(n7197), .I2(n7202), .O(n7708) );
  NAND_GATE U8082 ( .I1(n7198), .I2(n784), .O(n7202) );
  NAND_GATE U8083 ( .I1(n7200), .I2(n7199), .O(n7201) );
  NAND_GATE U8084 ( .I1(n7202), .I2(n7201), .O(n7711) );
  NAND_GATE U8085 ( .I1(n7708), .I2(n7714), .O(n7203) );
  NAND_GATE U8086 ( .I1(n7710), .I2(n7203), .O(n7703) );
  NAND_GATE U8087 ( .I1(B[16]), .I2(A[19]), .O(n7723) );
  INV_GATE U8088 ( .I1(n7723), .O(n7457) );
  NAND_GATE U8089 ( .I1(B[16]), .I2(A[18]), .O(n7738) );
  INV_GATE U8090 ( .I1(n7738), .O(n7443) );
  NAND_GATE U8091 ( .I1(B[16]), .I2(A[17]), .O(n7743) );
  INV_GATE U8092 ( .I1(n7743), .O(n7748) );
  NAND_GATE U8093 ( .I1(B[16]), .I2(A[16]), .O(n8055) );
  INV_GATE U8094 ( .I1(n8055), .O(n7759) );
  NAND_GATE U8095 ( .I1(n7205), .I2(n7204), .O(n7209) );
  INV_GATE U8096 ( .I1(n7218), .O(n7208) );
  NAND3_GATE U8097 ( .I1(n7209), .I2(n7208), .I3(n7210), .O(n7214) );
  NAND_GATE U8098 ( .I1(n7210), .I2(n7209), .O(n7211) );
  NAND_GATE U8099 ( .I1(n7218), .I2(n7211), .O(n7213) );
  NAND3_GATE U8100 ( .I1(n7214), .I2(n7213), .I3(n7212), .O(n7220) );
  OR_GATE U8101 ( .I1(n7216), .I2(n7215), .O(n7219) );
  NAND3_GATE U8102 ( .I1(n7220), .I2(n7219), .I3(n277), .O(n7757) );
  NAND_GATE U8103 ( .I1(n7759), .I2(n877), .O(n7415) );
  NAND_GATE U8104 ( .I1(B[16]), .I2(A[15]), .O(n7961) );
  INV_GATE U8105 ( .I1(n7961), .O(n7411) );
  NAND_GATE U8106 ( .I1(n7221), .I2(n7230), .O(n7228) );
  NAND_GATE U8107 ( .I1(n7225), .I2(n4), .O(n7222) );
  NAND_GATE U8108 ( .I1(n7223), .I2(n7222), .O(n7227) );
  NAND3_GATE U8109 ( .I1(n7225), .I2(n4), .I3(n7224), .O(n7226) );
  NAND3_GATE U8110 ( .I1(n7228), .I2(n7227), .I3(n7226), .O(n7232) );
  NAND_GATE U8111 ( .I1(n7232), .I2(n7231), .O(n7964) );
  NAND_GATE U8112 ( .I1(n7411), .I2(n7964), .O(n7966) );
  NAND_GATE U8113 ( .I1(n294), .I2(n7239), .O(n7235) );
  NAND3_GATE U8114 ( .I1(n7235), .I2(n7234), .I3(n7233), .O(n7242) );
  OR_GATE U8115 ( .I1(n7237), .I2(n7236), .O(n7241) );
  OR_GATE U8116 ( .I1(n7239), .I2(n7238), .O(n7240) );
  NAND3_GATE U8117 ( .I1(n7242), .I2(n7241), .I3(n7240), .O(n7955) );
  NAND_GATE U8118 ( .I1(B[16]), .I2(A[14]), .O(n7957) );
  INV_GATE U8119 ( .I1(n7957), .O(n7954) );
  NAND_GATE U8120 ( .I1(n293), .I2(n7954), .O(n7952) );
  NAND_GATE U8121 ( .I1(B[16]), .I2(A[13]), .O(n7945) );
  INV_GATE U8122 ( .I1(n7945), .O(n7402) );
  NAND_GATE U8123 ( .I1(B[16]), .I2(A[12]), .O(n7767) );
  INV_GATE U8124 ( .I1(n7767), .O(n7762) );
  NAND_GATE U8125 ( .I1(n7245), .I2(n7244), .O(n7248) );
  NAND_GATE U8126 ( .I1(n7075), .I2(n7248), .O(n7246) );
  NAND_GATE U8127 ( .I1(n7252), .I2(n7246), .O(n7251) );
  INV_GATE U8128 ( .I1(n7252), .O(n7247) );
  NAND3_GATE U8129 ( .I1(n7248), .I2(n7247), .I3(n7075), .O(n7250) );
  NAND3_GATE U8130 ( .I1(n7251), .I2(n7250), .I3(n7249), .O(n7258) );
  OR_GATE U8131 ( .I1(n7253), .I2(n7252), .O(n7257) );
  OR_GATE U8132 ( .I1(n7255), .I2(n7254), .O(n7256) );
  NAND_GATE U8133 ( .I1(n7762), .I2(n793), .O(n7770) );
  NAND_GATE U8134 ( .I1(B[16]), .I2(A[11]), .O(n7930) );
  INV_GATE U8135 ( .I1(n7930), .O(n7391) );
  NAND_GATE U8136 ( .I1(n7259), .I2(n1298), .O(n7263) );
  NAND_GATE U8137 ( .I1(n7261), .I2(n7260), .O(n7262) );
  NAND3_GATE U8138 ( .I1(n7263), .I2(n7262), .I3(n1294), .O(n7267) );
  NAND3_GATE U8139 ( .I1(n7267), .I2(n7266), .I3(n7265), .O(n7273) );
  NAND3_GATE U8140 ( .I1(n1294), .I2(n7268), .I3(n7270), .O(n7272) );
  OR_GATE U8141 ( .I1(n7270), .I2(n7269), .O(n7271) );
  NAND3_GATE U8142 ( .I1(n7273), .I2(n7272), .I3(n7271), .O(n7780) );
  INV_GATE U8143 ( .I1(n7780), .O(n7782) );
  NAND_GATE U8144 ( .I1(B[16]), .I2(A[10]), .O(n7778) );
  INV_GATE U8145 ( .I1(n7778), .O(n7777) );
  NAND_GATE U8146 ( .I1(n7782), .I2(n7777), .O(n7775) );
  NAND_GATE U8147 ( .I1(B[16]), .I2(A[8]), .O(n7797) );
  INV_GATE U8148 ( .I1(n7797), .O(n7794) );
  NAND_GATE U8149 ( .I1(n1043), .I2(n7280), .O(n7275) );
  NAND3_GATE U8150 ( .I1(n7276), .I2(n7275), .I3(n7274), .O(n7283) );
  OR_GATE U8151 ( .I1(n7278), .I2(n7277), .O(n7282) );
  OR_GATE U8152 ( .I1(n7280), .I2(n7279), .O(n7281) );
  NAND3_GATE U8153 ( .I1(n7283), .I2(n7282), .I3(n7281), .O(n7791) );
  INV_GATE U8154 ( .I1(n7791), .O(n7792) );
  NAND_GATE U8155 ( .I1(n7794), .I2(n7792), .O(n7366) );
  NAND_GATE U8156 ( .I1(B[16]), .I2(A[7]), .O(n7892) );
  INV_GATE U8157 ( .I1(n7892), .O(n7883) );
  NAND_GATE U8158 ( .I1(n1319), .I2(n7290), .O(n7286) );
  NAND3_GATE U8159 ( .I1(n7286), .I2(n7285), .I3(n7284), .O(n7293) );
  OR_GATE U8160 ( .I1(n7288), .I2(n7287), .O(n7292) );
  OR_GATE U8161 ( .I1(n7290), .I2(n7289), .O(n7291) );
  NAND3_GATE U8162 ( .I1(n7293), .I2(n7292), .I3(n7291), .O(n7804) );
  INV_GATE U8163 ( .I1(n7804), .O(n7807) );
  NAND_GATE U8164 ( .I1(B[16]), .I2(A[6]), .O(n7811) );
  INV_GATE U8165 ( .I1(n7811), .O(n7805) );
  NAND_GATE U8166 ( .I1(n7807), .I2(n7805), .O(n7802) );
  NAND_GATE U8167 ( .I1(B[16]), .I2(A[5]), .O(n7874) );
  INV_GATE U8168 ( .I1(n7874), .O(n7345) );
  OR_GATE U8169 ( .I1(n7294), .I2(n7299), .O(n7297) );
  OR_GATE U8170 ( .I1(n7298), .I2(n7295), .O(n7296) );
  AND_GATE U8171 ( .I1(n7297), .I2(n7296), .O(n7304) );
  NAND_GATE U8172 ( .I1(n1231), .I2(n7298), .O(n7302) );
  NAND3_GATE U8173 ( .I1(n7302), .I2(n7301), .I3(n7300), .O(n7303) );
  NAND_GATE U8174 ( .I1(n7304), .I2(n7303), .O(n7817) );
  NAND_GATE U8175 ( .I1(B[16]), .I2(A[4]), .O(n7823) );
  INV_GATE U8176 ( .I1(n7823), .O(n7818) );
  NAND_GATE U8177 ( .I1(n696), .I2(n7818), .O(n7814) );
  NAND_GATE U8178 ( .I1(B[16]), .I2(A[3]), .O(n7858) );
  INV_GATE U8179 ( .I1(n7858), .O(n7327) );
  NAND_GATE U8180 ( .I1(B[16]), .I2(A[2]), .O(n7837) );
  INV_GATE U8181 ( .I1(n7837), .O(n7831) );
  NAND_GATE U8182 ( .I1(n1429), .I2(A[0]), .O(n7305) );
  NAND_GATE U8183 ( .I1(n14241), .I2(n7305), .O(n7306) );
  NAND_GATE U8184 ( .I1(B[18]), .I2(n7306), .O(n7310) );
  NAND_GATE U8185 ( .I1(n1430), .I2(A[1]), .O(n7307) );
  NAND_GATE U8186 ( .I1(n724), .I2(n7307), .O(n7308) );
  NAND_GATE U8187 ( .I1(B[17]), .I2(n7308), .O(n7309) );
  NAND_GATE U8188 ( .I1(n7310), .I2(n7309), .O(n7833) );
  NAND_GATE U8189 ( .I1(n7831), .I2(n7833), .O(n7828) );
  NAND3_GATE U8190 ( .I1(B[16]), .I2(B[17]), .I3(n1254), .O(n7829) );
  INV_GATE U8191 ( .I1(n7829), .O(n7832) );
  INV_GATE U8192 ( .I1(n7833), .O(n7830) );
  NAND_GATE U8193 ( .I1(n7837), .I2(n7830), .O(n7311) );
  NAND_GATE U8194 ( .I1(n7832), .I2(n7311), .O(n7312) );
  NAND_GATE U8195 ( .I1(n7828), .I2(n7312), .O(n7857) );
  NAND_GATE U8196 ( .I1(n7327), .I2(n7857), .O(n7853) );
  OR_GATE U8197 ( .I1(n7314), .I2(n7313), .O(n7326) );
  NAND_GATE U8198 ( .I1(n7316), .I2(n7320), .O(n7324) );
  NAND_GATE U8199 ( .I1(n7318), .I2(n7317), .O(n7319) );
  NAND_GATE U8200 ( .I1(n7320), .I2(n7319), .O(n7321) );
  NAND_GATE U8201 ( .I1(n7322), .I2(n7321), .O(n7323) );
  NAND_GATE U8202 ( .I1(n7324), .I2(n7323), .O(n7325) );
  NAND_GATE U8203 ( .I1(n7326), .I2(n7325), .O(n7856) );
  NAND_GATE U8204 ( .I1(n7857), .I2(n7856), .O(n7328) );
  NAND3_GATE U8205 ( .I1(n7853), .I2(n7328), .I3(n7852), .O(n7819) );
  NAND_GATE U8206 ( .I1(n7817), .I2(n7823), .O(n7329) );
  NAND_GATE U8207 ( .I1(n7819), .I2(n7329), .O(n7330) );
  NAND_GATE U8208 ( .I1(n7814), .I2(n7330), .O(n7873) );
  NAND_GATE U8209 ( .I1(n7345), .I2(n7873), .O(n7868) );
  INV_GATE U8210 ( .I1(n7335), .O(n7332) );
  NAND_GATE U8211 ( .I1(n7333), .I2(n7332), .O(n7338) );
  NAND_GATE U8212 ( .I1(n7334), .I2(n7338), .O(n7342) );
  NAND_GATE U8213 ( .I1(n7336), .I2(n7335), .O(n7337) );
  NAND_GATE U8214 ( .I1(n7338), .I2(n7337), .O(n7339) );
  NAND_GATE U8215 ( .I1(n7340), .I2(n7339), .O(n7341) );
  NAND_GATE U8216 ( .I1(n7342), .I2(n7341), .O(n7343) );
  NAND_GATE U8217 ( .I1(n7344), .I2(n7343), .O(n7872) );
  NAND_GATE U8218 ( .I1(n7873), .I2(n7872), .O(n7346) );
  NAND_GATE U8219 ( .I1(n7345), .I2(n7872), .O(n7867) );
  NAND3_GATE U8220 ( .I1(n7868), .I2(n7346), .I3(n7867), .O(n7806) );
  NAND_GATE U8221 ( .I1(n7804), .I2(n7811), .O(n7347) );
  NAND_GATE U8222 ( .I1(n7806), .I2(n7347), .O(n7348) );
  NAND_GATE U8223 ( .I1(n7802), .I2(n7348), .O(n7887) );
  NAND_GATE U8224 ( .I1(n7883), .I2(n7887), .O(n7884) );
  INV_GATE U8225 ( .I1(n7358), .O(n7351) );
  NAND_GATE U8226 ( .I1(n7349), .I2(n7353), .O(n7356) );
  NAND_GATE U8227 ( .I1(n7352), .I2(n7351), .O(n7353) );
  NAND_GATE U8228 ( .I1(n7356), .I2(n7355), .O(n7361) );
  INV_GATE U8229 ( .I1(n7357), .O(n7359) );
  NAND_GATE U8230 ( .I1(n7359), .I2(n7358), .O(n7360) );
  NAND_GATE U8231 ( .I1(n7361), .I2(n7360), .O(n7888) );
  NAND_GATE U8232 ( .I1(n7887), .I2(n7888), .O(n7363) );
  NAND_GATE U8233 ( .I1(n7883), .I2(n7888), .O(n7362) );
  NAND3_GATE U8234 ( .I1(n7884), .I2(n7363), .I3(n7362), .O(n7793) );
  NAND_GATE U8235 ( .I1(n7797), .I2(n7791), .O(n7364) );
  NAND_GATE U8236 ( .I1(n7793), .I2(n7364), .O(n7365) );
  NAND_GATE U8237 ( .I1(n7366), .I2(n7365), .O(n7911) );
  INV_GATE U8238 ( .I1(n7371), .O(n7369) );
  NAND_GATE U8239 ( .I1(n7368), .I2(n7374), .O(n7901) );
  NAND_GATE U8240 ( .I1(n7370), .I2(n7369), .O(n7374) );
  NAND_GATE U8241 ( .I1(n7372), .I2(n7371), .O(n7373) );
  NAND_GATE U8242 ( .I1(n7374), .I2(n7373), .O(n7899) );
  NAND_GATE U8243 ( .I1(n7901), .I2(n7375), .O(n7376) );
  NAND_GATE U8244 ( .I1(n7903), .I2(n7376), .O(n7914) );
  NAND_GATE U8245 ( .I1(n7911), .I2(n7914), .O(n7378) );
  NAND_GATE U8246 ( .I1(B[16]), .I2(A[9]), .O(n7908) );
  INV_GATE U8247 ( .I1(n7908), .O(n7377) );
  NAND_GATE U8248 ( .I1(n7377), .I2(n7914), .O(n7912) );
  NAND_GATE U8249 ( .I1(n7377), .I2(n7911), .O(n7913) );
  NAND3_GATE U8250 ( .I1(n7378), .I2(n7912), .I3(n7913), .O(n7781) );
  NAND_GATE U8251 ( .I1(n7780), .I2(n7778), .O(n7379) );
  NAND_GATE U8252 ( .I1(n7781), .I2(n7379), .O(n7380) );
  NAND_GATE U8253 ( .I1(n7775), .I2(n7380), .O(n7926) );
  NAND_GATE U8254 ( .I1(n7391), .I2(n7926), .O(n7923) );
  NAND3_GATE U8255 ( .I1(n7382), .I2(n1346), .I3(n7381), .O(n7383) );
  NAND3_GATE U8256 ( .I1(n7385), .I2(n7384), .I3(n7383), .O(n7390) );
  INV_GATE U8257 ( .I1(n7386), .O(n7388) );
  NAND_GATE U8258 ( .I1(n7388), .I2(n7387), .O(n7389) );
  NAND_GATE U8259 ( .I1(n7390), .I2(n7389), .O(n7927) );
  NAND_GATE U8260 ( .I1(n7926), .I2(n7927), .O(n7392) );
  NAND_GATE U8261 ( .I1(n7391), .I2(n7927), .O(n7922) );
  NAND3_GATE U8262 ( .I1(n7923), .I2(n7392), .I3(n7922), .O(n7771) );
  NAND_GATE U8263 ( .I1(n7767), .I2(n396), .O(n7393) );
  NAND_GATE U8264 ( .I1(n7771), .I2(n7393), .O(n7394) );
  NAND_GATE U8265 ( .I1(n7770), .I2(n7394), .O(n7943) );
  NAND_GATE U8266 ( .I1(n7402), .I2(n7943), .O(n7937) );
  INV_GATE U8267 ( .I1(n7399), .O(n7396) );
  NAND_GATE U8268 ( .I1(n7397), .I2(n7396), .O(n7404) );
  NAND_GATE U8269 ( .I1(n7405), .I2(n7404), .O(n7400) );
  NAND3_GATE U8270 ( .I1(n7397), .I2(n7396), .I3(n7398), .O(n7401) );
  NAND3_GATE U8271 ( .I1(n757), .I2(n7399), .I3(n7398), .O(n7403) );
  NAND3_GATE U8272 ( .I1(n7400), .I2(n7401), .I3(n7403), .O(n7942) );
  NAND_GATE U8273 ( .I1(n7944), .I2(n7942), .O(n7940) );
  NAND_GATE U8274 ( .I1(n7943), .I2(n7940), .O(n7408) );
  AND3_GATE U8275 ( .I1(n7403), .I2(n7402), .I3(n7401), .O(n7407) );
  NAND3_GATE U8276 ( .I1(n7405), .I2(n7404), .I3(n7944), .O(n7406) );
  NAND_GATE U8277 ( .I1(n7407), .I2(n7406), .O(n7936) );
  NAND_GATE U8278 ( .I1(n7955), .I2(n7957), .O(n7409) );
  NAND_GATE U8279 ( .I1(n7956), .I2(n7409), .O(n7410) );
  NAND_GATE U8280 ( .I1(n7952), .I2(n7410), .O(n7967) );
  NAND_GATE U8281 ( .I1(n7964), .I2(n7967), .O(n7412) );
  NAND_GATE U8282 ( .I1(n7411), .I2(n7967), .O(n7965) );
  NAND3_GATE U8283 ( .I1(n7966), .I2(n7412), .I3(n7965), .O(n7758) );
  NAND_GATE U8284 ( .I1(n8055), .I2(n7757), .O(n7413) );
  NAND_GATE U8285 ( .I1(n7758), .I2(n7413), .O(n7414) );
  NAND_GATE U8286 ( .I1(n7415), .I2(n7414), .O(n7742) );
  NAND_GATE U8287 ( .I1(n7748), .I2(n7742), .O(n7746) );
  NAND_GATE U8288 ( .I1(n7418), .I2(n1290), .O(n7416) );
  NAND_GATE U8289 ( .I1(n7417), .I2(n7416), .O(n7422) );
  NAND_GATE U8290 ( .I1(n353), .I2(n7424), .O(n7421) );
  NAND3_GATE U8291 ( .I1(n7419), .I2(n1290), .I3(n7418), .O(n7420) );
  NAND3_GATE U8292 ( .I1(n7422), .I2(n7421), .I3(n7420), .O(n7427) );
  INV_GATE U8293 ( .I1(n7423), .O(n7425) );
  NAND_GATE U8294 ( .I1(n7425), .I2(n7424), .O(n7426) );
  NAND_GATE U8295 ( .I1(n7427), .I2(n7426), .O(n7749) );
  NAND_GATE U8296 ( .I1(n7748), .I2(n7749), .O(n7429) );
  NAND_GATE U8297 ( .I1(n7742), .I2(n7749), .O(n7428) );
  NAND3_GATE U8298 ( .I1(n7746), .I2(n7429), .I3(n7428), .O(n7735) );
  NAND_GATE U8299 ( .I1(n7443), .I2(n7735), .O(n7732) );
  INV_GATE U8300 ( .I1(n7436), .O(n7434) );
  NAND_GATE U8301 ( .I1(n7435), .I2(n7434), .O(n7432) );
  NAND3_GATE U8302 ( .I1(n7433), .I2(n7432), .I3(n7431), .O(n7442) );
  NAND_GATE U8303 ( .I1(n7437), .I2(n7436), .O(n7438) );
  NAND_GATE U8304 ( .I1(n7432), .I2(n7438), .O(n7439) );
  NAND_GATE U8305 ( .I1(n7440), .I2(n7439), .O(n7441) );
  NAND_GATE U8306 ( .I1(n7442), .I2(n7441), .O(n7734) );
  NAND_GATE U8307 ( .I1(n7443), .I2(n354), .O(n7731) );
  NAND_GATE U8308 ( .I1(n7735), .I2(n354), .O(n7444) );
  NAND3_GATE U8309 ( .I1(n7732), .I2(n7731), .I3(n7444), .O(n7724) );
  NAND_GATE U8310 ( .I1(n7457), .I2(n7724), .O(n7726) );
  NAND3_GATE U8311 ( .I1(n7454), .I2(n7445), .I3(n7446), .O(n7452) );
  NAND_GATE U8312 ( .I1(n7446), .I2(n7454), .O(n7447) );
  NAND_GATE U8313 ( .I1(n7448), .I2(n7447), .O(n7451) );
  NAND_GATE U8314 ( .I1(n7449), .I2(n307), .O(n7450) );
  NAND3_GATE U8315 ( .I1(n7452), .I2(n7451), .I3(n7450), .O(n7456) );
  OR_GATE U8316 ( .I1(n7454), .I2(n7453), .O(n7455) );
  NAND_GATE U8317 ( .I1(n7456), .I2(n7455), .O(n7727) );
  NAND_GATE U8318 ( .I1(n7457), .I2(n7727), .O(n7725) );
  NAND_GATE U8319 ( .I1(n7724), .I2(n7727), .O(n7458) );
  NAND3_GATE U8320 ( .I1(n7726), .I2(n7725), .I3(n7458), .O(n7716) );
  NAND_GATE U8321 ( .I1(n7459), .I2(n7716), .O(n7704) );
  NAND3_GATE U8322 ( .I1(n7705), .I2(n7704), .I3(n7460), .O(n7697) );
  NAND_GATE U8323 ( .I1(n7461), .I2(n7697), .O(n7692) );
  NAND_GATE U8324 ( .I1(n7696), .I2(n7697), .O(n7462) );
  NAND3_GATE U8325 ( .I1(n7693), .I2(n7692), .I3(n7462), .O(n7686) );
  NAND_GATE U8326 ( .I1(n7473), .I2(n7686), .O(n7682) );
  INV_GATE U8327 ( .I1(n7463), .O(n7464) );
  NAND_GATE U8328 ( .I1(n7464), .I2(n7467), .O(n7472) );
  NAND_GATE U8329 ( .I1(n7466), .I2(n7465), .O(n7470) );
  NAND_GATE U8330 ( .I1(n7470), .I2(n7469), .O(n7471) );
  NAND_GATE U8331 ( .I1(n7472), .I2(n7471), .O(n7685) );
  NAND_GATE U8332 ( .I1(n7686), .I2(n7685), .O(n7474) );
  NAND3_GATE U8333 ( .I1(n7682), .I2(n7681), .I3(n7474), .O(n7675) );
  NAND_GATE U8334 ( .I1(n7487), .I2(n7675), .O(n7671) );
  INV_GATE U8335 ( .I1(n7475), .O(n7476) );
  NAND_GATE U8336 ( .I1(n7476), .I2(n7479), .O(n7486) );
  NAND_GATE U8337 ( .I1(n7481), .I2(n809), .O(n7477) );
  NAND_GATE U8338 ( .I1(n7478), .I2(n7477), .O(n7484) );
  NAND_GATE U8339 ( .I1(n7484), .I2(n7483), .O(n7485) );
  NAND_GATE U8340 ( .I1(n7486), .I2(n7485), .O(n7674) );
  NAND_GATE U8341 ( .I1(n7487), .I2(n7674), .O(n7670) );
  NAND_GATE U8342 ( .I1(n7675), .I2(n7674), .O(n7488) );
  NAND3_GATE U8343 ( .I1(n7671), .I2(n7670), .I3(n7488), .O(n7664) );
  NAND_GATE U8344 ( .I1(n7502), .I2(n7664), .O(n7660) );
  INV_GATE U8345 ( .I1(n7489), .O(n7490) );
  NAND_GATE U8346 ( .I1(n7490), .I2(n7493), .O(n7501) );
  NAND_GATE U8347 ( .I1(n7492), .I2(n7495), .O(n7499) );
  NAND_GATE U8348 ( .I1(n833), .I2(n7493), .O(n7494) );
  NAND_GATE U8349 ( .I1(n7495), .I2(n7494), .O(n7496) );
  NAND_GATE U8350 ( .I1(n7497), .I2(n7496), .O(n7498) );
  NAND_GATE U8351 ( .I1(n7499), .I2(n7498), .O(n7500) );
  NAND_GATE U8352 ( .I1(n7501), .I2(n7500), .O(n7663) );
  NAND_GATE U8353 ( .I1(n7664), .I2(n7663), .O(n7503) );
  NAND3_GATE U8354 ( .I1(n7660), .I2(n7659), .I3(n7503), .O(n7654) );
  NAND_GATE U8355 ( .I1(n7517), .I2(n7654), .O(n7650) );
  INV_GATE U8356 ( .I1(n7504), .O(n7505) );
  NAND_GATE U8357 ( .I1(n7505), .I2(n7508), .O(n7516) );
  NAND_GATE U8358 ( .I1(n7507), .I2(n7510), .O(n7514) );
  NAND_GATE U8359 ( .I1(n910), .I2(n7508), .O(n7509) );
  NAND_GATE U8360 ( .I1(n7510), .I2(n7509), .O(n7511) );
  NAND_GATE U8361 ( .I1(n7512), .I2(n7511), .O(n7513) );
  NAND_GATE U8362 ( .I1(n7514), .I2(n7513), .O(n7515) );
  NAND_GATE U8363 ( .I1(n7516), .I2(n7515), .O(n7653) );
  NAND_GATE U8364 ( .I1(n7517), .I2(n7653), .O(n7649) );
  NAND_GATE U8365 ( .I1(n7654), .I2(n7653), .O(n7518) );
  NAND3_GATE U8366 ( .I1(n7650), .I2(n7649), .I3(n7518), .O(n7644) );
  NAND_GATE U8367 ( .I1(n7532), .I2(n7644), .O(n7640) );
  INV_GATE U8368 ( .I1(n7519), .O(n7520) );
  NAND_GATE U8369 ( .I1(n7520), .I2(n7523), .O(n7531) );
  NAND_GATE U8370 ( .I1(n7522), .I2(n7525), .O(n7529) );
  NAND_GATE U8371 ( .I1(n938), .I2(n7523), .O(n7524) );
  NAND_GATE U8372 ( .I1(n7525), .I2(n7524), .O(n7526) );
  NAND_GATE U8373 ( .I1(n7527), .I2(n7526), .O(n7528) );
  NAND_GATE U8374 ( .I1(n7529), .I2(n7528), .O(n7530) );
  NAND_GATE U8375 ( .I1(n7531), .I2(n7530), .O(n7643) );
  NAND_GATE U8376 ( .I1(n7532), .I2(n7643), .O(n7639) );
  NAND_GATE U8377 ( .I1(n7644), .I2(n7643), .O(n7533) );
  NAND3_GATE U8378 ( .I1(n7640), .I2(n7639), .I3(n7533), .O(n7634) );
  NAND_GATE U8379 ( .I1(n7547), .I2(n7634), .O(n7630) );
  INV_GATE U8380 ( .I1(n7534), .O(n7535) );
  NAND_GATE U8381 ( .I1(n7535), .I2(n7538), .O(n7546) );
  NAND_GATE U8382 ( .I1(n7537), .I2(n7540), .O(n7544) );
  NAND_GATE U8383 ( .I1(n318), .I2(n7538), .O(n7539) );
  NAND_GATE U8384 ( .I1(n7540), .I2(n7539), .O(n7541) );
  NAND_GATE U8385 ( .I1(n7542), .I2(n7541), .O(n7543) );
  NAND_GATE U8386 ( .I1(n7544), .I2(n7543), .O(n7545) );
  NAND_GATE U8387 ( .I1(n7546), .I2(n7545), .O(n7633) );
  NAND_GATE U8388 ( .I1(n7547), .I2(n7633), .O(n7629) );
  NAND_GATE U8389 ( .I1(n7634), .I2(n7633), .O(n7548) );
  NAND3_GATE U8390 ( .I1(n7630), .I2(n7629), .I3(n7548), .O(n7623) );
  NAND_GATE U8391 ( .I1(n7564), .I2(n7623), .O(n7619) );
  INV_GATE U8392 ( .I1(n7549), .O(n7550) );
  NAND_GATE U8393 ( .I1(n7550), .I2(n7554), .O(n7563) );
  INV_GATE U8394 ( .I1(n7554), .O(n7551) );
  NAND_GATE U8395 ( .I1(n7552), .I2(n7551), .O(n7557) );
  NAND_GATE U8396 ( .I1(n7553), .I2(n7557), .O(n7561) );
  NAND_GATE U8397 ( .I1(n7555), .I2(n7554), .O(n7556) );
  NAND_GATE U8398 ( .I1(n7557), .I2(n7556), .O(n7558) );
  NAND_GATE U8399 ( .I1(n7559), .I2(n7558), .O(n7560) );
  NAND_GATE U8400 ( .I1(n7561), .I2(n7560), .O(n7562) );
  NAND_GATE U8401 ( .I1(n7563), .I2(n7562), .O(n7622) );
  NAND_GATE U8402 ( .I1(n7564), .I2(n7622), .O(n7618) );
  NAND_GATE U8403 ( .I1(n7623), .I2(n7622), .O(n7565) );
  NAND3_GATE U8404 ( .I1(n7619), .I2(n7618), .I3(n7565), .O(n7612) );
  NAND_GATE U8405 ( .I1(n7581), .I2(n7612), .O(n7608) );
  INV_GATE U8406 ( .I1(n7566), .O(n7567) );
  NAND_GATE U8407 ( .I1(n7567), .I2(n7571), .O(n7580) );
  INV_GATE U8408 ( .I1(n7571), .O(n7568) );
  NAND_GATE U8409 ( .I1(n7569), .I2(n7568), .O(n7574) );
  NAND_GATE U8410 ( .I1(n7570), .I2(n7574), .O(n7578) );
  NAND_GATE U8411 ( .I1(n7572), .I2(n7571), .O(n7573) );
  NAND_GATE U8412 ( .I1(n7574), .I2(n7573), .O(n7575) );
  NAND_GATE U8413 ( .I1(n7576), .I2(n7575), .O(n7577) );
  NAND_GATE U8414 ( .I1(n7578), .I2(n7577), .O(n7579) );
  NAND_GATE U8415 ( .I1(n7580), .I2(n7579), .O(n7611) );
  NAND_GATE U8416 ( .I1(n7581), .I2(n7611), .O(n7607) );
  NAND_GATE U8417 ( .I1(n7612), .I2(n7611), .O(n7582) );
  NAND3_GATE U8418 ( .I1(n7608), .I2(n7607), .I3(n7582), .O(n7601) );
  NAND_GATE U8419 ( .I1(n7601), .I2(n7600), .O(n7584) );
  NAND_GATE U8420 ( .I1(n7583), .I2(n7601), .O(n7596) );
  AND3_GATE U8421 ( .I1(n7595), .I2(n7584), .I3(n7596), .O(n7591) );
  NAND_GATE U8422 ( .I1(n1428), .I2(A[31]), .O(n7590) );
  NAND_GATE U8423 ( .I1(n7591), .I2(n7590), .O(n7585) );
  NAND_GATE U8424 ( .I1(n7589), .I2(n7585), .O(n7594) );
  NAND_GATE U8425 ( .I1(n14808), .I2(n7594), .O(n7588) );
  INV_GATE U8426 ( .I1(n7594), .O(n14807) );
  NAND_GATE U8427 ( .I1(n7586), .I2(n14807), .O(n7587) );
  NAND_GATE U8428 ( .I1(n7588), .I2(n7587), .O(\A1[46] ) );
  INV_GATE U8429 ( .I1(n7589), .O(n7592) );
  NAND3_GATE U8430 ( .I1(n7592), .I2(n7591), .I3(n7590), .O(n7593) );
  NAND_GATE U8431 ( .I1(n7594), .I2(n7593), .O(n8003) );
  INV_GATE U8432 ( .I1(n8003), .O(n14810) );
  OR_GATE U8433 ( .I1(n7595), .I2(n7601), .O(n7598) );
  OR_GATE U8434 ( .I1(n7600), .I2(n7596), .O(n7597) );
  AND_GATE U8435 ( .I1(n7598), .I2(n7597), .O(n7606) );
  INV_GATE U8436 ( .I1(n7601), .O(n7599) );
  NAND_GATE U8437 ( .I1(n7599), .I2(n7600), .O(n7604) );
  NAND3_GATE U8438 ( .I1(n7604), .I2(n7603), .I3(n7602), .O(n7605) );
  OR_GATE U8439 ( .I1(n7607), .I2(n7612), .O(n7610) );
  OR_GATE U8440 ( .I1(n7611), .I2(n7608), .O(n7609) );
  AND_GATE U8441 ( .I1(n7610), .I2(n7609), .O(n7617) );
  NAND_GATE U8442 ( .I1(n990), .I2(n7611), .O(n7615) );
  NAND3_GATE U8443 ( .I1(n7615), .I2(n7614), .I3(n7613), .O(n7616) );
  NAND_GATE U8444 ( .I1(n7617), .I2(n7616), .O(n8012) );
  INV_GATE U8445 ( .I1(n8012), .O(n8015) );
  NAND_GATE U8446 ( .I1(B[15]), .I2(A[30]), .O(n8019) );
  INV_GATE U8447 ( .I1(n8019), .O(n8013) );
  NAND_GATE U8448 ( .I1(n8015), .I2(n8013), .O(n8009) );
  OR_GATE U8449 ( .I1(n7618), .I2(n7623), .O(n7621) );
  OR_GATE U8450 ( .I1(n7622), .I2(n7619), .O(n7620) );
  AND_GATE U8451 ( .I1(n7621), .I2(n7620), .O(n7628) );
  NAND_GATE U8452 ( .I1(n988), .I2(n7622), .O(n7626) );
  NAND3_GATE U8453 ( .I1(n7626), .I2(n7625), .I3(n7624), .O(n7627) );
  NAND_GATE U8454 ( .I1(n7628), .I2(n7627), .O(n8027) );
  INV_GATE U8455 ( .I1(n8027), .O(n8030) );
  NAND_GATE U8456 ( .I1(B[15]), .I2(A[29]), .O(n8034) );
  INV_GATE U8457 ( .I1(n8034), .O(n8028) );
  NAND_GATE U8458 ( .I1(n8030), .I2(n8028), .O(n8024) );
  OR_GATE U8459 ( .I1(n7629), .I2(n7634), .O(n7632) );
  OR_GATE U8460 ( .I1(n7633), .I2(n7630), .O(n7631) );
  NAND_GATE U8461 ( .I1(n983), .I2(n7633), .O(n7637) );
  NAND3_GATE U8462 ( .I1(n7637), .I2(n7636), .I3(n7635), .O(n7638) );
  NAND_GATE U8463 ( .I1(B[15]), .I2(A[28]), .O(n8427) );
  INV_GATE U8464 ( .I1(n8427), .O(n8423) );
  NAND_GATE U8465 ( .I1(n824), .I2(n8423), .O(n8420) );
  OR_GATE U8466 ( .I1(n7639), .I2(n7644), .O(n7642) );
  OR_GATE U8467 ( .I1(n7643), .I2(n7640), .O(n7641) );
  NAND_GATE U8468 ( .I1(n974), .I2(n7643), .O(n7647) );
  NAND3_GATE U8469 ( .I1(n7647), .I2(n7646), .I3(n7645), .O(n7648) );
  NAND_GATE U8470 ( .I1(B[15]), .I2(A[27]), .O(n8413) );
  INV_GATE U8471 ( .I1(n8413), .O(n8408) );
  NAND_GATE U8472 ( .I1(n763), .I2(n8408), .O(n8406) );
  OR_GATE U8473 ( .I1(n7649), .I2(n7654), .O(n7652) );
  OR_GATE U8474 ( .I1(n7653), .I2(n7650), .O(n7651) );
  NAND_GATE U8475 ( .I1(n963), .I2(n7653), .O(n7657) );
  NAND3_GATE U8476 ( .I1(n7657), .I2(n7656), .I3(n7655), .O(n7658) );
  NAND_GATE U8477 ( .I1(B[15]), .I2(A[26]), .O(n8399) );
  INV_GATE U8478 ( .I1(n8399), .O(n8394) );
  NAND_GATE U8479 ( .I1(n857), .I2(n8394), .O(n8391) );
  OR_GATE U8480 ( .I1(n7659), .I2(n7664), .O(n7662) );
  OR_GATE U8481 ( .I1(n7663), .I2(n7660), .O(n7661) );
  AND_GATE U8482 ( .I1(n7662), .I2(n7661), .O(n7669) );
  NAND_GATE U8483 ( .I1(n964), .I2(n7663), .O(n7667) );
  NAND3_GATE U8484 ( .I1(n7667), .I2(n7666), .I3(n7665), .O(n7668) );
  NAND_GATE U8485 ( .I1(n7669), .I2(n7668), .O(n8378) );
  NAND_GATE U8486 ( .I1(B[15]), .I2(A[25]), .O(n8384) );
  INV_GATE U8487 ( .I1(n8384), .O(n8379) );
  NAND_GATE U8488 ( .I1(n832), .I2(n8379), .O(n8376) );
  OR_GATE U8489 ( .I1(n7674), .I2(n7671), .O(n7672) );
  AND_GATE U8490 ( .I1(n7673), .I2(n7672), .O(n7680) );
  NAND_GATE U8491 ( .I1(n199), .I2(n7674), .O(n7678) );
  NAND3_GATE U8492 ( .I1(n7678), .I2(n7677), .I3(n7676), .O(n7679) );
  NAND_GATE U8493 ( .I1(n7680), .I2(n7679), .O(n8368) );
  INV_GATE U8494 ( .I1(n8368), .O(n8366) );
  NAND_GATE U8495 ( .I1(B[15]), .I2(A[24]), .O(n8369) );
  INV_GATE U8496 ( .I1(n8369), .O(n8364) );
  NAND_GATE U8497 ( .I1(n8366), .I2(n8364), .O(n8361) );
  OR_GATE U8498 ( .I1(n7681), .I2(n7686), .O(n7684) );
  OR_GATE U8499 ( .I1(n7685), .I2(n7682), .O(n7683) );
  AND_GATE U8500 ( .I1(n7684), .I2(n7683), .O(n7691) );
  NAND_GATE U8501 ( .I1(n955), .I2(n7685), .O(n7689) );
  NAND3_GATE U8502 ( .I1(n7689), .I2(n7688), .I3(n7687), .O(n7690) );
  NAND_GATE U8503 ( .I1(n7691), .I2(n7690), .O(n8351) );
  NAND_GATE U8504 ( .I1(B[15]), .I2(A[23]), .O(n8354) );
  INV_GATE U8505 ( .I1(n8354), .O(n8349) );
  NAND_GATE U8506 ( .I1(n701), .I2(n8349), .O(n8346) );
  NAND_GATE U8507 ( .I1(B[15]), .I2(A[22]), .O(n8336) );
  INV_GATE U8508 ( .I1(n8336), .O(n8332) );
  OR_GATE U8509 ( .I1(n7692), .I2(n7696), .O(n7695) );
  AND_GATE U8510 ( .I1(n7695), .I2(n7694), .O(n7702) );
  NAND_GATE U8511 ( .I1(n7696), .I2(n956), .O(n7699) );
  NAND3_GATE U8512 ( .I1(n7700), .I2(n7699), .I3(n7698), .O(n7701) );
  NAND_GATE U8513 ( .I1(n7702), .I2(n7701), .O(n8334) );
  NAND_GATE U8514 ( .I1(n8332), .I2(n590), .O(n8339) );
  NAND_GATE U8515 ( .I1(B[15]), .I2(A[21]), .O(n8320) );
  OR_GATE U8516 ( .I1(n7704), .I2(n7703), .O(n7707) );
  OR_GATE U8517 ( .I1(n7716), .I2(n7705), .O(n7706) );
  INV_GATE U8518 ( .I1(n7708), .O(n7709) );
  NAND_GATE U8519 ( .I1(n7710), .I2(n7709), .O(n7713) );
  NAND_GATE U8520 ( .I1(n7712), .I2(n7711), .O(n7714) );
  NAND3_GATE U8521 ( .I1(n7713), .I2(n309), .I3(n7714), .O(n7719) );
  NAND_GATE U8522 ( .I1(n7714), .I2(n7713), .O(n7715) );
  NAND_GATE U8523 ( .I1(n7716), .I2(n7715), .O(n7718) );
  NAND3_GATE U8524 ( .I1(n7719), .I2(n7718), .I3(n7717), .O(n7720) );
  NAND_GATE U8525 ( .I1(B[15]), .I2(A[20]), .O(n8308) );
  INV_GATE U8526 ( .I1(n8308), .O(n8306) );
  NAND_GATE U8527 ( .I1(n7724), .I2(n306), .O(n7722) );
  NAND3_GATE U8528 ( .I1(n7723), .I2(n7722), .I3(n7721), .O(n7730) );
  OR_GATE U8529 ( .I1(n7725), .I2(n7724), .O(n7729) );
  OR_GATE U8530 ( .I1(n7727), .I2(n7726), .O(n7728) );
  NAND3_GATE U8531 ( .I1(n7730), .I2(n7729), .I3(n7728), .O(n8310) );
  INV_GATE U8532 ( .I1(n8310), .O(n8307) );
  NAND_GATE U8533 ( .I1(n8306), .I2(n8307), .O(n8314) );
  NAND_GATE U8534 ( .I1(B[15]), .I2(A[19]), .O(n8559) );
  INV_GATE U8535 ( .I1(n8559), .O(n8039) );
  OR_GATE U8536 ( .I1(n7731), .I2(n7735), .O(n7741) );
  INV_GATE U8537 ( .I1(n7732), .O(n7733) );
  NAND_GATE U8538 ( .I1(n7733), .I2(n7734), .O(n7740) );
  NAND_GATE U8539 ( .I1(n7735), .I2(n7734), .O(n7737) );
  NAND3_GATE U8540 ( .I1(n7738), .I2(n7737), .I3(n7736), .O(n7739) );
  NAND3_GATE U8541 ( .I1(n7741), .I2(n7740), .I3(n7739), .O(n8043) );
  NAND_GATE U8542 ( .I1(n8039), .I2(n8041), .O(n7980) );
  NAND_GATE U8543 ( .I1(B[15]), .I2(A[18]), .O(n8569) );
  INV_GATE U8544 ( .I1(n8569), .O(n8052) );
  NAND_GATE U8545 ( .I1(n7742), .I2(n714), .O(n7745) );
  INV_GATE U8546 ( .I1(n7742), .O(n7750) );
  NAND_GATE U8547 ( .I1(n7750), .I2(n7749), .O(n7744) );
  NAND3_GATE U8548 ( .I1(n7745), .I2(n7744), .I3(n7743), .O(n7753) );
  INV_GATE U8549 ( .I1(n7746), .O(n7747) );
  NAND_GATE U8550 ( .I1(n7747), .I2(n714), .O(n7752) );
  NAND3_GATE U8551 ( .I1(n7750), .I2(n7749), .I3(n7748), .O(n7751) );
  NAND3_GATE U8552 ( .I1(n7753), .I2(n7752), .I3(n7751), .O(n8048) );
  NAND_GATE U8553 ( .I1(n8052), .I2(n8050), .O(n7977) );
  NAND_GATE U8554 ( .I1(B[15]), .I2(A[17]), .O(n8063) );
  INV_GATE U8555 ( .I1(n8063), .O(n7973) );
  NAND_GATE U8556 ( .I1(n877), .I2(n7758), .O(n7755) );
  INV_GATE U8557 ( .I1(n7758), .O(n7756) );
  NAND_GATE U8558 ( .I1(n7757), .I2(n7756), .O(n7754) );
  NAND_GATE U8559 ( .I1(n7755), .I2(n7754), .O(n8054) );
  NAND_GATE U8560 ( .I1(n7759), .I2(n7754), .O(n8056) );
  NAND_GATE U8561 ( .I1(n8060), .I2(n8056), .O(n7760) );
  NAND3_GATE U8562 ( .I1(n7759), .I2(n7758), .I3(n877), .O(n8057) );
  NAND_GATE U8563 ( .I1(n7760), .I2(n8057), .O(n8066) );
  NAND_GATE U8564 ( .I1(B[15]), .I2(A[16]), .O(n8594) );
  INV_GATE U8565 ( .I1(n8594), .O(n8078) );
  NAND_GATE U8566 ( .I1(B[15]), .I2(A[14]), .O(n8273) );
  INV_GATE U8567 ( .I1(n8273), .O(n8266) );
  INV_GATE U8568 ( .I1(n7771), .O(n7763) );
  NAND_GATE U8569 ( .I1(n396), .I2(n7763), .O(n7761) );
  NAND_GATE U8570 ( .I1(n7762), .I2(n7761), .O(n7769) );
  NAND_GATE U8571 ( .I1(n793), .I2(n7771), .O(n7765) );
  NAND_GATE U8572 ( .I1(n7765), .I2(n7764), .O(n7766) );
  NAND_GATE U8573 ( .I1(n7767), .I2(n7766), .O(n7768) );
  NAND_GATE U8574 ( .I1(n7769), .I2(n7768), .O(n7774) );
  INV_GATE U8575 ( .I1(n7770), .O(n7772) );
  NAND_GATE U8576 ( .I1(n7772), .I2(n7771), .O(n7773) );
  NAND_GATE U8577 ( .I1(n7774), .I2(n7773), .O(n8255) );
  NAND3_GATE U8578 ( .I1(A[13]), .I2(n8255), .I3(B[15]), .O(n8259) );
  NAND_GATE U8579 ( .I1(B[15]), .I2(A[12]), .O(n8248) );
  INV_GATE U8580 ( .I1(n8248), .O(n8084) );
  NAND_GATE U8581 ( .I1(B[15]), .I2(A[11]), .O(n8240) );
  INV_GATE U8582 ( .I1(n8240), .O(n7920) );
  INV_GATE U8583 ( .I1(n7781), .O(n7779) );
  NAND_GATE U8584 ( .I1(n7780), .I2(n7779), .O(n7776) );
  NAND_GATE U8585 ( .I1(n7777), .I2(n7776), .O(n7785) );
  NAND3_GATE U8586 ( .I1(n7780), .I2(n7779), .I3(n7778), .O(n7784) );
  NAND_GATE U8587 ( .I1(n7782), .I2(n7781), .O(n7783) );
  NAND3_GATE U8588 ( .I1(n7785), .I2(n7784), .I3(n7783), .O(n7786) );
  NAND_GATE U8589 ( .I1(n7787), .I2(n7786), .O(n8237) );
  NAND_GATE U8590 ( .I1(n7920), .I2(n8237), .O(n8233) );
  NAND_GATE U8591 ( .I1(B[15]), .I2(A[10]), .O(n8227) );
  INV_GATE U8592 ( .I1(n8227), .O(n8093) );
  INV_GATE U8593 ( .I1(n7793), .O(n7790) );
  NAND_GATE U8594 ( .I1(n7791), .I2(n7790), .O(n7788) );
  NAND_GATE U8595 ( .I1(n7789), .I2(n7788), .O(n7796) );
  NAND_GATE U8596 ( .I1(n7794), .I2(n7788), .O(n7799) );
  INV_GATE U8597 ( .I1(n7799), .O(n7795) );
  NAND3_GATE U8598 ( .I1(n7794), .I2(n7793), .I3(n7792), .O(n7801) );
  NAND_GATE U8599 ( .I1(n7795), .I2(n7801), .O(n8214) );
  NAND_GATE U8600 ( .I1(B[15]), .I2(A[9]), .O(n8217) );
  INV_GATE U8601 ( .I1(n8217), .O(n7897) );
  NAND3_GATE U8602 ( .I1(n7798), .I2(n8214), .I3(n7897), .O(n8212) );
  NAND_GATE U8603 ( .I1(n7797), .I2(n7796), .O(n7798) );
  NAND_GATE U8604 ( .I1(n7799), .I2(n7798), .O(n7800) );
  NAND_GATE U8605 ( .I1(n7801), .I2(n7800), .O(n8220) );
  NAND_GATE U8606 ( .I1(B[15]), .I2(A[8]), .O(n8105) );
  INV_GATE U8607 ( .I1(n8105), .O(n8108) );
  INV_GATE U8608 ( .I1(n7806), .O(n7803) );
  NAND_GATE U8609 ( .I1(n7804), .I2(n7803), .O(n7809) );
  NAND_GATE U8610 ( .I1(n7805), .I2(n7809), .O(n7813) );
  NAND_GATE U8611 ( .I1(n7807), .I2(n7806), .O(n7808) );
  NAND_GATE U8612 ( .I1(n7809), .I2(n7808), .O(n7810) );
  NAND_GATE U8613 ( .I1(n7811), .I2(n7810), .O(n7812) );
  NAND_GATE U8614 ( .I1(n7813), .I2(n7812), .O(n8203) );
  NAND_GATE U8615 ( .I1(n8202), .I2(n8203), .O(n8200) );
  NAND_GATE U8616 ( .I1(B[15]), .I2(A[6]), .O(n8124) );
  INV_GATE U8617 ( .I1(n8124), .O(n8118) );
  NAND_GATE U8618 ( .I1(B[15]), .I2(A[5]), .O(n8187) );
  INV_GATE U8619 ( .I1(n8187), .O(n7865) );
  INV_GATE U8620 ( .I1(n7814), .O(n7815) );
  NAND_GATE U8621 ( .I1(n7815), .I2(n7819), .O(n7827) );
  INV_GATE U8622 ( .I1(n7819), .O(n7816) );
  NAND_GATE U8623 ( .I1(n7817), .I2(n7816), .O(n7821) );
  NAND_GATE U8624 ( .I1(n7818), .I2(n7821), .O(n7825) );
  NAND_GATE U8625 ( .I1(n696), .I2(n7819), .O(n7820) );
  NAND_GATE U8626 ( .I1(n7821), .I2(n7820), .O(n7822) );
  NAND_GATE U8627 ( .I1(n7823), .I2(n7822), .O(n7824) );
  NAND_GATE U8628 ( .I1(n7825), .I2(n7824), .O(n7826) );
  NAND_GATE U8629 ( .I1(n7827), .I2(n7826), .O(n8185) );
  NAND_GATE U8630 ( .I1(n7865), .I2(n8185), .O(n8182) );
  NAND_GATE U8631 ( .I1(B[15]), .I2(A[4]), .O(n8138) );
  INV_GATE U8632 ( .I1(n8138), .O(n8132) );
  NAND_GATE U8633 ( .I1(B[15]), .I2(A[3]), .O(n8173) );
  INV_GATE U8634 ( .I1(n8173), .O(n7850) );
  OR_GATE U8635 ( .I1(n7829), .I2(n7828), .O(n7841) );
  NAND_GATE U8636 ( .I1(n7830), .I2(n7829), .O(n7835) );
  NAND_GATE U8637 ( .I1(n7831), .I2(n7835), .O(n7839) );
  NAND_GATE U8638 ( .I1(n7833), .I2(n7832), .O(n7834) );
  NAND_GATE U8639 ( .I1(n7835), .I2(n7834), .O(n7836) );
  NAND_GATE U8640 ( .I1(n7837), .I2(n7836), .O(n7838) );
  NAND_GATE U8641 ( .I1(n7839), .I2(n7838), .O(n7840) );
  NAND_GATE U8642 ( .I1(n7841), .I2(n7840), .O(n8171) );
  NAND_GATE U8643 ( .I1(n7850), .I2(n8171), .O(n8168) );
  NAND_GATE U8644 ( .I1(B[15]), .I2(A[2]), .O(n8152) );
  INV_GATE U8645 ( .I1(n8152), .O(n8146) );
  NAND_GATE U8646 ( .I1(n1428), .I2(A[0]), .O(n7842) );
  NAND_GATE U8647 ( .I1(n14241), .I2(n7842), .O(n7843) );
  NAND_GATE U8648 ( .I1(B[17]), .I2(n7843), .O(n7847) );
  NAND_GATE U8649 ( .I1(n1429), .I2(A[1]), .O(n7844) );
  NAND_GATE U8650 ( .I1(n724), .I2(n7844), .O(n7845) );
  NAND_GATE U8651 ( .I1(B[16]), .I2(n7845), .O(n7846) );
  NAND_GATE U8652 ( .I1(n7847), .I2(n7846), .O(n8148) );
  NAND_GATE U8653 ( .I1(n8146), .I2(n8148), .O(n8143) );
  NAND3_GATE U8654 ( .I1(B[15]), .I2(B[16]), .I3(n1254), .O(n8144) );
  INV_GATE U8655 ( .I1(n8144), .O(n8147) );
  INV_GATE U8656 ( .I1(n8148), .O(n8145) );
  NAND_GATE U8657 ( .I1(n8152), .I2(n8145), .O(n7848) );
  NAND_GATE U8658 ( .I1(n8147), .I2(n7848), .O(n7849) );
  NAND_GATE U8659 ( .I1(n8143), .I2(n7849), .O(n8172) );
  NAND_GATE U8660 ( .I1(n8171), .I2(n8172), .O(n7851) );
  NAND_GATE U8661 ( .I1(n7850), .I2(n8172), .O(n8167) );
  NAND3_GATE U8662 ( .I1(n8168), .I2(n7851), .I3(n8167), .O(n8134) );
  NAND_GATE U8663 ( .I1(n8132), .I2(n8134), .O(n8129) );
  OR_GATE U8664 ( .I1(n7852), .I2(n7857), .O(n7855) );
  OR_GATE U8665 ( .I1(n7856), .I2(n7853), .O(n7854) );
  AND_GATE U8666 ( .I1(n7855), .I2(n7854), .O(n7862) );
  NAND_GATE U8667 ( .I1(n1236), .I2(n7856), .O(n7860) );
  NAND3_GATE U8668 ( .I1(n7860), .I2(n7859), .I3(n7858), .O(n7861) );
  NAND_GATE U8669 ( .I1(n7862), .I2(n7861), .O(n8130) );
  INV_GATE U8670 ( .I1(n8130), .O(n8133) );
  INV_GATE U8671 ( .I1(n8134), .O(n8131) );
  NAND_GATE U8672 ( .I1(n8138), .I2(n8131), .O(n7863) );
  NAND_GATE U8673 ( .I1(n8133), .I2(n7863), .O(n7864) );
  NAND_GATE U8674 ( .I1(n8129), .I2(n7864), .O(n8186) );
  NAND_GATE U8675 ( .I1(n8185), .I2(n8186), .O(n7866) );
  NAND_GATE U8676 ( .I1(n7865), .I2(n8186), .O(n8181) );
  NAND3_GATE U8677 ( .I1(n8182), .I2(n7866), .I3(n8181), .O(n8120) );
  NAND_GATE U8678 ( .I1(n8118), .I2(n8120), .O(n8115) );
  OR_GATE U8679 ( .I1(n7872), .I2(n7868), .O(n7869) );
  AND_GATE U8680 ( .I1(n7870), .I2(n7869), .O(n7878) );
  INV_GATE U8681 ( .I1(n7873), .O(n7871) );
  NAND_GATE U8682 ( .I1(n7871), .I2(n7872), .O(n7876) );
  NAND_GATE U8683 ( .I1(n7873), .I2(n1315), .O(n7875) );
  NAND3_GATE U8684 ( .I1(n7876), .I2(n7875), .I3(n7874), .O(n7877) );
  NAND_GATE U8685 ( .I1(n7878), .I2(n7877), .O(n8116) );
  INV_GATE U8686 ( .I1(n8116), .O(n8119) );
  INV_GATE U8687 ( .I1(n8120), .O(n8117) );
  NAND_GATE U8688 ( .I1(n8124), .I2(n8117), .O(n7879) );
  NAND_GATE U8689 ( .I1(n8119), .I2(n7879), .O(n7880) );
  NAND_GATE U8690 ( .I1(n8115), .I2(n7880), .O(n8201) );
  NAND_GATE U8691 ( .I1(n8200), .I2(n8201), .O(n7882) );
  NAND_GATE U8692 ( .I1(B[15]), .I2(A[7]), .O(n8204) );
  INV_GATE U8693 ( .I1(n8204), .O(n7881) );
  NAND_GATE U8694 ( .I1(n7881), .I2(n8201), .O(n8195) );
  NAND_GATE U8695 ( .I1(n7881), .I2(n8200), .O(n8196) );
  NAND3_GATE U8696 ( .I1(n7882), .I2(n8195), .I3(n8196), .O(n8102) );
  NAND_GATE U8697 ( .I1(n8108), .I2(n8102), .O(n8111) );
  INV_GATE U8698 ( .I1(n7887), .O(n7889) );
  NAND3_GATE U8699 ( .I1(n7889), .I2(n7883), .I3(n7888), .O(n7886) );
  OR_GATE U8700 ( .I1(n7888), .I2(n7884), .O(n7885) );
  AND_GATE U8701 ( .I1(n7886), .I2(n7885), .O(n7894) );
  NAND_GATE U8702 ( .I1(n7889), .I2(n7888), .O(n7890) );
  NAND3_GATE U8703 ( .I1(n7892), .I2(n7891), .I3(n7890), .O(n7893) );
  NAND_GATE U8704 ( .I1(n7894), .I2(n7893), .O(n8112) );
  INV_GATE U8705 ( .I1(n8112), .O(n8101) );
  INV_GATE U8706 ( .I1(n8102), .O(n8106) );
  NAND_GATE U8707 ( .I1(n8105), .I2(n8106), .O(n7895) );
  NAND_GATE U8708 ( .I1(n8101), .I2(n7895), .O(n7896) );
  NAND_GATE U8709 ( .I1(n8111), .I2(n7896), .O(n8216) );
  NAND_GATE U8710 ( .I1(n8220), .I2(n8216), .O(n7898) );
  NAND_GATE U8711 ( .I1(n7897), .I2(n8216), .O(n8221) );
  NAND3_GATE U8712 ( .I1(n8212), .I2(n7898), .I3(n8221), .O(n8099) );
  NAND_GATE U8713 ( .I1(n8093), .I2(n8099), .O(n8094) );
  NAND_GATE U8714 ( .I1(n7900), .I2(n7899), .O(n7905) );
  INV_GATE U8715 ( .I1(n7911), .O(n7904) );
  INV_GATE U8716 ( .I1(n7901), .O(n7902) );
  NAND_GATE U8717 ( .I1(n7903), .I2(n7902), .O(n7906) );
  NAND3_GATE U8718 ( .I1(n7905), .I2(n7904), .I3(n7906), .O(n7910) );
  NAND_GATE U8719 ( .I1(n7906), .I2(n7905), .O(n7907) );
  NAND_GATE U8720 ( .I1(n7911), .I2(n7907), .O(n7909) );
  NAND3_GATE U8721 ( .I1(n7910), .I2(n7909), .I3(n7908), .O(n7917) );
  OR_GATE U8722 ( .I1(n7912), .I2(n7911), .O(n7916) );
  OR_GATE U8723 ( .I1(n7914), .I2(n7913), .O(n7915) );
  NAND3_GATE U8724 ( .I1(n7917), .I2(n7916), .I3(n7915), .O(n8096) );
  INV_GATE U8725 ( .I1(n8096), .O(n8098) );
  INV_GATE U8726 ( .I1(n8099), .O(n8097) );
  NAND_GATE U8727 ( .I1(n8227), .I2(n8097), .O(n7918) );
  NAND_GATE U8728 ( .I1(n8098), .I2(n7918), .O(n7919) );
  NAND_GATE U8729 ( .I1(n8094), .I2(n7919), .O(n8238) );
  NAND_GATE U8730 ( .I1(n8237), .I2(n8238), .O(n7921) );
  NAND_GATE U8731 ( .I1(n7920), .I2(n8238), .O(n8232) );
  NAND3_GATE U8732 ( .I1(n8233), .I2(n7921), .I3(n8232), .O(n8088) );
  NAND_GATE U8733 ( .I1(n8084), .I2(n8088), .O(n8085) );
  OR_GATE U8734 ( .I1(n7922), .I2(n7926), .O(n7925) );
  OR_GATE U8735 ( .I1(n7927), .I2(n7923), .O(n7924) );
  NAND_GATE U8736 ( .I1(n1032), .I2(n7927), .O(n7928) );
  NAND3_GATE U8737 ( .I1(n7930), .I2(n7929), .I3(n7928), .O(n7931) );
  INV_GATE U8738 ( .I1(n8089), .O(n8087) );
  INV_GATE U8739 ( .I1(n8088), .O(n8090) );
  NAND_GATE U8740 ( .I1(n8248), .I2(n8090), .O(n7932) );
  NAND_GATE U8741 ( .I1(n8087), .I2(n7932), .O(n7933) );
  NAND_GATE U8742 ( .I1(n8085), .I2(n7933), .O(n8260) );
  NAND_GATE U8743 ( .I1(n8255), .I2(n8260), .O(n7935) );
  NAND_GATE U8744 ( .I1(B[15]), .I2(A[13]), .O(n8258) );
  INV_GATE U8745 ( .I1(n8258), .O(n7934) );
  NAND_GATE U8746 ( .I1(n8260), .I2(n7934), .O(n8254) );
  NAND3_GATE U8747 ( .I1(n8259), .I2(n7935), .I3(n8254), .O(n8269) );
  NAND_GATE U8748 ( .I1(n8266), .I2(n8269), .O(n8276) );
  OR_GATE U8749 ( .I1(n7936), .I2(n7943), .O(n7939) );
  OR_GATE U8750 ( .I1(n7940), .I2(n7937), .O(n7938) );
  AND_GATE U8751 ( .I1(n7939), .I2(n7938), .O(n7949) );
  INV_GATE U8752 ( .I1(n7943), .O(n7941) );
  NAND_GATE U8753 ( .I1(n7941), .I2(n7940), .O(n7947) );
  NAND3_GATE U8754 ( .I1(n7944), .I2(n7943), .I3(n7942), .O(n7946) );
  NAND3_GATE U8755 ( .I1(n7947), .I2(n7946), .I3(n7945), .O(n7948) );
  NAND_GATE U8756 ( .I1(n7949), .I2(n7948), .O(n8267) );
  INV_GATE U8757 ( .I1(n8267), .O(n8277) );
  NAND_GATE U8758 ( .I1(n8273), .I2(n8268), .O(n7950) );
  NAND_GATE U8759 ( .I1(n8277), .I2(n7950), .O(n7951) );
  NAND_GATE U8760 ( .I1(n8276), .I2(n7951), .O(n8288) );
  NAND_GATE U8761 ( .I1(n7955), .I2(n761), .O(n7953) );
  NAND_GATE U8762 ( .I1(n7954), .I2(n7953), .O(n7958) );
  NAND_GATE U8763 ( .I1(n8289), .I2(n8287), .O(n8285) );
  NAND_GATE U8764 ( .I1(n8288), .I2(n8285), .O(n7960) );
  NAND_GATE U8765 ( .I1(B[15]), .I2(A[15]), .O(n8290) );
  INV_GATE U8766 ( .I1(n8290), .O(n8281) );
  NAND_GATE U8767 ( .I1(n8281), .I2(n8285), .O(n7959) );
  NAND_GATE U8768 ( .I1(n8281), .I2(n8288), .O(n8282) );
  NAND3_GATE U8769 ( .I1(n7960), .I2(n7959), .I3(n8282), .O(n8073) );
  NAND_GATE U8770 ( .I1(n8078), .I2(n8073), .O(n8079) );
  NAND3_GATE U8771 ( .I1(n7963), .I2(n7962), .I3(n7961), .O(n7970) );
  OR_GATE U8772 ( .I1(n7965), .I2(n7964), .O(n7969) );
  OR_GATE U8773 ( .I1(n7967), .I2(n7966), .O(n7968) );
  NAND3_GATE U8774 ( .I1(n7970), .I2(n7969), .I3(n7968), .O(n8076) );
  INV_GATE U8775 ( .I1(n8076), .O(n8080) );
  INV_GATE U8776 ( .I1(n8073), .O(n8077) );
  NAND_GATE U8777 ( .I1(n8594), .I2(n8077), .O(n7971) );
  NAND_GATE U8778 ( .I1(n8080), .I2(n7971), .O(n7972) );
  NAND_GATE U8779 ( .I1(n8079), .I2(n7972), .O(n8069) );
  NAND_GATE U8780 ( .I1(n8066), .I2(n8069), .O(n7974) );
  NAND_GATE U8781 ( .I1(n7973), .I2(n8069), .O(n8067) );
  NAND_GATE U8782 ( .I1(n8569), .I2(n8048), .O(n7975) );
  NAND_GATE U8783 ( .I1(n8051), .I2(n7975), .O(n7976) );
  NAND_GATE U8784 ( .I1(n7977), .I2(n7976), .O(n8040) );
  NAND_GATE U8785 ( .I1(n8559), .I2(n8043), .O(n7978) );
  NAND_GATE U8786 ( .I1(n8040), .I2(n7978), .O(n7979) );
  NAND_GATE U8787 ( .I1(n7980), .I2(n7979), .O(n8315) );
  NAND_GATE U8788 ( .I1(n8308), .I2(n8310), .O(n7981) );
  NAND_GATE U8789 ( .I1(n8315), .I2(n7981), .O(n7982) );
  NAND_GATE U8790 ( .I1(n8314), .I2(n7982), .O(n8326) );
  NAND_GATE U8791 ( .I1(n8320), .I2(n8322), .O(n7983) );
  NAND_GATE U8792 ( .I1(n8336), .I2(n8334), .O(n7984) );
  NAND_GATE U8793 ( .I1(n8340), .I2(n7984), .O(n7985) );
  NAND_GATE U8794 ( .I1(n8339), .I2(n7985), .O(n8350) );
  NAND_GATE U8795 ( .I1(n8351), .I2(n8354), .O(n7986) );
  NAND_GATE U8796 ( .I1(n8350), .I2(n7986), .O(n7987) );
  NAND_GATE U8797 ( .I1(n8346), .I2(n7987), .O(n8365) );
  NAND_GATE U8798 ( .I1(n8368), .I2(n8369), .O(n7988) );
  NAND_GATE U8799 ( .I1(n8365), .I2(n7988), .O(n7989) );
  NAND_GATE U8800 ( .I1(n8361), .I2(n7989), .O(n8380) );
  NAND_GATE U8801 ( .I1(n8378), .I2(n8384), .O(n7990) );
  NAND_GATE U8802 ( .I1(n8380), .I2(n7990), .O(n7991) );
  NAND_GATE U8803 ( .I1(n8376), .I2(n7991), .O(n8395) );
  NAND_GATE U8804 ( .I1(n8393), .I2(n8399), .O(n7992) );
  NAND_GATE U8805 ( .I1(n8395), .I2(n7992), .O(n7993) );
  NAND_GATE U8806 ( .I1(n8391), .I2(n7993), .O(n8409) );
  NAND_GATE U8807 ( .I1(n8409), .I2(n7994), .O(n7995) );
  NAND_GATE U8808 ( .I1(n8406), .I2(n7995), .O(n8424) );
  NAND_GATE U8809 ( .I1(n8422), .I2(n8427), .O(n7996) );
  NAND_GATE U8810 ( .I1(n8424), .I2(n7996), .O(n7997) );
  NAND_GATE U8811 ( .I1(n8420), .I2(n7997), .O(n8029) );
  NAND_GATE U8812 ( .I1(n8027), .I2(n8034), .O(n7998) );
  NAND_GATE U8813 ( .I1(n8029), .I2(n7998), .O(n7999) );
  NAND_GATE U8814 ( .I1(n8024), .I2(n7999), .O(n8014) );
  NAND_GATE U8815 ( .I1(n8012), .I2(n8019), .O(n8000) );
  NAND_GATE U8816 ( .I1(n8014), .I2(n8000), .O(n8002) );
  NAND_GATE U8817 ( .I1(n1427), .I2(A[31]), .O(n8001) );
  NAND3_GATE U8818 ( .I1(n8009), .I2(n8002), .I3(n8001), .O(n8006) );
  NAND_GATE U8819 ( .I1(n404), .I2(n8006), .O(n8008) );
  NAND_GATE U8820 ( .I1(n14810), .I2(n8008), .O(n8005) );
  INV_GATE U8821 ( .I1(n8008), .O(n14809) );
  NAND_GATE U8822 ( .I1(n8003), .I2(n14809), .O(n8004) );
  NAND_GATE U8823 ( .I1(n8005), .I2(n8004), .O(\A1[45] ) );
  NAND_GATE U8824 ( .I1(n8008), .I2(n8007), .O(n8437) );
  INV_GATE U8825 ( .I1(n8437), .O(n14812) );
  INV_GATE U8826 ( .I1(n8009), .O(n8010) );
  NAND_GATE U8827 ( .I1(n8010), .I2(n8014), .O(n8023) );
  INV_GATE U8828 ( .I1(n8014), .O(n8011) );
  NAND_GATE U8829 ( .I1(n8012), .I2(n8011), .O(n8017) );
  NAND_GATE U8830 ( .I1(n8013), .I2(n8017), .O(n8021) );
  NAND_GATE U8831 ( .I1(n8015), .I2(n8014), .O(n8016) );
  NAND_GATE U8832 ( .I1(n8017), .I2(n8016), .O(n8018) );
  NAND_GATE U8833 ( .I1(n8019), .I2(n8018), .O(n8020) );
  NAND_GATE U8834 ( .I1(n8021), .I2(n8020), .O(n8022) );
  NAND_GATE U8835 ( .I1(n8023), .I2(n8022), .O(n8440) );
  NAND_GATE U8836 ( .I1(n1425), .I2(A[30]), .O(n8451) );
  INV_GATE U8837 ( .I1(n8451), .O(n8434) );
  INV_GATE U8838 ( .I1(n8024), .O(n8025) );
  NAND_GATE U8839 ( .I1(n8025), .I2(n8029), .O(n8038) );
  INV_GATE U8840 ( .I1(n8029), .O(n8026) );
  NAND_GATE U8841 ( .I1(n8027), .I2(n8026), .O(n8032) );
  NAND_GATE U8842 ( .I1(n8028), .I2(n8032), .O(n8036) );
  NAND_GATE U8843 ( .I1(n8030), .I2(n8029), .O(n8031) );
  NAND_GATE U8844 ( .I1(n8032), .I2(n8031), .O(n8033) );
  NAND_GATE U8845 ( .I1(n8034), .I2(n8033), .O(n8035) );
  NAND_GATE U8846 ( .I1(n8036), .I2(n8035), .O(n8037) );
  NAND_GATE U8847 ( .I1(n8038), .I2(n8037), .O(n8449) );
  NAND_GATE U8848 ( .I1(n8434), .I2(n8449), .O(n8445) );
  NAND_GATE U8849 ( .I1(n1425), .I2(A[29]), .O(n8462) );
  INV_GATE U8850 ( .I1(n8462), .O(n8432) );
  NAND_GATE U8851 ( .I1(n1425), .I2(A[28]), .O(n8472) );
  INV_GATE U8852 ( .I1(n8472), .O(n8418) );
  NAND_GATE U8853 ( .I1(n1425), .I2(A[27]), .O(n8482) );
  INV_GATE U8854 ( .I1(n8482), .O(n8404) );
  NAND_GATE U8855 ( .I1(n1425), .I2(A[26]), .O(n8493) );
  INV_GATE U8856 ( .I1(n8493), .O(n8389) );
  NAND_GATE U8857 ( .I1(n1425), .I2(A[25]), .O(n8504) );
  INV_GATE U8858 ( .I1(n8504), .O(n8374) );
  NAND_GATE U8859 ( .I1(n1425), .I2(A[24]), .O(n8515) );
  INV_GATE U8860 ( .I1(n8515), .O(n8359) );
  NAND_GATE U8861 ( .I1(n1425), .I2(A[23]), .O(n8527) );
  INV_GATE U8862 ( .I1(n8527), .O(n8344) );
  NAND_GATE U8863 ( .I1(n1425), .I2(A[22]), .O(n8538) );
  INV_GATE U8864 ( .I1(n8538), .O(n8329) );
  NAND_GATE U8865 ( .I1(n1425), .I2(A[21]), .O(n8549) );
  INV_GATE U8866 ( .I1(n8549), .O(n8541) );
  NAND_GATE U8867 ( .I1(n1425), .I2(A[20]), .O(n8565) );
  INV_GATE U8868 ( .I1(n8565), .O(n8303) );
  NAND3_GATE U8869 ( .I1(n8039), .I2(n8040), .I3(n8041), .O(n8557) );
  INV_GATE U8870 ( .I1(n8040), .O(n8042) );
  NAND_GATE U8871 ( .I1(n8039), .I2(n8044), .O(n8555) );
  NAND_GATE U8872 ( .I1(n8041), .I2(n8040), .O(n8045) );
  NAND_GATE U8873 ( .I1(n8043), .I2(n8042), .O(n8044) );
  NAND_GATE U8874 ( .I1(n8045), .I2(n8044), .O(n8558) );
  NAND_GATE U8875 ( .I1(n8555), .I2(n8561), .O(n8046) );
  NAND_GATE U8876 ( .I1(n8557), .I2(n8046), .O(n8552) );
  NAND_GATE U8877 ( .I1(n1425), .I2(A[19]), .O(n8579) );
  INV_GATE U8878 ( .I1(n8579), .O(n8301) );
  NAND_GATE U8879 ( .I1(n8050), .I2(n8051), .O(n8047) );
  NAND_GATE U8880 ( .I1(n8049), .I2(n8047), .O(n8568) );
  NAND_GATE U8881 ( .I1(n8048), .I2(n1283), .O(n8049) );
  NAND_GATE U8882 ( .I1(n8052), .I2(n8049), .O(n8570) );
  NAND_GATE U8883 ( .I1(n8576), .I2(n8570), .O(n8053) );
  NAND3_GATE U8884 ( .I1(n8052), .I2(n8051), .I3(n8050), .O(n8571) );
  NAND_GATE U8885 ( .I1(n8053), .I2(n8571), .O(n8582) );
  NAND_GATE U8886 ( .I1(n8301), .I2(n8582), .O(n8580) );
  NAND_GATE U8887 ( .I1(n1425), .I2(A[18]), .O(n8587) );
  INV_GATE U8888 ( .I1(n8587), .O(n8841) );
  NAND_GATE U8889 ( .I1(n8055), .I2(n8054), .O(n8060) );
  INV_GATE U8890 ( .I1(n8069), .O(n8059) );
  INV_GATE U8891 ( .I1(n8056), .O(n8058) );
  NAND_GATE U8892 ( .I1(n8058), .I2(n8057), .O(n8061) );
  NAND3_GATE U8893 ( .I1(n8060), .I2(n8059), .I3(n8061), .O(n8065) );
  NAND_GATE U8894 ( .I1(n8061), .I2(n8060), .O(n8062) );
  NAND_GATE U8895 ( .I1(n8069), .I2(n8062), .O(n8064) );
  NAND3_GATE U8896 ( .I1(n8065), .I2(n8064), .I3(n8063), .O(n8072) );
  OR_GATE U8897 ( .I1(n8067), .I2(n8066), .O(n8071) );
  OR_GATE U8898 ( .I1(n8069), .I2(n8068), .O(n8070) );
  NAND3_GATE U8899 ( .I1(n8072), .I2(n8071), .I3(n8070), .O(n8590) );
  NAND_GATE U8900 ( .I1(n8841), .I2(n876), .O(n8588) );
  NAND_GATE U8901 ( .I1(n1425), .I2(A[17]), .O(n8600) );
  INV_GATE U8902 ( .I1(n8600), .O(n8297) );
  NAND_GATE U8903 ( .I1(n8073), .I2(n8080), .O(n8075) );
  NAND_GATE U8904 ( .I1(n8077), .I2(n8076), .O(n8074) );
  NAND_GATE U8905 ( .I1(n8075), .I2(n8074), .O(n8593) );
  INV_GATE U8906 ( .I1(n8079), .O(n8081) );
  NAND_GATE U8907 ( .I1(n8081), .I2(n8080), .O(n8595) );
  NAND_GATE U8908 ( .I1(n8082), .I2(n8595), .O(n8605) );
  NAND_GATE U8909 ( .I1(n1425), .I2(A[16]), .O(n8940) );
  INV_GATE U8910 ( .I1(n8940), .O(n8833) );
  NAND_GATE U8911 ( .I1(n1425), .I2(A[14]), .O(n8623) );
  INV_GATE U8912 ( .I1(n8623), .O(n8610) );
  NAND_GATE U8913 ( .I1(n8090), .I2(n8089), .O(n8083) );
  NAND_GATE U8914 ( .I1(n8084), .I2(n8083), .O(n8249) );
  INV_GATE U8915 ( .I1(n8085), .O(n8086) );
  NAND_GATE U8916 ( .I1(n8086), .I2(n8087), .O(n8251) );
  NAND_GATE U8917 ( .I1(n8088), .I2(n8087), .O(n8091) );
  NAND_GATE U8918 ( .I1(n8091), .I2(n8083), .O(n8247) );
  NAND_GATE U8919 ( .I1(n8248), .I2(n8247), .O(n8798) );
  NAND4_GATE U8920 ( .I1(A[13]), .I2(n8797), .I3(n1425), .I4(n8798), .O(n8803)
         );
  NAND_GATE U8921 ( .I1(n1425), .I2(A[12]), .O(n8788) );
  INV_GATE U8922 ( .I1(n8788), .O(n8782) );
  NAND_GATE U8923 ( .I1(n8097), .I2(n8096), .O(n8092) );
  INV_GATE U8924 ( .I1(n8094), .O(n8095) );
  NAND_GATE U8925 ( .I1(n8095), .I2(n8098), .O(n8229) );
  NAND_GATE U8926 ( .I1(n1392), .I2(n8229), .O(n8768) );
  NAND_GATE U8927 ( .I1(n8099), .I2(n8098), .O(n8100) );
  NAND_GATE U8928 ( .I1(n8092), .I2(n8100), .O(n8226) );
  NAND_GATE U8929 ( .I1(n8227), .I2(n8226), .O(n8767) );
  NAND4_GATE U8930 ( .I1(A[11]), .I2(n8768), .I3(n1425), .I4(n8767), .O(n8774)
         );
  NAND_GATE U8931 ( .I1(n1425), .I2(A[10]), .O(n8757) );
  INV_GATE U8932 ( .I1(n8757), .O(n8632) );
  NAND_GATE U8933 ( .I1(n8102), .I2(n8101), .O(n8103) );
  NAND_GATE U8934 ( .I1(n8103), .I2(n8107), .O(n8104) );
  NAND_GATE U8935 ( .I1(n8105), .I2(n8104), .O(n8110) );
  NAND_GATE U8936 ( .I1(n8106), .I2(n8112), .O(n8107) );
  NAND_GATE U8937 ( .I1(n8108), .I2(n8107), .O(n8109) );
  NAND_GATE U8938 ( .I1(n8110), .I2(n8109), .O(n8114) );
  OR_GATE U8939 ( .I1(n8112), .I2(n8111), .O(n8113) );
  NAND_GATE U8940 ( .I1(n8114), .I2(n8113), .O(n8745) );
  NAND_GATE U8941 ( .I1(n1425), .I2(A[8]), .O(n8643) );
  INV_GATE U8942 ( .I1(n8643), .O(n8638) );
  NAND_GATE U8943 ( .I1(n1425), .I2(A[7]), .O(n8735) );
  INV_GATE U8944 ( .I1(n8735), .O(n8193) );
  OR_GATE U8945 ( .I1(n8116), .I2(n8115), .O(n8128) );
  NAND_GATE U8946 ( .I1(n8117), .I2(n8116), .O(n8122) );
  NAND_GATE U8947 ( .I1(n8118), .I2(n8122), .O(n8126) );
  NAND_GATE U8948 ( .I1(n8120), .I2(n8119), .O(n8121) );
  NAND_GATE U8949 ( .I1(n8122), .I2(n8121), .O(n8123) );
  NAND_GATE U8950 ( .I1(n8124), .I2(n8123), .O(n8125) );
  NAND_GATE U8951 ( .I1(n8126), .I2(n8125), .O(n8127) );
  NAND_GATE U8952 ( .I1(n8128), .I2(n8127), .O(n8733) );
  NAND_GATE U8953 ( .I1(n1425), .I2(A[6]), .O(n8657) );
  INV_GATE U8954 ( .I1(n8657), .O(n8651) );
  NAND_GATE U8955 ( .I1(n1425), .I2(A[5]), .O(n8721) );
  INV_GATE U8956 ( .I1(n8721), .O(n8179) );
  OR_GATE U8957 ( .I1(n8130), .I2(n8129), .O(n8142) );
  NAND_GATE U8958 ( .I1(n8131), .I2(n8130), .O(n8136) );
  NAND_GATE U8959 ( .I1(n8132), .I2(n8136), .O(n8140) );
  NAND_GATE U8960 ( .I1(n8134), .I2(n8133), .O(n8135) );
  NAND_GATE U8961 ( .I1(n8136), .I2(n8135), .O(n8137) );
  NAND_GATE U8962 ( .I1(n8138), .I2(n8137), .O(n8139) );
  NAND_GATE U8963 ( .I1(n8140), .I2(n8139), .O(n8141) );
  NAND_GATE U8964 ( .I1(n8142), .I2(n8141), .O(n8719) );
  NAND_GATE U8965 ( .I1(n8179), .I2(n8719), .O(n8716) );
  NAND_GATE U8966 ( .I1(n1425), .I2(A[4]), .O(n8671) );
  INV_GATE U8967 ( .I1(n8671), .O(n8665) );
  NAND_GATE U8968 ( .I1(n1425), .I2(A[3]), .O(n8706) );
  INV_GATE U8969 ( .I1(n8706), .O(n8165) );
  OR_GATE U8970 ( .I1(n8144), .I2(n8143), .O(n8156) );
  NAND_GATE U8971 ( .I1(n8145), .I2(n8144), .O(n8150) );
  NAND_GATE U8972 ( .I1(n8146), .I2(n8150), .O(n8154) );
  NAND_GATE U8973 ( .I1(n8148), .I2(n8147), .O(n8149) );
  NAND_GATE U8974 ( .I1(n8150), .I2(n8149), .O(n8151) );
  NAND_GATE U8975 ( .I1(n8152), .I2(n8151), .O(n8153) );
  NAND_GATE U8976 ( .I1(n8154), .I2(n8153), .O(n8155) );
  NAND_GATE U8977 ( .I1(n8156), .I2(n8155), .O(n8704) );
  NAND_GATE U8978 ( .I1(n8165), .I2(n8704), .O(n8701) );
  NAND_GATE U8979 ( .I1(n1425), .I2(A[2]), .O(n8685) );
  INV_GATE U8980 ( .I1(n8685), .O(n8679) );
  NAND3_GATE U8981 ( .I1(B[14]), .I2(B[15]), .I3(n1254), .O(n8678) );
  INV_GATE U8982 ( .I1(n8678), .O(n8681) );
  NAND_GATE U8983 ( .I1(n8679), .I2(n8681), .O(n8676) );
  NAND_GATE U8984 ( .I1(n1427), .I2(A[0]), .O(n8157) );
  NAND_GATE U8985 ( .I1(n14241), .I2(n8157), .O(n8158) );
  NAND_GATE U8986 ( .I1(B[16]), .I2(n8158), .O(n8162) );
  NAND_GATE U8987 ( .I1(n1428), .I2(A[1]), .O(n8159) );
  NAND_GATE U8988 ( .I1(n724), .I2(n8159), .O(n8160) );
  NAND_GATE U8989 ( .I1(B[15]), .I2(n8160), .O(n8161) );
  NAND_GATE U8990 ( .I1(n8162), .I2(n8161), .O(n8680) );
  NAND_GATE U8991 ( .I1(n8685), .I2(n8678), .O(n8163) );
  NAND_GATE U8992 ( .I1(n8680), .I2(n8163), .O(n8164) );
  NAND_GATE U8993 ( .I1(n8676), .I2(n8164), .O(n8705) );
  NAND_GATE U8994 ( .I1(n8704), .I2(n8705), .O(n8166) );
  NAND_GATE U8995 ( .I1(n8165), .I2(n8705), .O(n8700) );
  NAND3_GATE U8996 ( .I1(n8701), .I2(n8166), .I3(n8700), .O(n8667) );
  NAND_GATE U8997 ( .I1(n8665), .I2(n8667), .O(n8662) );
  OR_GATE U8998 ( .I1(n8167), .I2(n8171), .O(n8170) );
  OR_GATE U8999 ( .I1(n8172), .I2(n8168), .O(n8169) );
  NAND_GATE U9000 ( .I1(n8171), .I2(n1237), .O(n8175) );
  NAND3_GATE U9001 ( .I1(n8175), .I2(n8174), .I3(n8173), .O(n8176) );
  INV_GATE U9002 ( .I1(n8663), .O(n8666) );
  INV_GATE U9003 ( .I1(n8667), .O(n8664) );
  NAND_GATE U9004 ( .I1(n8671), .I2(n8664), .O(n8177) );
  NAND_GATE U9005 ( .I1(n8666), .I2(n8177), .O(n8178) );
  NAND_GATE U9006 ( .I1(n8662), .I2(n8178), .O(n8720) );
  NAND_GATE U9007 ( .I1(n8719), .I2(n8720), .O(n8180) );
  NAND_GATE U9008 ( .I1(n8179), .I2(n8720), .O(n8715) );
  NAND3_GATE U9009 ( .I1(n8716), .I2(n8180), .I3(n8715), .O(n8653) );
  NAND_GATE U9010 ( .I1(n8651), .I2(n8653), .O(n8648) );
  OR_GATE U9011 ( .I1(n8181), .I2(n8185), .O(n8184) );
  OR_GATE U9012 ( .I1(n8186), .I2(n8182), .O(n8183) );
  NAND_GATE U9013 ( .I1(n8185), .I2(n1134), .O(n8189) );
  NAND3_GATE U9014 ( .I1(n8189), .I2(n8188), .I3(n8187), .O(n8190) );
  INV_GATE U9015 ( .I1(n8649), .O(n8652) );
  INV_GATE U9016 ( .I1(n8653), .O(n8650) );
  NAND_GATE U9017 ( .I1(n8657), .I2(n8650), .O(n8191) );
  NAND_GATE U9018 ( .I1(n8652), .I2(n8191), .O(n8192) );
  NAND_GATE U9019 ( .I1(n8648), .I2(n8192), .O(n8734) );
  NAND_GATE U9020 ( .I1(n8733), .I2(n8734), .O(n8194) );
  NAND_GATE U9021 ( .I1(n8193), .I2(n8734), .O(n8729) );
  NAND3_GATE U9022 ( .I1(n8730), .I2(n8194), .I3(n8729), .O(n8639) );
  NAND_GATE U9023 ( .I1(n8638), .I2(n8639), .O(n8635) );
  OR_GATE U9024 ( .I1(n8195), .I2(n8200), .O(n8198) );
  OR_GATE U9025 ( .I1(n8201), .I2(n8196), .O(n8197) );
  AND_GATE U9026 ( .I1(n8198), .I2(n8197), .O(n8208) );
  INV_GATE U9027 ( .I1(n8201), .O(n8199) );
  NAND_GATE U9028 ( .I1(n8200), .I2(n8199), .O(n8206) );
  NAND3_GATE U9029 ( .I1(n8203), .I2(n8202), .I3(n8201), .O(n8205) );
  NAND3_GATE U9030 ( .I1(n8206), .I2(n8205), .I3(n8204), .O(n8207) );
  NAND_GATE U9031 ( .I1(n8208), .I2(n8207), .O(n8636) );
  INV_GATE U9032 ( .I1(n8639), .O(n8637) );
  NAND_GATE U9033 ( .I1(n8745), .I2(n8750), .O(n8211) );
  NAND_GATE U9034 ( .I1(n1425), .I2(A[9]), .O(n8748) );
  INV_GATE U9035 ( .I1(n8748), .O(n8210) );
  NAND_GATE U9036 ( .I1(n8750), .I2(n8210), .O(n8744) );
  NAND3_GATE U9037 ( .I1(n8749), .I2(n8211), .I3(n8744), .O(n8627) );
  NAND_GATE U9038 ( .I1(n8632), .I2(n8627), .O(n8769) );
  OR_GATE U9039 ( .I1(n8216), .I2(n8212), .O(n8224) );
  INV_GATE U9040 ( .I1(n8216), .O(n8213) );
  NAND3_GATE U9041 ( .I1(n8213), .I2(n7798), .I3(n8214), .O(n8219) );
  NAND_GATE U9042 ( .I1(n7798), .I2(n8214), .O(n8215) );
  NAND_GATE U9043 ( .I1(n8216), .I2(n8215), .O(n8218) );
  NAND3_GATE U9044 ( .I1(n8219), .I2(n8218), .I3(n8217), .O(n8223) );
  OR_GATE U9045 ( .I1(n8221), .I2(n8220), .O(n8222) );
  NAND3_GATE U9046 ( .I1(n8224), .I2(n8223), .I3(n8222), .O(n8630) );
  INV_GATE U9047 ( .I1(n8630), .O(n8633) );
  INV_GATE U9048 ( .I1(n8627), .O(n8631) );
  NAND_GATE U9049 ( .I1(n8757), .I2(n8631), .O(n8225) );
  NAND_GATE U9050 ( .I1(n8633), .I2(n8225), .O(n8770) );
  NAND_GATE U9051 ( .I1(n8769), .I2(n8770), .O(n8775) );
  NAND_GATE U9052 ( .I1(n8229), .I2(n8228), .O(n8764) );
  NAND_GATE U9053 ( .I1(n8775), .I2(n8764), .O(n8231) );
  NAND_GATE U9054 ( .I1(n1425), .I2(A[11]), .O(n8773) );
  INV_GATE U9055 ( .I1(n8773), .O(n8230) );
  NAND_GATE U9056 ( .I1(n8775), .I2(n8230), .O(n8765) );
  NAND3_GATE U9057 ( .I1(n8774), .I2(n8231), .I3(n8765), .O(n8784) );
  NAND_GATE U9058 ( .I1(n8782), .I2(n8784), .O(n8791) );
  OR_GATE U9059 ( .I1(n8232), .I2(n8237), .O(n8235) );
  OR_GATE U9060 ( .I1(n8238), .I2(n8233), .O(n8234) );
  AND_GATE U9061 ( .I1(n8235), .I2(n8234), .O(n8244) );
  INV_GATE U9062 ( .I1(n8238), .O(n8236) );
  NAND_GATE U9063 ( .I1(n8237), .I2(n8236), .O(n8242) );
  INV_GATE U9064 ( .I1(n8237), .O(n8239) );
  NAND_GATE U9065 ( .I1(n8239), .I2(n8238), .O(n8241) );
  NAND3_GATE U9066 ( .I1(n8242), .I2(n8241), .I3(n8240), .O(n8243) );
  NAND_GATE U9067 ( .I1(n8244), .I2(n8243), .O(n8792) );
  NAND_GATE U9068 ( .I1(n8788), .I2(n8783), .O(n8245) );
  NAND_GATE U9069 ( .I1(n1297), .I2(n8245), .O(n8246) );
  NAND_GATE U9070 ( .I1(n8791), .I2(n8246), .O(n8804) );
  NAND_GATE U9071 ( .I1(n8249), .I2(n8798), .O(n8250) );
  NAND_GATE U9072 ( .I1(n8251), .I2(n8250), .O(n8805) );
  NAND_GATE U9073 ( .I1(n8804), .I2(n8805), .O(n8253) );
  NAND_GATE U9074 ( .I1(n1425), .I2(A[13]), .O(n8802) );
  INV_GATE U9075 ( .I1(n8802), .O(n8252) );
  NAND_GATE U9076 ( .I1(n8804), .I2(n8252), .O(n8806) );
  NAND3_GATE U9077 ( .I1(n8803), .I2(n8253), .I3(n8806), .O(n8615) );
  NAND_GATE U9078 ( .I1(n8610), .I2(n8615), .O(n8611) );
  OR_GATE U9079 ( .I1(n8254), .I2(n8255), .O(n8263) );
  NAND_GATE U9080 ( .I1(n8255), .I2(n1002), .O(n8256) );
  NAND3_GATE U9081 ( .I1(n8258), .I2(n8257), .I3(n8256), .O(n8262) );
  OR_GATE U9082 ( .I1(n8260), .I2(n8259), .O(n8261) );
  NAND3_GATE U9083 ( .I1(n8263), .I2(n8262), .I3(n8261), .O(n8616) );
  INV_GATE U9084 ( .I1(n8616), .O(n8614) );
  NAND_GATE U9085 ( .I1(n8623), .I2(n8617), .O(n8264) );
  NAND_GATE U9086 ( .I1(n8614), .I2(n8264), .O(n8265) );
  NAND_GATE U9087 ( .I1(n8611), .I2(n8265), .O(n8820) );
  NAND_GATE U9088 ( .I1(n8266), .I2(n8271), .O(n8275) );
  NAND_GATE U9089 ( .I1(n8268), .I2(n8267), .O(n8271) );
  NAND_GATE U9090 ( .I1(n8271), .I2(n8270), .O(n8272) );
  NAND_GATE U9091 ( .I1(n8273), .I2(n8272), .O(n8274) );
  NAND_GATE U9092 ( .I1(n8275), .I2(n8274), .O(n8818) );
  INV_GATE U9093 ( .I1(n8276), .O(n8278) );
  NAND_GATE U9094 ( .I1(n8278), .I2(n8277), .O(n8819) );
  NAND_GATE U9095 ( .I1(n8818), .I2(n8819), .O(n8821) );
  NAND_GATE U9096 ( .I1(n8820), .I2(n8821), .O(n8280) );
  NAND_GATE U9097 ( .I1(n1425), .I2(A[15]), .O(n8825) );
  INV_GATE U9098 ( .I1(n8825), .O(n8815) );
  NAND_GATE U9099 ( .I1(n8821), .I2(n8815), .O(n8279) );
  NAND_GATE U9100 ( .I1(n8820), .I2(n8815), .O(n8814) );
  NAND_GATE U9101 ( .I1(n8833), .I2(n395), .O(n8834) );
  INV_GATE U9102 ( .I1(n8288), .O(n8286) );
  NAND3_GATE U9103 ( .I1(n8286), .I2(n8281), .I3(n8285), .O(n8284) );
  OR_GATE U9104 ( .I1(n8285), .I2(n8282), .O(n8283) );
  AND_GATE U9105 ( .I1(n8284), .I2(n8283), .O(n8294) );
  NAND_GATE U9106 ( .I1(n8286), .I2(n8285), .O(n8292) );
  NAND3_GATE U9107 ( .I1(n8289), .I2(n8288), .I3(n8287), .O(n8291) );
  NAND3_GATE U9108 ( .I1(n8292), .I2(n8291), .I3(n8290), .O(n8293) );
  NAND_GATE U9109 ( .I1(n8294), .I2(n8293), .O(n8832) );
  NAND_GATE U9110 ( .I1(n8940), .I2(n1386), .O(n8295) );
  NAND_GATE U9111 ( .I1(n292), .I2(n8295), .O(n8296) );
  NAND_GATE U9112 ( .I1(n8834), .I2(n8296), .O(n8604) );
  NAND_GATE U9113 ( .I1(n8605), .I2(n8604), .O(n8298) );
  NAND_GATE U9114 ( .I1(n8297), .I2(n8604), .O(n8606) );
  NAND3_GATE U9115 ( .I1(n8603), .I2(n8298), .I3(n8606), .O(n8589) );
  NAND_GATE U9116 ( .I1(n8587), .I2(n8590), .O(n8299) );
  NAND_GATE U9117 ( .I1(n8589), .I2(n8299), .O(n8300) );
  NAND_GATE U9118 ( .I1(n8588), .I2(n8300), .O(n8581) );
  NAND_GATE U9119 ( .I1(n8582), .I2(n8581), .O(n8302) );
  NAND_GATE U9120 ( .I1(n8301), .I2(n8581), .O(n8583) );
  NAND3_GATE U9121 ( .I1(n8580), .I2(n8302), .I3(n8583), .O(n8564) );
  NAND_GATE U9122 ( .I1(n8552), .I2(n8564), .O(n8304) );
  NAND_GATE U9123 ( .I1(n8303), .I2(n8564), .O(n8553) );
  NAND3_GATE U9124 ( .I1(n8554), .I2(n8304), .I3(n8553), .O(n8544) );
  NAND_GATE U9125 ( .I1(n8541), .I2(n8544), .O(n8540) );
  INV_GATE U9126 ( .I1(n8315), .O(n8309) );
  NAND_GATE U9127 ( .I1(n8310), .I2(n8309), .O(n8305) );
  NAND_GATE U9128 ( .I1(n8306), .I2(n8305), .O(n8313) );
  NAND_GATE U9129 ( .I1(n8307), .I2(n8315), .O(n8312) );
  NAND3_GATE U9130 ( .I1(n8310), .I2(n8309), .I3(n8308), .O(n8311) );
  NAND3_GATE U9131 ( .I1(n8313), .I2(n8312), .I3(n8311), .O(n8317) );
  NAND_GATE U9132 ( .I1(n8317), .I2(n8316), .O(n8545) );
  NAND_GATE U9133 ( .I1(n8544), .I2(n8545), .O(n8319) );
  NAND_GATE U9134 ( .I1(n8541), .I2(n8545), .O(n8318) );
  NAND3_GATE U9135 ( .I1(n8540), .I2(n8319), .I3(n8318), .O(n8534) );
  NAND_GATE U9136 ( .I1(n8329), .I2(n8534), .O(n8531) );
  INV_GATE U9137 ( .I1(n8326), .O(n8321) );
  NAND3_GATE U9138 ( .I1(n8322), .I2(n8321), .I3(n8320), .O(n8323) );
  NAND3_GATE U9139 ( .I1(n8325), .I2(n8324), .I3(n8323), .O(n8328) );
  NAND_GATE U9140 ( .I1(n1289), .I2(n8326), .O(n8327) );
  NAND_GATE U9141 ( .I1(n8328), .I2(n8327), .O(n8535) );
  NAND_GATE U9142 ( .I1(n8329), .I2(n8535), .O(n8530) );
  NAND_GATE U9143 ( .I1(n8534), .I2(n8535), .O(n8330) );
  NAND3_GATE U9144 ( .I1(n8531), .I2(n8530), .I3(n8330), .O(n8524) );
  NAND_GATE U9145 ( .I1(n8344), .I2(n8524), .O(n8520) );
  INV_GATE U9146 ( .I1(n8340), .O(n8333) );
  NAND_GATE U9147 ( .I1(n8334), .I2(n8333), .O(n8331) );
  NAND_GATE U9148 ( .I1(n8332), .I2(n8331), .O(n8338) );
  NAND_GATE U9149 ( .I1(n590), .I2(n8340), .O(n8335) );
  NAND_GATE U9150 ( .I1(n8338), .I2(n8337), .O(n8343) );
  INV_GATE U9151 ( .I1(n8339), .O(n8341) );
  NAND_GATE U9152 ( .I1(n8341), .I2(n8340), .O(n8342) );
  NAND_GATE U9153 ( .I1(n8343), .I2(n8342), .O(n8523) );
  NAND_GATE U9154 ( .I1(n8344), .I2(n8523), .O(n8519) );
  NAND_GATE U9155 ( .I1(n8524), .I2(n8523), .O(n8345) );
  NAND3_GATE U9156 ( .I1(n8520), .I2(n8519), .I3(n8345), .O(n8514) );
  NAND_GATE U9157 ( .I1(n8359), .I2(n8514), .O(n8510) );
  INV_GATE U9158 ( .I1(n8346), .O(n8347) );
  NAND_GATE U9159 ( .I1(n8347), .I2(n8350), .O(n8358) );
  NAND_GATE U9160 ( .I1(n8351), .I2(n305), .O(n8348) );
  NAND_GATE U9161 ( .I1(n8349), .I2(n8348), .O(n8356) );
  NAND_GATE U9162 ( .I1(n701), .I2(n8350), .O(n8352) );
  NAND_GATE U9163 ( .I1(n8352), .I2(n8348), .O(n8353) );
  NAND_GATE U9164 ( .I1(n8354), .I2(n8353), .O(n8355) );
  NAND_GATE U9165 ( .I1(n8356), .I2(n8355), .O(n8357) );
  NAND_GATE U9166 ( .I1(n8358), .I2(n8357), .O(n8513) );
  NAND_GATE U9167 ( .I1(n8514), .I2(n8513), .O(n8360) );
  NAND3_GATE U9168 ( .I1(n8510), .I2(n8509), .I3(n8360), .O(n8503) );
  NAND_GATE U9169 ( .I1(n8374), .I2(n8503), .O(n8499) );
  INV_GATE U9170 ( .I1(n8361), .O(n8362) );
  NAND_GATE U9171 ( .I1(n8362), .I2(n8365), .O(n8373) );
  INV_GATE U9172 ( .I1(n8365), .O(n8367) );
  NAND_GATE U9173 ( .I1(n8368), .I2(n8367), .O(n8363) );
  NAND_GATE U9174 ( .I1(n8364), .I2(n8363), .O(n8371) );
  NAND_GATE U9175 ( .I1(n8371), .I2(n8370), .O(n8372) );
  NAND_GATE U9176 ( .I1(n8373), .I2(n8372), .O(n8502) );
  NAND_GATE U9177 ( .I1(n8503), .I2(n8502), .O(n8375) );
  NAND3_GATE U9178 ( .I1(n8499), .I2(n8498), .I3(n8375), .O(n8492) );
  NAND_GATE U9179 ( .I1(n8389), .I2(n8492), .O(n8488) );
  INV_GATE U9180 ( .I1(n8380), .O(n8377) );
  NAND_GATE U9181 ( .I1(n8378), .I2(n8377), .O(n8382) );
  NAND_GATE U9182 ( .I1(n8379), .I2(n8382), .O(n8386) );
  NAND_GATE U9183 ( .I1(n832), .I2(n8380), .O(n8381) );
  NAND_GATE U9184 ( .I1(n8382), .I2(n8381), .O(n8383) );
  NAND_GATE U9185 ( .I1(n8384), .I2(n8383), .O(n8385) );
  NAND_GATE U9186 ( .I1(n8386), .I2(n8385), .O(n8387) );
  NAND_GATE U9187 ( .I1(n8388), .I2(n8387), .O(n8491) );
  NAND_GATE U9188 ( .I1(n8389), .I2(n8491), .O(n8487) );
  NAND_GATE U9189 ( .I1(n8492), .I2(n8491), .O(n8390) );
  NAND3_GATE U9190 ( .I1(n8488), .I2(n8487), .I3(n8390), .O(n8481) );
  NAND_GATE U9191 ( .I1(n8404), .I2(n8481), .O(n8477) );
  INV_GATE U9192 ( .I1(n8391), .O(n8392) );
  NAND_GATE U9193 ( .I1(n8392), .I2(n8395), .O(n8403) );
  NAND_GATE U9194 ( .I1(n8394), .I2(n8397), .O(n8401) );
  NAND_GATE U9195 ( .I1(n857), .I2(n8395), .O(n8396) );
  NAND_GATE U9196 ( .I1(n8397), .I2(n8396), .O(n8398) );
  NAND_GATE U9197 ( .I1(n8399), .I2(n8398), .O(n8400) );
  NAND_GATE U9198 ( .I1(n8401), .I2(n8400), .O(n8402) );
  NAND_GATE U9199 ( .I1(n8403), .I2(n8402), .O(n8480) );
  NAND_GATE U9200 ( .I1(n8481), .I2(n8480), .O(n8405) );
  NAND3_GATE U9201 ( .I1(n8477), .I2(n8476), .I3(n8405), .O(n8471) );
  NAND_GATE U9202 ( .I1(n8418), .I2(n8471), .O(n8467) );
  INV_GATE U9203 ( .I1(n8406), .O(n8407) );
  NAND_GATE U9204 ( .I1(n8407), .I2(n8409), .O(n8417) );
  NAND_GATE U9205 ( .I1(n8408), .I2(n8411), .O(n8415) );
  NAND_GATE U9206 ( .I1(n763), .I2(n8409), .O(n8410) );
  NAND_GATE U9207 ( .I1(n8411), .I2(n8410), .O(n8412) );
  NAND_GATE U9208 ( .I1(n8413), .I2(n8412), .O(n8414) );
  NAND_GATE U9209 ( .I1(n8415), .I2(n8414), .O(n8416) );
  NAND_GATE U9210 ( .I1(n8417), .I2(n8416), .O(n8470) );
  NAND_GATE U9211 ( .I1(n8418), .I2(n8470), .O(n8466) );
  NAND_GATE U9212 ( .I1(n8471), .I2(n8470), .O(n8419) );
  NAND3_GATE U9213 ( .I1(n8467), .I2(n8466), .I3(n8419), .O(n8461) );
  NAND_GATE U9214 ( .I1(n8432), .I2(n8461), .O(n8457) );
  INV_GATE U9215 ( .I1(n8420), .O(n8421) );
  NAND_GATE U9216 ( .I1(n8421), .I2(n8424), .O(n8431) );
  NAND_GATE U9217 ( .I1(n8423), .I2(n8426), .O(n8429) );
  NAND_GATE U9218 ( .I1(n824), .I2(n8424), .O(n8425) );
  NAND_GATE U9219 ( .I1(n8429), .I2(n8428), .O(n8430) );
  NAND_GATE U9220 ( .I1(n8431), .I2(n8430), .O(n8460) );
  NAND_GATE U9221 ( .I1(n8432), .I2(n8460), .O(n8456) );
  NAND_GATE U9222 ( .I1(n8461), .I2(n8460), .O(n8433) );
  NAND3_GATE U9223 ( .I1(n8457), .I2(n8456), .I3(n8433), .O(n8450) );
  NAND_GATE U9224 ( .I1(n8450), .I2(n8449), .O(n8435) );
  NAND_GATE U9225 ( .I1(n8434), .I2(n8450), .O(n8446) );
  AND3_GATE U9226 ( .I1(n8445), .I2(n8435), .I3(n8446), .O(n8442) );
  NAND_GATE U9227 ( .I1(n1426), .I2(A[31]), .O(n8441) );
  NAND_GATE U9228 ( .I1(n8442), .I2(n8441), .O(n8436) );
  NAND_GATE U9229 ( .I1(n8440), .I2(n8436), .O(n8444) );
  NAND_GATE U9230 ( .I1(n14812), .I2(n8444), .O(n8439) );
  INV_GATE U9231 ( .I1(n8444), .O(n14811) );
  NAND_GATE U9232 ( .I1(n8439), .I2(n8438), .O(\A1[44] ) );
  NAND_GATE U9233 ( .I1(n8444), .I2(n8443), .O(n8876) );
  OR_GATE U9234 ( .I1(n232), .I2(n221), .O(n8448) );
  OR_GATE U9235 ( .I1(n8449), .I2(n8446), .O(n8447) );
  AND_GATE U9236 ( .I1(n8448), .I2(n8447), .O(n8455) );
  NAND_GATE U9237 ( .I1(n989), .I2(n8449), .O(n8453) );
  NAND3_GATE U9238 ( .I1(n8453), .I2(n8452), .I3(n8451), .O(n8454) );
  NAND_GATE U9239 ( .I1(n8455), .I2(n8454), .O(n8881) );
  OR_GATE U9240 ( .I1(n8456), .I2(n8461), .O(n8459) );
  OR_GATE U9241 ( .I1(n8460), .I2(n8457), .O(n8458) );
  NAND_GATE U9242 ( .I1(n984), .I2(n8460), .O(n8464) );
  NAND3_GATE U9243 ( .I1(n8464), .I2(n8463), .I3(n8462), .O(n8465) );
  NAND_GATE U9244 ( .I1(B[13]), .I2(A[30]), .O(n8890) );
  INV_GATE U9245 ( .I1(n8890), .O(n8887) );
  NAND_GATE U9246 ( .I1(n799), .I2(n8887), .O(n8884) );
  OR_GATE U9247 ( .I1(n8466), .I2(n8471), .O(n8469) );
  OR_GATE U9248 ( .I1(n8470), .I2(n8467), .O(n8468) );
  NAND_GATE U9249 ( .I1(n975), .I2(n8470), .O(n8474) );
  NAND3_GATE U9250 ( .I1(n8474), .I2(n8473), .I3(n8472), .O(n8475) );
  NAND_GATE U9251 ( .I1(B[13]), .I2(A[29]), .O(n8901) );
  INV_GATE U9252 ( .I1(n8901), .O(n8898) );
  NAND_GATE U9253 ( .I1(n726), .I2(n8898), .O(n8895) );
  OR_GATE U9254 ( .I1(n8476), .I2(n8481), .O(n8479) );
  OR_GATE U9255 ( .I1(n8480), .I2(n8477), .O(n8478) );
  AND_GATE U9256 ( .I1(n8479), .I2(n8478), .O(n8486) );
  NAND_GATE U9257 ( .I1(n965), .I2(n8480), .O(n8484) );
  NAND3_GATE U9258 ( .I1(n8484), .I2(n8483), .I3(n8482), .O(n8485) );
  NAND_GATE U9259 ( .I1(n8486), .I2(n8485), .O(n9278) );
  NAND_GATE U9260 ( .I1(B[13]), .I2(A[28]), .O(n9284) );
  INV_GATE U9261 ( .I1(n9284), .O(n9279) );
  NAND_GATE U9262 ( .I1(n831), .I2(n9279), .O(n9277) );
  OR_GATE U9263 ( .I1(n8491), .I2(n8488), .O(n8489) );
  AND_GATE U9264 ( .I1(n8490), .I2(n8489), .O(n8497) );
  NAND_GATE U9265 ( .I1(n8492), .I2(n1336), .O(n8494) );
  NAND3_GATE U9266 ( .I1(n8495), .I2(n8494), .I3(n8493), .O(n8496) );
  NAND_GATE U9267 ( .I1(n8497), .I2(n8496), .O(n9264) );
  NAND_GATE U9268 ( .I1(B[13]), .I2(A[27]), .O(n9270) );
  INV_GATE U9269 ( .I1(n9270), .O(n9265) );
  NAND_GATE U9270 ( .I1(n901), .I2(n9265), .O(n9262) );
  OR_GATE U9271 ( .I1(n8498), .I2(n8503), .O(n8501) );
  OR_GATE U9272 ( .I1(n8502), .I2(n8499), .O(n8500) );
  AND_GATE U9273 ( .I1(n8501), .I2(n8500), .O(n8508) );
  NAND_GATE U9274 ( .I1(n594), .I2(n8502), .O(n8506) );
  NAND3_GATE U9275 ( .I1(n8506), .I2(n8505), .I3(n8504), .O(n8507) );
  NAND_GATE U9276 ( .I1(n8508), .I2(n8507), .O(n9253) );
  NAND_GATE U9277 ( .I1(B[13]), .I2(A[26]), .O(n9254) );
  INV_GATE U9278 ( .I1(n9254), .O(n9250) );
  NAND_GATE U9279 ( .I1(n807), .I2(n9250), .O(n9247) );
  OR_GATE U9280 ( .I1(n8509), .I2(n8514), .O(n8512) );
  OR_GATE U9281 ( .I1(n8513), .I2(n8510), .O(n8511) );
  NAND_GATE U9282 ( .I1(n954), .I2(n8513), .O(n8517) );
  NAND3_GATE U9283 ( .I1(n8517), .I2(n8516), .I3(n8515), .O(n8518) );
  NAND_GATE U9284 ( .I1(B[13]), .I2(A[25]), .O(n9240) );
  NAND_GATE U9285 ( .I1(n9237), .I2(n601), .O(n9233) );
  NAND_GATE U9286 ( .I1(B[13]), .I2(A[24]), .O(n9223) );
  INV_GATE U9287 ( .I1(n9223), .O(n9216) );
  OR_GATE U9288 ( .I1(n8523), .I2(n8520), .O(n8521) );
  AND_GATE U9289 ( .I1(n8522), .I2(n8521), .O(n8529) );
  NAND_GATE U9290 ( .I1(n957), .I2(n8523), .O(n8526) );
  NAND3_GATE U9291 ( .I1(n8527), .I2(n8526), .I3(n8525), .O(n8528) );
  NAND_GATE U9292 ( .I1(n8529), .I2(n8528), .O(n9219) );
  NAND_GATE U9293 ( .I1(n9216), .I2(n9217), .O(n9226) );
  NAND_GATE U9294 ( .I1(B[13]), .I2(A[23]), .O(n9375) );
  INV_GATE U9295 ( .I1(n9375), .O(n8907) );
  OR_GATE U9296 ( .I1(n8530), .I2(n8534), .O(n8533) );
  OR_GATE U9297 ( .I1(n8535), .I2(n8531), .O(n8532) );
  NAND_GATE U9298 ( .I1(n994), .I2(n8535), .O(n8536) );
  NAND3_GATE U9299 ( .I1(n8538), .I2(n8537), .I3(n8536), .O(n8539) );
  INV_GATE U9300 ( .I1(n8910), .O(n8909) );
  NAND_GATE U9301 ( .I1(n8907), .I2(n8909), .O(n8906) );
  NAND_GATE U9302 ( .I1(B[13]), .I2(A[22]), .O(n9384) );
  INV_GATE U9303 ( .I1(n9384), .O(n8920) );
  OR_GATE U9304 ( .I1(n8545), .I2(n8540), .O(n8543) );
  INV_GATE U9305 ( .I1(n8544), .O(n8546) );
  NAND3_GATE U9306 ( .I1(n8541), .I2(n8546), .I3(n8545), .O(n8542) );
  AND_GATE U9307 ( .I1(n8543), .I2(n8542), .O(n8551) );
  NAND_GATE U9308 ( .I1(n8544), .I2(n705), .O(n8548) );
  NAND_GATE U9309 ( .I1(n8546), .I2(n8545), .O(n8547) );
  NAND3_GATE U9310 ( .I1(n8549), .I2(n8548), .I3(n8547), .O(n8550) );
  NAND_GATE U9311 ( .I1(n8551), .I2(n8550), .O(n8916) );
  NAND_GATE U9312 ( .I1(n8920), .I2(n8918), .O(n8858) );
  NAND_GATE U9313 ( .I1(B[13]), .I2(A[21]), .O(n9410) );
  INV_GATE U9314 ( .I1(n9410), .O(n9203) );
  INV_GATE U9315 ( .I1(n8564), .O(n8560) );
  INV_GATE U9316 ( .I1(n8555), .O(n8556) );
  NAND_GATE U9317 ( .I1(n8557), .I2(n8556), .O(n8562) );
  NAND_GATE U9318 ( .I1(n8559), .I2(n8558), .O(n8561) );
  NAND3_GATE U9319 ( .I1(n8562), .I2(n8561), .I3(n8560), .O(n8567) );
  NAND_GATE U9320 ( .I1(n8562), .I2(n8561), .O(n8563) );
  NAND_GATE U9321 ( .I1(n8564), .I2(n8563), .O(n8566) );
  NAND3_GATE U9322 ( .I1(n8567), .I2(n8566), .I3(n8565), .O(n8853) );
  NAND3_GATE U9323 ( .I1(n8851), .I2(n8852), .I3(n8853), .O(n9205) );
  NAND_GATE U9324 ( .I1(n9203), .I2(n351), .O(n8855) );
  NAND_GATE U9325 ( .I1(B[13]), .I2(A[20]), .O(n9428) );
  NAND_GATE U9326 ( .I1(n8569), .I2(n8568), .O(n8576) );
  INV_GATE U9327 ( .I1(n8570), .O(n8572) );
  NAND_GATE U9328 ( .I1(n8572), .I2(n8571), .O(n8575) );
  NAND_GATE U9329 ( .I1(n8576), .I2(n8575), .O(n8573) );
  NAND_GATE U9330 ( .I1(n8581), .I2(n8573), .O(n8578) );
  INV_GATE U9331 ( .I1(n8581), .O(n8574) );
  NAND3_GATE U9332 ( .I1(n8576), .I2(n8575), .I3(n8574), .O(n8577) );
  NAND3_GATE U9333 ( .I1(n8579), .I2(n8578), .I3(n8577), .O(n8586) );
  OR_GATE U9334 ( .I1(n8581), .I2(n8580), .O(n8585) );
  OR_GATE U9335 ( .I1(n8583), .I2(n8582), .O(n8584) );
  NAND3_GATE U9336 ( .I1(n8586), .I2(n8585), .I3(n8584), .O(n8923) );
  NAND3_GATE U9337 ( .I1(n8587), .I2(n8589), .I3(n876), .O(n8844) );
  NAND3_GATE U9338 ( .I1(n8590), .I2(n1363), .I3(n8587), .O(n8843) );
  AND_GATE U9339 ( .I1(n8844), .I2(n8843), .O(n8592) );
  NAND_GATE U9340 ( .I1(n8590), .I2(n1363), .O(n8840) );
  NAND_GATE U9341 ( .I1(B[13]), .I2(A[19]), .O(n8935) );
  INV_GATE U9342 ( .I1(n8935), .O(n8847) );
  NAND3_GATE U9343 ( .I1(n8592), .I2(n8591), .I3(n8847), .O(n8927) );
  NAND_GATE U9344 ( .I1(B[13]), .I2(A[18]), .O(n9186) );
  INV_GATE U9345 ( .I1(n9186), .O(n9184) );
  NAND_GATE U9346 ( .I1(n8594), .I2(n8593), .O(n8597) );
  INV_GATE U9347 ( .I1(n8604), .O(n8596) );
  NAND_GATE U9348 ( .I1(n1362), .I2(n8595), .O(n8598) );
  NAND3_GATE U9349 ( .I1(n8597), .I2(n8596), .I3(n8598), .O(n8602) );
  NAND_GATE U9350 ( .I1(n8598), .I2(n8597), .O(n8599) );
  NAND_GATE U9351 ( .I1(n8604), .I2(n8599), .O(n8601) );
  NAND3_GATE U9352 ( .I1(n8602), .I2(n8601), .I3(n8600), .O(n8609) );
  OR_GATE U9353 ( .I1(n8604), .I2(n8603), .O(n8608) );
  OR_GATE U9354 ( .I1(n8606), .I2(n8605), .O(n8607) );
  NAND3_GATE U9355 ( .I1(n8609), .I2(n8608), .I3(n8607), .O(n9188) );
  INV_GATE U9356 ( .I1(n9188), .O(n9185) );
  NAND_GATE U9357 ( .I1(n9184), .I2(n9185), .O(n9192) );
  NAND_GATE U9358 ( .I1(B[13]), .I2(A[17]), .O(n8955) );
  INV_GATE U9359 ( .I1(n8955), .O(n8836) );
  NAND_GATE U9360 ( .I1(B[13]), .I2(A[16]), .O(n9166) );
  INV_GATE U9361 ( .I1(n9166), .O(n9169) );
  NAND_GATE U9362 ( .I1(n8610), .I2(n8618), .O(n8624) );
  INV_GATE U9363 ( .I1(n8624), .O(n8613) );
  INV_GATE U9364 ( .I1(n8611), .O(n8612) );
  NAND_GATE U9365 ( .I1(n8612), .I2(n8614), .O(n8626) );
  NAND_GATE U9366 ( .I1(n8613), .I2(n8626), .O(n8621) );
  NAND_GATE U9367 ( .I1(n8615), .I2(n8614), .O(n8619) );
  NAND_GATE U9368 ( .I1(n8617), .I2(n8616), .O(n8618) );
  NAND_GATE U9369 ( .I1(n8619), .I2(n8618), .O(n8622) );
  NAND_GATE U9370 ( .I1(n8623), .I2(n8622), .O(n8620) );
  NAND_GATE U9371 ( .I1(B[13]), .I2(A[15]), .O(n9161) );
  INV_GATE U9372 ( .I1(n9161), .O(n8812) );
  NAND3_GATE U9373 ( .I1(n8621), .I2(n8620), .I3(n8812), .O(n9153) );
  NAND_GATE U9374 ( .I1(n8624), .I2(n8620), .O(n8625) );
  NAND_GATE U9375 ( .I1(n8626), .I2(n8625), .O(n9158) );
  NAND_GATE U9376 ( .I1(B[13]), .I2(A[14]), .O(n8962) );
  INV_GATE U9377 ( .I1(n8962), .O(n8959) );
  NAND_GATE U9378 ( .I1(B[13]), .I2(A[13]), .O(n9143) );
  INV_GATE U9379 ( .I1(n9143), .O(n8781) );
  NAND_GATE U9380 ( .I1(B[13]), .I2(A[12]), .O(n8975) );
  INV_GATE U9381 ( .I1(n8975), .O(n8976) );
  NAND_GATE U9382 ( .I1(n8627), .I2(n8633), .O(n8629) );
  NAND_GATE U9383 ( .I1(n8631), .I2(n8630), .O(n8628) );
  NAND_GATE U9384 ( .I1(n8629), .I2(n8628), .O(n8756) );
  NAND_GATE U9385 ( .I1(n8757), .I2(n8756), .O(n9127) );
  INV_GATE U9386 ( .I1(n8769), .O(n8634) );
  NAND_GATE U9387 ( .I1(n8634), .I2(n8633), .O(n8761) );
  NAND_GATE U9388 ( .I1(n795), .I2(n8761), .O(n9126) );
  NAND_GATE U9389 ( .I1(B[13]), .I2(A[11]), .O(n9130) );
  INV_GATE U9390 ( .I1(n9130), .O(n8762) );
  NAND3_GATE U9391 ( .I1(n9127), .I2(n9126), .I3(n8762), .O(n9122) );
  NAND_GATE U9392 ( .I1(B[13]), .I2(A[10]), .O(n8986) );
  INV_GATE U9393 ( .I1(n8986), .O(n8989) );
  NAND_GATE U9394 ( .I1(B[13]), .I2(A[9]), .O(n9111) );
  INV_GATE U9395 ( .I1(n9111), .O(n8742) );
  OR_GATE U9396 ( .I1(n8636), .I2(n8635), .O(n8647) );
  NAND_GATE U9397 ( .I1(n8637), .I2(n8636), .O(n8641) );
  NAND_GATE U9398 ( .I1(n8638), .I2(n8641), .O(n8645) );
  NAND_GATE U9399 ( .I1(n8641), .I2(n8640), .O(n8642) );
  NAND_GATE U9400 ( .I1(n8643), .I2(n8642), .O(n8644) );
  NAND_GATE U9401 ( .I1(n8645), .I2(n8644), .O(n8646) );
  NAND_GATE U9402 ( .I1(n8647), .I2(n8646), .O(n9109) );
  NAND_GATE U9403 ( .I1(B[13]), .I2(A[8]), .O(n9005) );
  INV_GATE U9404 ( .I1(n9005), .O(n8999) );
  NAND_GATE U9405 ( .I1(B[13]), .I2(A[7]), .O(n9097) );
  INV_GATE U9406 ( .I1(n9097), .O(n8727) );
  OR_GATE U9407 ( .I1(n8649), .I2(n8648), .O(n8661) );
  NAND_GATE U9408 ( .I1(n8650), .I2(n8649), .O(n8655) );
  NAND_GATE U9409 ( .I1(n8651), .I2(n8655), .O(n8659) );
  NAND_GATE U9410 ( .I1(n8655), .I2(n8654), .O(n8656) );
  NAND_GATE U9411 ( .I1(n8657), .I2(n8656), .O(n8658) );
  NAND_GATE U9412 ( .I1(n8659), .I2(n8658), .O(n8660) );
  NAND_GATE U9413 ( .I1(n8661), .I2(n8660), .O(n9095) );
  NAND_GATE U9414 ( .I1(n8727), .I2(n9095), .O(n9092) );
  NAND_GATE U9415 ( .I1(B[13]), .I2(A[6]), .O(n9019) );
  INV_GATE U9416 ( .I1(n9019), .O(n9013) );
  NAND_GATE U9417 ( .I1(B[13]), .I2(A[5]), .O(n9083) );
  INV_GATE U9418 ( .I1(n9083), .O(n8713) );
  OR_GATE U9419 ( .I1(n8663), .I2(n8662), .O(n8675) );
  NAND_GATE U9420 ( .I1(n8664), .I2(n8663), .O(n8669) );
  NAND_GATE U9421 ( .I1(n8665), .I2(n8669), .O(n8673) );
  NAND_GATE U9422 ( .I1(n8667), .I2(n8666), .O(n8668) );
  NAND_GATE U9423 ( .I1(n8669), .I2(n8668), .O(n8670) );
  NAND_GATE U9424 ( .I1(n8671), .I2(n8670), .O(n8672) );
  NAND_GATE U9425 ( .I1(n8673), .I2(n8672), .O(n8674) );
  NAND_GATE U9426 ( .I1(n8675), .I2(n8674), .O(n9081) );
  NAND_GATE U9427 ( .I1(n8713), .I2(n9081), .O(n9078) );
  NAND_GATE U9428 ( .I1(B[13]), .I2(A[4]), .O(n9033) );
  INV_GATE U9429 ( .I1(n9033), .O(n9027) );
  NAND_GATE U9430 ( .I1(B[13]), .I2(A[3]), .O(n9068) );
  INV_GATE U9431 ( .I1(n9068), .O(n8698) );
  INV_GATE U9432 ( .I1(n8676), .O(n8677) );
  NAND_GATE U9433 ( .I1(n8677), .I2(n8680), .O(n8689) );
  NAND_GATE U9434 ( .I1(n8679), .I2(n8683), .O(n8687) );
  NAND_GATE U9435 ( .I1(n8681), .I2(n8680), .O(n8682) );
  NAND_GATE U9436 ( .I1(n8683), .I2(n8682), .O(n8684) );
  NAND_GATE U9437 ( .I1(n8685), .I2(n8684), .O(n8686) );
  NAND_GATE U9438 ( .I1(n8687), .I2(n8686), .O(n8688) );
  NAND_GATE U9439 ( .I1(n8689), .I2(n8688), .O(n9066) );
  NAND_GATE U9440 ( .I1(n8698), .I2(n9066), .O(n9063) );
  NAND_GATE U9441 ( .I1(B[13]), .I2(A[2]), .O(n9047) );
  INV_GATE U9442 ( .I1(n9047), .O(n9041) );
  NAND3_GATE U9443 ( .I1(B[13]), .I2(n1425), .I3(n1254), .O(n9040) );
  INV_GATE U9444 ( .I1(n9040), .O(n9043) );
  NAND_GATE U9445 ( .I1(n9041), .I2(n9043), .O(n9038) );
  NAND_GATE U9446 ( .I1(n1426), .I2(A[0]), .O(n8690) );
  NAND_GATE U9447 ( .I1(n14241), .I2(n8690), .O(n8691) );
  NAND_GATE U9448 ( .I1(B[15]), .I2(n8691), .O(n8695) );
  NAND_GATE U9449 ( .I1(n1427), .I2(A[1]), .O(n8692) );
  NAND_GATE U9450 ( .I1(n724), .I2(n8692), .O(n8693) );
  NAND_GATE U9451 ( .I1(n1425), .I2(n8693), .O(n8694) );
  NAND_GATE U9452 ( .I1(n8695), .I2(n8694), .O(n9042) );
  NAND_GATE U9453 ( .I1(n9047), .I2(n9040), .O(n8696) );
  NAND_GATE U9454 ( .I1(n9042), .I2(n8696), .O(n8697) );
  NAND_GATE U9455 ( .I1(n9038), .I2(n8697), .O(n9067) );
  NAND_GATE U9456 ( .I1(n9066), .I2(n9067), .O(n8699) );
  NAND_GATE U9457 ( .I1(n8698), .I2(n9067), .O(n9062) );
  NAND3_GATE U9458 ( .I1(n9063), .I2(n8699), .I3(n9062), .O(n9029) );
  NAND_GATE U9459 ( .I1(n9027), .I2(n9029), .O(n9024) );
  OR_GATE U9460 ( .I1(n8700), .I2(n8704), .O(n8703) );
  OR_GATE U9461 ( .I1(n8705), .I2(n8701), .O(n8702) );
  AND_GATE U9462 ( .I1(n8703), .I2(n8702), .O(n8710) );
  NAND_GATE U9463 ( .I1(n8704), .I2(n1238), .O(n8708) );
  NAND3_GATE U9464 ( .I1(n8708), .I2(n8707), .I3(n8706), .O(n8709) );
  NAND_GATE U9465 ( .I1(n8710), .I2(n8709), .O(n9025) );
  INV_GATE U9466 ( .I1(n9025), .O(n9028) );
  INV_GATE U9467 ( .I1(n9029), .O(n9026) );
  NAND_GATE U9468 ( .I1(n9033), .I2(n9026), .O(n8711) );
  NAND_GATE U9469 ( .I1(n9028), .I2(n8711), .O(n8712) );
  NAND_GATE U9470 ( .I1(n9024), .I2(n8712), .O(n9082) );
  NAND_GATE U9471 ( .I1(n9081), .I2(n9082), .O(n8714) );
  NAND_GATE U9472 ( .I1(n8713), .I2(n9082), .O(n9077) );
  NAND3_GATE U9473 ( .I1(n9078), .I2(n8714), .I3(n9077), .O(n9015) );
  NAND_GATE U9474 ( .I1(n9013), .I2(n9015), .O(n9010) );
  OR_GATE U9475 ( .I1(n8715), .I2(n8719), .O(n8718) );
  OR_GATE U9476 ( .I1(n8720), .I2(n8716), .O(n8717) );
  NAND_GATE U9477 ( .I1(n8719), .I2(n1155), .O(n8723) );
  NAND3_GATE U9478 ( .I1(n8723), .I2(n8722), .I3(n8721), .O(n8724) );
  INV_GATE U9479 ( .I1(n9011), .O(n9014) );
  INV_GATE U9480 ( .I1(n9015), .O(n9012) );
  NAND_GATE U9481 ( .I1(n9019), .I2(n9012), .O(n8725) );
  NAND_GATE U9482 ( .I1(n9014), .I2(n8725), .O(n8726) );
  NAND_GATE U9483 ( .I1(n9010), .I2(n8726), .O(n9096) );
  NAND_GATE U9484 ( .I1(n9095), .I2(n9096), .O(n8728) );
  NAND_GATE U9485 ( .I1(n8727), .I2(n9096), .O(n9091) );
  NAND3_GATE U9486 ( .I1(n9092), .I2(n8728), .I3(n9091), .O(n9001) );
  NAND_GATE U9487 ( .I1(n8999), .I2(n9001), .O(n8996) );
  OR_GATE U9488 ( .I1(n8729), .I2(n8733), .O(n8732) );
  OR_GATE U9489 ( .I1(n8734), .I2(n8730), .O(n8731) );
  AND_GATE U9490 ( .I1(n8732), .I2(n8731), .O(n8739) );
  NAND_GATE U9491 ( .I1(n8733), .I2(n1012), .O(n8737) );
  NAND3_GATE U9492 ( .I1(n8737), .I2(n8736), .I3(n8735), .O(n8738) );
  NAND_GATE U9493 ( .I1(n8739), .I2(n8738), .O(n8997) );
  INV_GATE U9494 ( .I1(n8997), .O(n9000) );
  INV_GATE U9495 ( .I1(n9001), .O(n8998) );
  NAND_GATE U9496 ( .I1(n9005), .I2(n8998), .O(n8740) );
  NAND_GATE U9497 ( .I1(n9000), .I2(n8740), .O(n8741) );
  NAND_GATE U9498 ( .I1(n8996), .I2(n8741), .O(n9110) );
  NAND_GATE U9499 ( .I1(n9109), .I2(n9110), .O(n8743) );
  NAND_GATE U9500 ( .I1(n8742), .I2(n9110), .O(n9105) );
  NAND3_GATE U9501 ( .I1(n9106), .I2(n8743), .I3(n9105), .O(n8982) );
  NAND_GATE U9502 ( .I1(n8989), .I2(n8982), .O(n8992) );
  OR_GATE U9503 ( .I1(n8744), .I2(n8745), .O(n8753) );
  NAND_GATE U9504 ( .I1(n8745), .I2(n1317), .O(n8746) );
  NAND3_GATE U9505 ( .I1(n8748), .I2(n8747), .I3(n8746), .O(n8752) );
  OR_GATE U9506 ( .I1(n8750), .I2(n8749), .O(n8751) );
  INV_GATE U9507 ( .I1(n8982), .O(n8987) );
  NAND_GATE U9508 ( .I1(n8986), .I2(n8987), .O(n8754) );
  NAND_GATE U9509 ( .I1(n802), .I2(n8754), .O(n8755) );
  NAND_GATE U9510 ( .I1(n8992), .I2(n8755), .O(n9129) );
  NAND_GATE U9511 ( .I1(n8759), .I2(n8758), .O(n8760) );
  NAND_GATE U9512 ( .I1(n8761), .I2(n8760), .O(n9120) );
  NAND_GATE U9513 ( .I1(n9129), .I2(n9120), .O(n8763) );
  NAND_GATE U9514 ( .I1(n8762), .I2(n9129), .O(n9121) );
  NAND3_GATE U9515 ( .I1(n9122), .I2(n8763), .I3(n9121), .O(n8971) );
  NAND_GATE U9516 ( .I1(n8976), .I2(n8971), .O(n8979) );
  OR_GATE U9517 ( .I1(n8765), .I2(n8764), .O(n8778) );
  NAND_GATE U9518 ( .I1(n8768), .I2(n8767), .O(n8766) );
  NAND_GATE U9519 ( .I1(n8775), .I2(n8766), .O(n8772) );
  NAND4_GATE U9520 ( .I1(n8770), .I2(n8769), .I3(n8768), .I4(n8767), .O(n8771)
         );
  NAND3_GATE U9521 ( .I1(n8773), .I2(n8772), .I3(n8771), .O(n8777) );
  OR_GATE U9522 ( .I1(n8775), .I2(n8774), .O(n8776) );
  NAND3_GATE U9523 ( .I1(n8778), .I2(n8777), .I3(n8776), .O(n8980) );
  INV_GATE U9524 ( .I1(n8980), .O(n8970) );
  NAND_GATE U9525 ( .I1(n8975), .I2(n690), .O(n8779) );
  NAND_GATE U9526 ( .I1(n8970), .I2(n8779), .O(n8780) );
  NAND_GATE U9527 ( .I1(n8979), .I2(n8780), .O(n9144) );
  NAND_GATE U9528 ( .I1(n8781), .I2(n9144), .O(n9139) );
  NAND_GATE U9529 ( .I1(n8782), .I2(n8786), .O(n8790) );
  NAND_GATE U9530 ( .I1(n8783), .I2(n8792), .O(n8786) );
  NAND_GATE U9531 ( .I1(n8784), .I2(n1297), .O(n8785) );
  NAND_GATE U9532 ( .I1(n8786), .I2(n8785), .O(n8787) );
  NAND_GATE U9533 ( .I1(n8788), .I2(n8787), .O(n8789) );
  NAND_GATE U9534 ( .I1(n8790), .I2(n8789), .O(n8794) );
  OR_GATE U9535 ( .I1(n8792), .I2(n8791), .O(n8793) );
  NAND_GATE U9536 ( .I1(n8794), .I2(n8793), .O(n9140) );
  NAND_GATE U9537 ( .I1(n9144), .I2(n9140), .O(n8795) );
  NAND3_GATE U9538 ( .I1(A[13]), .I2(n9140), .I3(B[13]), .O(n9145) );
  NAND_GATE U9539 ( .I1(n8959), .I2(n8961), .O(n8966) );
  NAND_GATE U9540 ( .I1(n8797), .I2(n8798), .O(n8796) );
  NAND_GATE U9541 ( .I1(n8804), .I2(n8796), .O(n8801) );
  INV_GATE U9542 ( .I1(n8804), .O(n8799) );
  NAND3_GATE U9543 ( .I1(n8799), .I2(n8798), .I3(n8797), .O(n8800) );
  NAND3_GATE U9544 ( .I1(n8802), .I2(n8801), .I3(n8800), .O(n8809) );
  OR_GATE U9545 ( .I1(n8804), .I2(n8803), .O(n8808) );
  OR_GATE U9546 ( .I1(n8806), .I2(n8805), .O(n8807) );
  NAND3_GATE U9547 ( .I1(n8809), .I2(n8808), .I3(n8807), .O(n8967) );
  INV_GATE U9548 ( .I1(n8967), .O(n8960) );
  NAND_GATE U9549 ( .I1(n8962), .I2(n762), .O(n8810) );
  NAND_GATE U9550 ( .I1(n8960), .I2(n8810), .O(n8811) );
  NAND_GATE U9551 ( .I1(n8966), .I2(n8811), .O(n9157) );
  NAND_GATE U9552 ( .I1(n9158), .I2(n9157), .O(n8813) );
  NAND_GATE U9553 ( .I1(n8812), .I2(n9157), .O(n9154) );
  NAND3_GATE U9554 ( .I1(n9153), .I2(n8813), .I3(n9154), .O(n9171) );
  NAND_GATE U9555 ( .I1(n9169), .I2(n9171), .O(n9175) );
  OR_GATE U9556 ( .I1(n8814), .I2(n8821), .O(n8817) );
  INV_GATE U9557 ( .I1(n8820), .O(n8822) );
  NAND3_GATE U9558 ( .I1(n8822), .I2(n8815), .I3(n8821), .O(n8816) );
  AND_GATE U9559 ( .I1(n8817), .I2(n8816), .O(n8827) );
  NAND3_GATE U9560 ( .I1(n8820), .I2(n8819), .I3(n8818), .O(n8824) );
  NAND_GATE U9561 ( .I1(n8822), .I2(n8821), .O(n8823) );
  NAND3_GATE U9562 ( .I1(n8825), .I2(n8824), .I3(n8823), .O(n8826) );
  NAND_GATE U9563 ( .I1(n8827), .I2(n8826), .O(n9176) );
  INV_GATE U9564 ( .I1(n9176), .O(n9170) );
  NAND_GATE U9565 ( .I1(n9166), .I2(n9167), .O(n8828) );
  NAND_GATE U9566 ( .I1(n9170), .I2(n8828), .O(n8829) );
  NAND_GATE U9567 ( .I1(n9175), .I2(n8829), .O(n8950) );
  NAND_GATE U9568 ( .I1(n8836), .I2(n8950), .O(n8944) );
  NAND_GATE U9569 ( .I1(n395), .I2(n292), .O(n8831) );
  NAND_GATE U9570 ( .I1(n1386), .I2(n8832), .O(n8830) );
  NAND_GATE U9571 ( .I1(n8831), .I2(n8830), .O(n8939) );
  NAND_GATE U9572 ( .I1(n8940), .I2(n8939), .O(n8947) );
  NAND_GATE U9573 ( .I1(n8833), .I2(n8830), .O(n8941) );
  INV_GATE U9574 ( .I1(n8941), .O(n8835) );
  NAND_GATE U9575 ( .I1(n8835), .I2(n8943), .O(n8948) );
  NAND3_GATE U9576 ( .I1(n8947), .I2(n8948), .I3(n8950), .O(n8837) );
  NAND3_GATE U9577 ( .I1(n8947), .I2(n8948), .I3(n8836), .O(n8938) );
  NAND3_GATE U9578 ( .I1(n8944), .I2(n8837), .I3(n8938), .O(n9193) );
  NAND_GATE U9579 ( .I1(n9186), .I2(n9188), .O(n8838) );
  NAND_GATE U9580 ( .I1(n9193), .I2(n8838), .O(n8839) );
  NAND_GATE U9581 ( .I1(n9192), .I2(n8839), .O(n8932) );
  NAND_GATE U9582 ( .I1(n8841), .I2(n8840), .O(n8842) );
  NAND3_GATE U9583 ( .I1(n8844), .I2(n8843), .I3(n8842), .O(n8845) );
  NAND_GATE U9584 ( .I1(n8846), .I2(n8845), .O(n8931) );
  NAND_GATE U9585 ( .I1(n8932), .I2(n8931), .O(n8848) );
  NAND_GATE U9586 ( .I1(n8847), .I2(n8932), .O(n8928) );
  NAND3_GATE U9587 ( .I1(n8927), .I2(n8848), .I3(n8928), .O(n8924) );
  NAND_GATE U9588 ( .I1(n9428), .I2(n8923), .O(n8849) );
  NAND_GATE U9589 ( .I1(n8924), .I2(n8849), .O(n8850) );
  NAND_GATE U9590 ( .I1(n8922), .I2(n8850), .O(n9207) );
  NAND4_GATE U9591 ( .I1(n8853), .I2(n8852), .I3(n8851), .I4(n9207), .O(n8854)
         );
  NAND_GATE U9592 ( .I1(n9203), .I2(n9207), .O(n9204) );
  NAND_GATE U9593 ( .I1(n9384), .I2(n8916), .O(n8856) );
  NAND_GATE U9594 ( .I1(n8919), .I2(n8856), .O(n8857) );
  NAND_GATE U9595 ( .I1(n8858), .I2(n8857), .O(n8908) );
  NAND_GATE U9596 ( .I1(n9375), .I2(n8910), .O(n8859) );
  NAND_GATE U9597 ( .I1(n8908), .I2(n8859), .O(n8860) );
  NAND_GATE U9598 ( .I1(n8906), .I2(n8860), .O(n9227) );
  NAND_GATE U9599 ( .I1(n9223), .I2(n9219), .O(n8861) );
  NAND_GATE U9600 ( .I1(n9227), .I2(n8861), .O(n8862) );
  NAND_GATE U9601 ( .I1(n9226), .I2(n8862), .O(n9236) );
  NAND_GATE U9602 ( .I1(n9239), .I2(n9240), .O(n8863) );
  NAND_GATE U9603 ( .I1(n9236), .I2(n8863), .O(n8864) );
  NAND_GATE U9604 ( .I1(n9233), .I2(n8864), .O(n9251) );
  NAND_GATE U9605 ( .I1(n9253), .I2(n9254), .O(n8865) );
  NAND_GATE U9606 ( .I1(n9251), .I2(n8865), .O(n8866) );
  NAND_GATE U9607 ( .I1(n9247), .I2(n8866), .O(n9266) );
  NAND_GATE U9608 ( .I1(n9264), .I2(n9270), .O(n8867) );
  NAND_GATE U9609 ( .I1(n9266), .I2(n8867), .O(n8868) );
  NAND_GATE U9610 ( .I1(n9278), .I2(n9284), .O(n8869) );
  NAND_GATE U9611 ( .I1(n9280), .I2(n8869), .O(n8870) );
  NAND_GATE U9612 ( .I1(n9277), .I2(n8870), .O(n8899) );
  NAND_GATE U9613 ( .I1(n8897), .I2(n8901), .O(n8871) );
  NAND_GATE U9614 ( .I1(n8899), .I2(n8871), .O(n8872) );
  NAND_GATE U9615 ( .I1(n8895), .I2(n8872), .O(n8888) );
  NAND_GATE U9616 ( .I1(n8886), .I2(n8890), .O(n8873) );
  NAND_GATE U9617 ( .I1(n8888), .I2(n8873), .O(n8875) );
  NAND_GATE U9618 ( .I1(n1424), .I2(A[31]), .O(n8874) );
  NAND3_GATE U9619 ( .I1(n8884), .I2(n8875), .I3(n8874), .O(n8879) );
  INV_GATE U9620 ( .I1(n8883), .O(n14813) );
  NAND_GATE U9621 ( .I1(n8876), .I2(n14813), .O(n8877) );
  NAND_GATE U9622 ( .I1(n8878), .I2(n8877), .O(\A1[43] ) );
  INV_GATE U9623 ( .I1(n8879), .O(n8880) );
  NAND_GATE U9624 ( .I1(n8881), .I2(n8880), .O(n8882) );
  NAND_GATE U9625 ( .I1(n8883), .I2(n8882), .O(n9293) );
  INV_GATE U9626 ( .I1(n9293), .O(n14815) );
  INV_GATE U9627 ( .I1(n8884), .O(n8885) );
  NAND_GATE U9628 ( .I1(n8885), .I2(n8888), .O(n8894) );
  NAND_GATE U9629 ( .I1(n8887), .I2(n8889), .O(n8892) );
  NAND_GATE U9630 ( .I1(n8892), .I2(n8891), .O(n8893) );
  NAND_GATE U9631 ( .I1(n8894), .I2(n8893), .O(n9296) );
  NAND_GATE U9632 ( .I1(n1422), .I2(A[30]), .O(n9307) );
  INV_GATE U9633 ( .I1(n9307), .O(n9290) );
  INV_GATE U9634 ( .I1(n8895), .O(n8896) );
  NAND_GATE U9635 ( .I1(n8896), .I2(n8899), .O(n8905) );
  NAND_GATE U9636 ( .I1(n8898), .I2(n8900), .O(n8903) );
  NAND_GATE U9637 ( .I1(n8903), .I2(n8902), .O(n8904) );
  NAND_GATE U9638 ( .I1(n8905), .I2(n8904), .O(n9305) );
  NAND_GATE U9639 ( .I1(n1422), .I2(A[29]), .O(n9319) );
  INV_GATE U9640 ( .I1(n9319), .O(n9288) );
  NAND_GATE U9641 ( .I1(n1422), .I2(A[28]), .O(n9324) );
  INV_GATE U9642 ( .I1(n9324), .O(n9275) );
  NAND_GATE U9643 ( .I1(n1422), .I2(A[27]), .O(n9342) );
  INV_GATE U9644 ( .I1(n9342), .O(n9334) );
  NAND_GATE U9645 ( .I1(n1422), .I2(A[26]), .O(n9345) );
  INV_GATE U9646 ( .I1(n9345), .O(n9245) );
  NAND_GATE U9647 ( .I1(n1422), .I2(A[25]), .O(n9363) );
  INV_GATE U9648 ( .I1(n9363), .O(n9231) );
  NAND_GATE U9649 ( .I1(n1422), .I2(A[24]), .O(n9379) );
  INV_GATE U9650 ( .I1(n9379), .O(n9214) );
  NAND_GATE U9651 ( .I1(n8907), .I2(n8911), .O(n9371) );
  NAND_GATE U9652 ( .I1(n8909), .I2(n8908), .O(n8912) );
  NAND_GATE U9653 ( .I1(n8910), .I2(n1018), .O(n8911) );
  NAND_GATE U9654 ( .I1(n8912), .I2(n8911), .O(n9374) );
  NAND_GATE U9655 ( .I1(n9375), .I2(n9374), .O(n8913) );
  NAND_GATE U9656 ( .I1(n9371), .I2(n8913), .O(n8914) );
  NAND_GATE U9657 ( .I1(n9373), .I2(n8914), .O(n9366) );
  NAND_GATE U9658 ( .I1(n9214), .I2(n9366), .O(n9368) );
  NAND_GATE U9659 ( .I1(n1422), .I2(A[23]), .O(n9393) );
  INV_GATE U9660 ( .I1(n9393), .O(n9212) );
  NAND_GATE U9661 ( .I1(n8918), .I2(n8919), .O(n8915) );
  NAND_GATE U9662 ( .I1(n8915), .I2(n8917), .O(n9383) );
  NAND_GATE U9663 ( .I1(n8916), .I2(n352), .O(n8917) );
  NAND_GATE U9664 ( .I1(n8920), .I2(n8917), .O(n9385) );
  NAND_GATE U9665 ( .I1(n9388), .I2(n9385), .O(n8921) );
  NAND3_GATE U9666 ( .I1(n8920), .I2(n8919), .I3(n8918), .O(n9386) );
  NAND_GATE U9667 ( .I1(n8921), .I2(n9386), .O(n9396) );
  NAND_GATE U9668 ( .I1(n9212), .I2(n9396), .O(n9394) );
  NAND_GATE U9669 ( .I1(n1422), .I2(A[22]), .O(n9416) );
  INV_GATE U9670 ( .I1(n9416), .O(n9210) );
  NAND_GATE U9671 ( .I1(n1422), .I2(A[21]), .O(n9433) );
  INV_GATE U9672 ( .I1(n9433), .O(n9200) );
  NAND_GATE U9673 ( .I1(n1276), .I2(n9423), .O(n9430) );
  NAND_GATE U9674 ( .I1(n8923), .I2(n1017), .O(n8926) );
  NAND_GATE U9675 ( .I1(n8926), .I2(n8925), .O(n9427) );
  NAND_GATE U9676 ( .I1(n9428), .I2(n9427), .O(n9201) );
  NAND3_GATE U9677 ( .I1(n9200), .I2(n9430), .I3(n9201), .O(n9426) );
  NAND_GATE U9678 ( .I1(n1422), .I2(A[20]), .O(n9757) );
  INV_GATE U9679 ( .I1(n9757), .O(n9684) );
  OR_GATE U9680 ( .I1(n8932), .I2(n8927), .O(n8930) );
  OR_GATE U9681 ( .I1(n8928), .I2(n8931), .O(n8929) );
  AND_GATE U9682 ( .I1(n8930), .I2(n8929), .O(n8937) );
  NAND_GATE U9683 ( .I1(n1024), .I2(n8931), .O(n8934) );
  NAND3_GATE U9684 ( .I1(n8935), .I2(n8934), .I3(n8933), .O(n8936) );
  NAND_GATE U9685 ( .I1(n8937), .I2(n8936), .O(n9687) );
  NAND_GATE U9686 ( .I1(n9684), .I2(n875), .O(n9683) );
  NAND_GATE U9687 ( .I1(n1422), .I2(A[19]), .O(n9441) );
  INV_GATE U9688 ( .I1(n9441), .O(n9196) );
  NAND_GATE U9689 ( .I1(n1422), .I2(A[18]), .O(n9776) );
  INV_GATE U9690 ( .I1(n9776), .O(n9671) );
  OR_GATE U9691 ( .I1(n8938), .I2(n8950), .O(n8946) );
  NAND_GATE U9692 ( .I1(n8941), .I2(n8947), .O(n8942) );
  NAND_GATE U9693 ( .I1(n8943), .I2(n8942), .O(n8951) );
  OR_GATE U9694 ( .I1(n8951), .I2(n8944), .O(n8945) );
  AND_GATE U9695 ( .I1(n8946), .I2(n8945), .O(n8957) );
  NAND_GATE U9696 ( .I1(n8948), .I2(n8947), .O(n8949) );
  NAND_GATE U9697 ( .I1(n8950), .I2(n8949), .O(n8954) );
  INV_GATE U9698 ( .I1(n8950), .O(n8952) );
  NAND_GATE U9699 ( .I1(n8952), .I2(n8951), .O(n8953) );
  NAND3_GATE U9700 ( .I1(n8955), .I2(n8954), .I3(n8953), .O(n8956) );
  NAND_GATE U9701 ( .I1(n8957), .I2(n8956), .O(n9675) );
  NAND_GATE U9702 ( .I1(n9671), .I2(n394), .O(n9672) );
  NAND_GATE U9703 ( .I1(n1422), .I2(A[17]), .O(n9457) );
  INV_GATE U9704 ( .I1(n9457), .O(n9179) );
  NAND_GATE U9705 ( .I1(n1422), .I2(A[16]), .O(n9797) );
  INV_GATE U9706 ( .I1(n9797), .O(n9664) );
  NAND_GATE U9707 ( .I1(n762), .I2(n8967), .O(n8958) );
  NAND_GATE U9708 ( .I1(n8959), .I2(n8958), .O(n8965) );
  NAND_GATE U9709 ( .I1(n8961), .I2(n8960), .O(n8964) );
  NAND3_GATE U9710 ( .I1(n762), .I2(n8962), .I3(n8967), .O(n8963) );
  NAND3_GATE U9711 ( .I1(n8965), .I2(n8964), .I3(n8963), .O(n8969) );
  OR_GATE U9712 ( .I1(n8967), .I2(n8966), .O(n8968) );
  NAND_GATE U9713 ( .I1(n8969), .I2(n8968), .O(n9646) );
  NAND3_GATE U9714 ( .I1(A[15]), .I2(n9646), .I3(n1422), .O(n9650) );
  NAND_GATE U9715 ( .I1(n1422), .I2(A[14]), .O(n9469) );
  INV_GATE U9716 ( .I1(n9469), .O(n9463) );
  NAND_GATE U9717 ( .I1(n1422), .I2(A[13]), .O(n9633) );
  INV_GATE U9718 ( .I1(n9633), .O(n9137) );
  NAND_GATE U9719 ( .I1(n8971), .I2(n8970), .O(n8973) );
  NAND_GATE U9720 ( .I1(n690), .I2(n8980), .O(n8972) );
  NAND_GATE U9721 ( .I1(n8973), .I2(n8972), .O(n8974) );
  NAND_GATE U9722 ( .I1(n8975), .I2(n8974), .O(n8978) );
  NAND_GATE U9723 ( .I1(n8976), .I2(n8972), .O(n8977) );
  OR_GATE U9724 ( .I1(n8980), .I2(n8979), .O(n8981) );
  NAND_GATE U9725 ( .I1(n1422), .I2(A[12]), .O(n9989) );
  INV_GATE U9726 ( .I1(n9989), .O(n9478) );
  NAND_GATE U9727 ( .I1(n8982), .I2(n802), .O(n8984) );
  NAND_GATE U9728 ( .I1(n8984), .I2(n8983), .O(n8985) );
  NAND_GATE U9729 ( .I1(n8986), .I2(n8985), .O(n8991) );
  NAND_GATE U9730 ( .I1(n8987), .I2(n8993), .O(n8988) );
  NAND_GATE U9731 ( .I1(n8989), .I2(n8988), .O(n8990) );
  NAND_GATE U9732 ( .I1(n8991), .I2(n8990), .O(n8995) );
  OR_GATE U9733 ( .I1(n8993), .I2(n8992), .O(n8994) );
  NAND_GATE U9734 ( .I1(n8995), .I2(n8994), .O(n9618) );
  NAND3_GATE U9735 ( .I1(A[11]), .I2(n9618), .I3(n1422), .O(n9622) );
  NAND_GATE U9736 ( .I1(n1422), .I2(A[10]), .O(n9488) );
  INV_GATE U9737 ( .I1(n9488), .O(n9482) );
  NAND_GATE U9738 ( .I1(n1422), .I2(A[9]), .O(n9609) );
  INV_GATE U9739 ( .I1(n9609), .O(n9103) );
  OR_GATE U9740 ( .I1(n8997), .I2(n8996), .O(n9009) );
  NAND_GATE U9741 ( .I1(n8998), .I2(n8997), .O(n9003) );
  NAND_GATE U9742 ( .I1(n8999), .I2(n9003), .O(n9007) );
  NAND_GATE U9743 ( .I1(n9001), .I2(n9000), .O(n9002) );
  NAND_GATE U9744 ( .I1(n9003), .I2(n9002), .O(n9004) );
  NAND_GATE U9745 ( .I1(n9005), .I2(n9004), .O(n9006) );
  NAND_GATE U9746 ( .I1(n9007), .I2(n9006), .O(n9008) );
  NAND_GATE U9747 ( .I1(n9009), .I2(n9008), .O(n9607) );
  NAND_GATE U9748 ( .I1(n9103), .I2(n9607), .O(n9603) );
  NAND_GATE U9749 ( .I1(n1422), .I2(A[8]), .O(n9502) );
  INV_GATE U9750 ( .I1(n9502), .O(n9496) );
  NAND_GATE U9751 ( .I1(n1422), .I2(A[7]), .O(n9594) );
  INV_GATE U9752 ( .I1(n9594), .O(n9089) );
  OR_GATE U9753 ( .I1(n9011), .I2(n9010), .O(n9023) );
  NAND_GATE U9754 ( .I1(n9012), .I2(n9011), .O(n9017) );
  NAND_GATE U9755 ( .I1(n9013), .I2(n9017), .O(n9021) );
  NAND_GATE U9756 ( .I1(n9015), .I2(n9014), .O(n9016) );
  NAND_GATE U9757 ( .I1(n9017), .I2(n9016), .O(n9018) );
  NAND_GATE U9758 ( .I1(n9019), .I2(n9018), .O(n9020) );
  NAND_GATE U9759 ( .I1(n9021), .I2(n9020), .O(n9022) );
  NAND_GATE U9760 ( .I1(n9023), .I2(n9022), .O(n9592) );
  NAND_GATE U9761 ( .I1(n9089), .I2(n9592), .O(n9589) );
  NAND_GATE U9762 ( .I1(n1422), .I2(A[6]), .O(n9516) );
  INV_GATE U9763 ( .I1(n9516), .O(n9510) );
  NAND_GATE U9764 ( .I1(n1422), .I2(A[5]), .O(n9580) );
  INV_GATE U9765 ( .I1(n9580), .O(n9075) );
  OR_GATE U9766 ( .I1(n9025), .I2(n9024), .O(n9037) );
  NAND_GATE U9767 ( .I1(n9026), .I2(n9025), .O(n9031) );
  NAND_GATE U9768 ( .I1(n9027), .I2(n9031), .O(n9035) );
  NAND_GATE U9769 ( .I1(n9029), .I2(n9028), .O(n9030) );
  NAND_GATE U9770 ( .I1(n9031), .I2(n9030), .O(n9032) );
  NAND_GATE U9771 ( .I1(n9033), .I2(n9032), .O(n9034) );
  NAND_GATE U9772 ( .I1(n9035), .I2(n9034), .O(n9036) );
  NAND_GATE U9773 ( .I1(n9037), .I2(n9036), .O(n9578) );
  NAND_GATE U9774 ( .I1(n9075), .I2(n9578), .O(n9575) );
  NAND_GATE U9775 ( .I1(n1422), .I2(A[4]), .O(n9530) );
  INV_GATE U9776 ( .I1(n9530), .O(n9524) );
  INV_GATE U9777 ( .I1(n9038), .O(n9039) );
  NAND_GATE U9778 ( .I1(n9039), .I2(n9042), .O(n9051) );
  NAND_GATE U9779 ( .I1(n9041), .I2(n9045), .O(n9049) );
  NAND_GATE U9780 ( .I1(n9043), .I2(n9042), .O(n9044) );
  NAND_GATE U9781 ( .I1(n9045), .I2(n9044), .O(n9046) );
  NAND_GATE U9782 ( .I1(n9047), .I2(n9046), .O(n9048) );
  NAND_GATE U9783 ( .I1(n9049), .I2(n9048), .O(n9050) );
  NAND_GATE U9784 ( .I1(n9051), .I2(n9050), .O(n9539) );
  NAND_GATE U9785 ( .I1(n1424), .I2(A[0]), .O(n9052) );
  NAND_GATE U9786 ( .I1(n14241), .I2(n9052), .O(n9053) );
  NAND_GATE U9787 ( .I1(n1425), .I2(n9053), .O(n9057) );
  NAND_GATE U9788 ( .I1(n1426), .I2(A[1]), .O(n9054) );
  NAND_GATE U9789 ( .I1(n724), .I2(n9054), .O(n9055) );
  NAND_GATE U9790 ( .I1(B[13]), .I2(n9055), .O(n9056) );
  NAND_GATE U9791 ( .I1(n9057), .I2(n9056), .O(n9551) );
  NAND_GATE U9792 ( .I1(n1422), .I2(A[2]), .O(n9555) );
  NAND3_GATE U9793 ( .I1(n1422), .I2(B[13]), .I3(n1254), .O(n9548) );
  NAND_GATE U9794 ( .I1(n9555), .I2(n9548), .O(n9058) );
  NAND_GATE U9795 ( .I1(n9551), .I2(n9058), .O(n9059) );
  INV_GATE U9796 ( .I1(n9555), .O(n9549) );
  INV_GATE U9797 ( .I1(n9548), .O(n9550) );
  NAND_GATE U9798 ( .I1(n9549), .I2(n9550), .O(n9546) );
  NAND_GATE U9799 ( .I1(n9059), .I2(n9546), .O(n9540) );
  NAND_GATE U9800 ( .I1(n9539), .I2(n9540), .O(n9061) );
  NAND_GATE U9801 ( .I1(n1422), .I2(A[3]), .O(n9541) );
  INV_GATE U9802 ( .I1(n9541), .O(n9060) );
  NAND_GATE U9803 ( .I1(n9539), .I2(n9060), .O(n9536) );
  NAND_GATE U9804 ( .I1(n9540), .I2(n9060), .O(n9535) );
  NAND3_GATE U9805 ( .I1(n9061), .I2(n9536), .I3(n9535), .O(n9526) );
  NAND_GATE U9806 ( .I1(n9524), .I2(n9526), .O(n9521) );
  OR_GATE U9807 ( .I1(n9062), .I2(n9066), .O(n9065) );
  OR_GATE U9808 ( .I1(n9067), .I2(n9063), .O(n9064) );
  AND_GATE U9809 ( .I1(n9065), .I2(n9064), .O(n9072) );
  NAND_GATE U9810 ( .I1(n9066), .I2(n1239), .O(n9070) );
  NAND3_GATE U9811 ( .I1(n9070), .I2(n9069), .I3(n9068), .O(n9071) );
  NAND_GATE U9812 ( .I1(n9072), .I2(n9071), .O(n9522) );
  INV_GATE U9813 ( .I1(n9522), .O(n9525) );
  INV_GATE U9814 ( .I1(n9526), .O(n9523) );
  NAND_GATE U9815 ( .I1(n9530), .I2(n9523), .O(n9073) );
  NAND_GATE U9816 ( .I1(n9525), .I2(n9073), .O(n9074) );
  NAND_GATE U9817 ( .I1(n9521), .I2(n9074), .O(n9579) );
  NAND_GATE U9818 ( .I1(n9578), .I2(n9579), .O(n9076) );
  NAND_GATE U9819 ( .I1(n9075), .I2(n9579), .O(n9574) );
  NAND3_GATE U9820 ( .I1(n9575), .I2(n9076), .I3(n9574), .O(n9512) );
  NAND_GATE U9821 ( .I1(n9510), .I2(n9512), .O(n9507) );
  OR_GATE U9822 ( .I1(n9077), .I2(n9081), .O(n9080) );
  OR_GATE U9823 ( .I1(n9082), .I2(n9078), .O(n9079) );
  NAND_GATE U9824 ( .I1(n9081), .I2(n1166), .O(n9085) );
  NAND3_GATE U9825 ( .I1(n9085), .I2(n9084), .I3(n9083), .O(n9086) );
  INV_GATE U9826 ( .I1(n9508), .O(n9511) );
  INV_GATE U9827 ( .I1(n9512), .O(n9509) );
  NAND_GATE U9828 ( .I1(n9516), .I2(n9509), .O(n9087) );
  NAND_GATE U9829 ( .I1(n9511), .I2(n9087), .O(n9088) );
  NAND_GATE U9830 ( .I1(n9507), .I2(n9088), .O(n9593) );
  NAND_GATE U9831 ( .I1(n9592), .I2(n9593), .O(n9090) );
  NAND_GATE U9832 ( .I1(n9089), .I2(n9593), .O(n9588) );
  NAND3_GATE U9833 ( .I1(n9589), .I2(n9090), .I3(n9588), .O(n9498) );
  NAND_GATE U9834 ( .I1(n9496), .I2(n9498), .O(n9493) );
  OR_GATE U9835 ( .I1(n9091), .I2(n9095), .O(n9094) );
  OR_GATE U9836 ( .I1(n9096), .I2(n9092), .O(n9093) );
  NAND_GATE U9837 ( .I1(n9095), .I2(n1040), .O(n9099) );
  NAND3_GATE U9838 ( .I1(n9099), .I2(n9098), .I3(n9097), .O(n9100) );
  INV_GATE U9839 ( .I1(n9494), .O(n9497) );
  INV_GATE U9840 ( .I1(n9498), .O(n9495) );
  NAND_GATE U9841 ( .I1(n9502), .I2(n9495), .O(n9101) );
  NAND_GATE U9842 ( .I1(n9497), .I2(n9101), .O(n9102) );
  NAND_GATE U9843 ( .I1(n9493), .I2(n9102), .O(n9608) );
  NAND_GATE U9844 ( .I1(n9607), .I2(n9608), .O(n9104) );
  NAND_GATE U9845 ( .I1(n9103), .I2(n9608), .O(n9602) );
  NAND_GATE U9846 ( .I1(n9482), .I2(n9484), .O(n9480) );
  OR_GATE U9847 ( .I1(n9105), .I2(n9109), .O(n9108) );
  OR_GATE U9848 ( .I1(n9110), .I2(n9106), .O(n9107) );
  AND_GATE U9849 ( .I1(n9108), .I2(n9107), .O(n9115) );
  NAND_GATE U9850 ( .I1(n9109), .I2(n1010), .O(n9113) );
  NAND3_GATE U9851 ( .I1(n9113), .I2(n9112), .I3(n9111), .O(n9114) );
  NAND_GATE U9852 ( .I1(n9115), .I2(n9114), .O(n9481) );
  INV_GATE U9853 ( .I1(n9481), .O(n9483) );
  NAND_GATE U9854 ( .I1(n9488), .I2(n826), .O(n9116) );
  NAND_GATE U9855 ( .I1(n9483), .I2(n9116), .O(n9117) );
  NAND_GATE U9856 ( .I1(n9480), .I2(n9117), .O(n9623) );
  NAND_GATE U9857 ( .I1(n9618), .I2(n9623), .O(n9119) );
  NAND_GATE U9858 ( .I1(n1422), .I2(A[11]), .O(n9619) );
  INV_GATE U9859 ( .I1(n9619), .O(n9118) );
  NAND_GATE U9860 ( .I1(n9623), .I2(n9118), .O(n9617) );
  NAND3_GATE U9861 ( .I1(n9622), .I2(n9119), .I3(n9617), .O(n9473) );
  NAND_GATE U9862 ( .I1(n9478), .I2(n9473), .O(n9479) );
  OR_GATE U9863 ( .I1(n9121), .I2(n9120), .O(n9124) );
  OR_GATE U9864 ( .I1(n9129), .I2(n9122), .O(n9123) );
  AND_GATE U9865 ( .I1(n9124), .I2(n9123), .O(n9134) );
  INV_GATE U9866 ( .I1(n9129), .O(n9125) );
  NAND3_GATE U9867 ( .I1(n9125), .I2(n9127), .I3(n9126), .O(n9132) );
  NAND_GATE U9868 ( .I1(n9127), .I2(n9126), .O(n9128) );
  NAND_GATE U9869 ( .I1(n9129), .I2(n9128), .O(n9131) );
  NAND3_GATE U9870 ( .I1(n9132), .I2(n9131), .I3(n9130), .O(n9133) );
  NAND_GATE U9871 ( .I1(n9134), .I2(n9133), .O(n9476) );
  NAND_GATE U9872 ( .I1(n9989), .I2(n9477), .O(n9135) );
  NAND_GATE U9873 ( .I1(n679), .I2(n9135), .O(n9136) );
  NAND_GATE U9874 ( .I1(n9479), .I2(n9136), .O(n9635) );
  NAND_GATE U9875 ( .I1(n9137), .I2(n9635), .O(n9637) );
  NAND3_GATE U9876 ( .I1(n9634), .I2(n9138), .I3(n9637), .O(n9459) );
  NAND_GATE U9877 ( .I1(n9463), .I2(n9459), .O(n9464) );
  OR_GATE U9878 ( .I1(n9140), .I2(n9139), .O(n9148) );
  NAND_GATE U9879 ( .I1(n1030), .I2(n9140), .O(n9141) );
  NAND3_GATE U9880 ( .I1(n9143), .I2(n9142), .I3(n9141), .O(n9147) );
  OR_GATE U9881 ( .I1(n9145), .I2(n9144), .O(n9146) );
  NAND3_GATE U9882 ( .I1(n9148), .I2(n9147), .I3(n9146), .O(n9462) );
  INV_GATE U9883 ( .I1(n9462), .O(n9465) );
  NAND_GATE U9884 ( .I1(n9469), .I2(n362), .O(n9149) );
  NAND_GATE U9885 ( .I1(n9465), .I2(n9149), .O(n9150) );
  NAND_GATE U9886 ( .I1(n9464), .I2(n9150), .O(n9651) );
  NAND_GATE U9887 ( .I1(n9646), .I2(n9651), .O(n9152) );
  NAND_GATE U9888 ( .I1(n1422), .I2(A[15]), .O(n9649) );
  INV_GATE U9889 ( .I1(n9649), .O(n9151) );
  NAND_GATE U9890 ( .I1(n9651), .I2(n9151), .O(n9645) );
  NAND3_GATE U9891 ( .I1(n9650), .I2(n9152), .I3(n9645), .O(n9659) );
  NAND_GATE U9892 ( .I1(n9664), .I2(n9659), .O(n9657) );
  OR_GATE U9893 ( .I1(n9157), .I2(n9153), .O(n9156) );
  OR_GATE U9894 ( .I1(n9154), .I2(n9158), .O(n9155) );
  AND_GATE U9895 ( .I1(n9156), .I2(n9155), .O(n9163) );
  NAND_GATE U9896 ( .I1(n9158), .I2(n1318), .O(n9159) );
  NAND3_GATE U9897 ( .I1(n9161), .I2(n9160), .I3(n9159), .O(n9162) );
  NAND_GATE U9898 ( .I1(n9163), .I2(n9162), .O(n9661) );
  INV_GATE U9899 ( .I1(n9659), .O(n9662) );
  NAND_GATE U9900 ( .I1(n9797), .I2(n9662), .O(n9164) );
  NAND_GATE U9901 ( .I1(n640), .I2(n9164), .O(n9165) );
  NAND_GATE U9902 ( .I1(n9657), .I2(n9165), .O(n9453) );
  NAND_GATE U9903 ( .I1(n9179), .I2(n9453), .O(n9450) );
  NAND3_GATE U9904 ( .I1(n9176), .I2(n9166), .I3(n9167), .O(n9174) );
  NAND_GATE U9905 ( .I1(n9167), .I2(n9176), .O(n9168) );
  NAND_GATE U9906 ( .I1(n9169), .I2(n9168), .O(n9173) );
  NAND_GATE U9907 ( .I1(n9171), .I2(n9170), .O(n9172) );
  NAND3_GATE U9908 ( .I1(n9174), .I2(n9173), .I3(n9172), .O(n9178) );
  OR_GATE U9909 ( .I1(n9176), .I2(n9175), .O(n9177) );
  NAND_GATE U9910 ( .I1(n9178), .I2(n9177), .O(n9454) );
  NAND_GATE U9911 ( .I1(n9453), .I2(n9454), .O(n9180) );
  NAND_GATE U9912 ( .I1(n9179), .I2(n9454), .O(n9449) );
  NAND3_GATE U9913 ( .I1(n9450), .I2(n9180), .I3(n9449), .O(n9676) );
  NAND_GATE U9914 ( .I1(n9776), .I2(n9675), .O(n9181) );
  NAND_GATE U9915 ( .I1(n9676), .I2(n9181), .O(n9182) );
  NAND_GATE U9916 ( .I1(n9196), .I2(n9442), .O(n9444) );
  INV_GATE U9917 ( .I1(n9193), .O(n9187) );
  NAND_GATE U9918 ( .I1(n9188), .I2(n9187), .O(n9183) );
  NAND_GATE U9919 ( .I1(n9184), .I2(n9183), .O(n9191) );
  NAND_GATE U9920 ( .I1(n9185), .I2(n9193), .O(n9190) );
  NAND3_GATE U9921 ( .I1(n9188), .I2(n9187), .I3(n9186), .O(n9189) );
  NAND3_GATE U9922 ( .I1(n9191), .I2(n9190), .I3(n9189), .O(n9195) );
  NAND_GATE U9923 ( .I1(n9195), .I2(n9194), .O(n9445) );
  NAND_GATE U9924 ( .I1(n9196), .I2(n9445), .O(n9443) );
  NAND_GATE U9925 ( .I1(n9442), .I2(n9445), .O(n9197) );
  NAND3_GATE U9926 ( .I1(n9444), .I2(n9443), .I3(n9197), .O(n9685) );
  NAND_GATE U9927 ( .I1(n9757), .I2(n9687), .O(n9198) );
  NAND_GATE U9928 ( .I1(n9685), .I2(n9198), .O(n9199) );
  NAND_GATE U9929 ( .I1(n9683), .I2(n9199), .O(n9432) );
  NAND_GATE U9930 ( .I1(n9200), .I2(n9432), .O(n9422) );
  NAND3_GATE U9931 ( .I1(n9430), .I2(n9432), .I3(n9201), .O(n9202) );
  NAND3_GATE U9932 ( .I1(n9426), .I2(n9422), .I3(n9202), .O(n9415) );
  NAND_GATE U9933 ( .I1(n9210), .I2(n9415), .O(n9403) );
  INV_GATE U9934 ( .I1(n9207), .O(n9206) );
  NAND_GATE U9935 ( .I1(n9203), .I2(n9209), .O(n9402) );
  NAND_GATE U9936 ( .I1(n9206), .I2(n9205), .O(n9209) );
  NAND_GATE U9937 ( .I1(n9207), .I2(n351), .O(n9208) );
  NAND_GATE U9938 ( .I1(n9209), .I2(n9208), .O(n9409) );
  NAND3_GATE U9939 ( .I1(n9210), .I2(n9413), .I3(n9412), .O(n9401) );
  NAND3_GATE U9940 ( .I1(n9415), .I2(n9413), .I3(n9412), .O(n9211) );
  NAND3_GATE U9941 ( .I1(n9403), .I2(n9401), .I3(n9211), .O(n9395) );
  NAND_GATE U9942 ( .I1(n9396), .I2(n9395), .O(n9213) );
  NAND_GATE U9943 ( .I1(n9212), .I2(n9395), .O(n9397) );
  NAND3_GATE U9944 ( .I1(n9394), .I2(n9213), .I3(n9397), .O(n9378) );
  NAND_GATE U9945 ( .I1(n9214), .I2(n9378), .O(n9367) );
  NAND_GATE U9946 ( .I1(n9366), .I2(n9378), .O(n9215) );
  NAND3_GATE U9947 ( .I1(n9368), .I2(n9367), .I3(n9215), .O(n9360) );
  NAND_GATE U9948 ( .I1(n9231), .I2(n9360), .O(n9355) );
  INV_GATE U9949 ( .I1(n9227), .O(n9218) );
  NAND_GATE U9950 ( .I1(n9216), .I2(n9220), .O(n9225) );
  NAND_GATE U9951 ( .I1(n9217), .I2(n9227), .O(n9221) );
  NAND_GATE U9952 ( .I1(n9219), .I2(n9218), .O(n9220) );
  NAND_GATE U9953 ( .I1(n9221), .I2(n9220), .O(n9222) );
  NAND_GATE U9954 ( .I1(n9223), .I2(n9222), .O(n9224) );
  NAND_GATE U9955 ( .I1(n9225), .I2(n9224), .O(n9230) );
  INV_GATE U9956 ( .I1(n9226), .O(n9228) );
  NAND_GATE U9957 ( .I1(n9228), .I2(n9227), .O(n9229) );
  NAND_GATE U9958 ( .I1(n9230), .I2(n9229), .O(n9359) );
  NAND_GATE U9959 ( .I1(n9231), .I2(n9359), .O(n9356) );
  NAND_GATE U9960 ( .I1(n9360), .I2(n9359), .O(n9232) );
  NAND3_GATE U9961 ( .I1(n9355), .I2(n9356), .I3(n9232), .O(n9348) );
  NAND_GATE U9962 ( .I1(n9245), .I2(n9348), .O(n9350) );
  INV_GATE U9963 ( .I1(n9233), .O(n9234) );
  NAND_GATE U9964 ( .I1(n9234), .I2(n9236), .O(n9244) );
  NAND_GATE U9965 ( .I1(n9239), .I2(n9238), .O(n9235) );
  NAND_GATE U9966 ( .I1(n601), .I2(n9235), .O(n9242) );
  NAND_GATE U9967 ( .I1(n9242), .I2(n9241), .O(n9243) );
  NAND_GATE U9968 ( .I1(n9244), .I2(n9243), .O(n9351) );
  NAND_GATE U9969 ( .I1(n9245), .I2(n9351), .O(n9349) );
  NAND_GATE U9970 ( .I1(n9348), .I2(n9351), .O(n9246) );
  NAND3_GATE U9971 ( .I1(n9350), .I2(n9349), .I3(n9246), .O(n9337) );
  NAND_GATE U9972 ( .I1(n9334), .I2(n9337), .O(n9261) );
  INV_GATE U9973 ( .I1(n9247), .O(n9248) );
  NAND_GATE U9974 ( .I1(n9248), .I2(n9251), .O(n9258) );
  NAND_GATE U9975 ( .I1(n9253), .I2(n9252), .O(n9249) );
  NAND_GATE U9976 ( .I1(n9250), .I2(n9249), .O(n9256) );
  NAND_GATE U9977 ( .I1(n9256), .I2(n9255), .O(n9257) );
  NAND_GATE U9978 ( .I1(n9258), .I2(n9257), .O(n9338) );
  NAND_GATE U9979 ( .I1(n9334), .I2(n9338), .O(n9260) );
  NAND_GATE U9980 ( .I1(n9337), .I2(n9338), .O(n9259) );
  NAND3_GATE U9981 ( .I1(n9261), .I2(n9260), .I3(n9259), .O(n9327) );
  NAND_GATE U9982 ( .I1(n9275), .I2(n9327), .O(n9329) );
  INV_GATE U9983 ( .I1(n9262), .O(n9263) );
  NAND_GATE U9984 ( .I1(n9263), .I2(n9266), .O(n9274) );
  NAND_GATE U9985 ( .I1(n9265), .I2(n9268), .O(n9272) );
  NAND_GATE U9986 ( .I1(n901), .I2(n9266), .O(n9267) );
  NAND_GATE U9987 ( .I1(n9268), .I2(n9267), .O(n9269) );
  NAND_GATE U9988 ( .I1(n9270), .I2(n9269), .O(n9271) );
  NAND_GATE U9989 ( .I1(n9272), .I2(n9271), .O(n9273) );
  NAND_GATE U9990 ( .I1(n9274), .I2(n9273), .O(n9330) );
  NAND_GATE U9991 ( .I1(n9275), .I2(n9330), .O(n9328) );
  NAND_GATE U9992 ( .I1(n9327), .I2(n9330), .O(n9276) );
  NAND3_GATE U9993 ( .I1(n9329), .I2(n9328), .I3(n9276), .O(n9318) );
  NAND_GATE U9994 ( .I1(n9288), .I2(n9318), .O(n9313) );
  NAND_GATE U9995 ( .I1(n9278), .I2(n858), .O(n9282) );
  NAND_GATE U9996 ( .I1(n9279), .I2(n9282), .O(n9286) );
  NAND_GATE U9997 ( .I1(n831), .I2(n9280), .O(n9281) );
  NAND_GATE U9998 ( .I1(n9282), .I2(n9281), .O(n9283) );
  NAND_GATE U9999 ( .I1(n9284), .I2(n9283), .O(n9285) );
  NAND_GATE U10000 ( .I1(n9318), .I2(n9317), .O(n9289) );
  NAND3_GATE U10001 ( .I1(n9313), .I2(n9312), .I3(n9289), .O(n9306) );
  NAND_GATE U10002 ( .I1(n9306), .I2(n9305), .O(n9291) );
  NAND_GATE U10003 ( .I1(n9290), .I2(n9306), .O(n9302) );
  AND3_GATE U10004 ( .I1(n9301), .I2(n9291), .I3(n9302), .O(n9298) );
  NAND_GATE U10005 ( .I1(n1423), .I2(A[31]), .O(n9297) );
  NAND_GATE U10006 ( .I1(n9298), .I2(n9297), .O(n9292) );
  NAND_GATE U10007 ( .I1(n9296), .I2(n9292), .O(n9300) );
  INV_GATE U10008 ( .I1(n9300), .O(n14814) );
  NAND_GATE U10009 ( .I1(n9293), .I2(n14814), .O(n9294) );
  NAND_GATE U10010 ( .I1(n9295), .I2(n9294), .O(\A1[42] ) );
  NAND_GATE U10011 ( .I1(n9300), .I2(n9299), .O(n9712) );
  INV_GATE U10012 ( .I1(n9712), .O(n14817) );
  OR_GATE U10013 ( .I1(n9301), .I2(n9306), .O(n9304) );
  OR_GATE U10014 ( .I1(n9305), .I2(n9302), .O(n9303) );
  AND_GATE U10015 ( .I1(n9304), .I2(n9303), .O(n9311) );
  NAND_GATE U10016 ( .I1(n976), .I2(n9305), .O(n9309) );
  NAND3_GATE U10017 ( .I1(n9309), .I2(n9308), .I3(n9307), .O(n9310) );
  OR_GATE U10018 ( .I1(n9312), .I2(n9318), .O(n9315) );
  OR_GATE U10019 ( .I1(n9317), .I2(n9313), .O(n9314) );
  AND_GATE U10020 ( .I1(n9315), .I2(n9314), .O(n9323) );
  INV_GATE U10021 ( .I1(n9318), .O(n9316) );
  NAND_GATE U10022 ( .I1(n9316), .I2(n9317), .O(n9321) );
  NAND_GATE U10023 ( .I1(n9318), .I2(n835), .O(n9320) );
  NAND3_GATE U10024 ( .I1(n9321), .I2(n9320), .I3(n9319), .O(n9322) );
  NAND_GATE U10025 ( .I1(n9323), .I2(n9322), .O(n9721) );
  NAND_GATE U10026 ( .I1(B[11]), .I2(A[30]), .O(n9726) );
  INV_GATE U10027 ( .I1(n9726), .O(n9722) );
  NAND_GATE U10028 ( .I1(n1331), .I2(n9722), .O(n9718) );
  NAND_GATE U10029 ( .I1(n1337), .I2(n9330), .O(n9326) );
  NAND3_GATE U10030 ( .I1(n9326), .I2(n9325), .I3(n9324), .O(n9333) );
  OR_GATE U10031 ( .I1(n9328), .I2(n9327), .O(n9332) );
  OR_GATE U10032 ( .I1(n9330), .I2(n9329), .O(n9331) );
  NAND3_GATE U10033 ( .I1(n9333), .I2(n9332), .I3(n9331), .O(n9733) );
  NAND_GATE U10034 ( .I1(B[11]), .I2(A[29]), .O(n9740) );
  INV_GATE U10035 ( .I1(n9740), .O(n9734) );
  NAND_GATE U10036 ( .I1(n9736), .I2(n9734), .O(n9731) );
  NAND3_GATE U10037 ( .I1(n9337), .I2(n814), .I3(n9334), .O(n9336) );
  INV_GATE U10038 ( .I1(n9337), .O(n9339) );
  NAND3_GATE U10039 ( .I1(n9338), .I2(n9339), .I3(n9334), .O(n9335) );
  AND_GATE U10040 ( .I1(n9336), .I2(n9335), .O(n9344) );
  NAND_GATE U10041 ( .I1(n9257), .I2(n597), .O(n9341) );
  NAND_GATE U10042 ( .I1(n9339), .I2(n9338), .O(n9340) );
  NAND3_GATE U10043 ( .I1(n9342), .I2(n9341), .I3(n9340), .O(n9343) );
  NAND_GATE U10044 ( .I1(n9344), .I2(n9343), .O(n10137) );
  NAND_GATE U10045 ( .I1(B[11]), .I2(A[28]), .O(n10138) );
  INV_GATE U10046 ( .I1(n10138), .O(n10135) );
  NAND_GATE U10047 ( .I1(n806), .I2(n10135), .O(n10132) );
  NAND_GATE U10048 ( .I1(n603), .I2(n9351), .O(n9347) );
  NAND3_GATE U10049 ( .I1(n9347), .I2(n9346), .I3(n9345), .O(n9354) );
  OR_GATE U10050 ( .I1(n9349), .I2(n9348), .O(n9353) );
  OR_GATE U10051 ( .I1(n9351), .I2(n9350), .O(n9352) );
  NAND3_GATE U10052 ( .I1(n9354), .I2(n9353), .I3(n9352), .O(n9750) );
  NAND_GATE U10053 ( .I1(B[11]), .I2(A[27]), .O(n9751) );
  INV_GATE U10054 ( .I1(n9751), .O(n9748) );
  NAND_GATE U10055 ( .I1(n742), .I2(n9748), .O(n9745) );
  NAND_GATE U10056 ( .I1(B[11]), .I2(A[26]), .O(n10119) );
  OR_GATE U10057 ( .I1(n9359), .I2(n9355), .O(n9358) );
  AND_GATE U10058 ( .I1(n9358), .I2(n9357), .O(n9365) );
  NAND_GATE U10059 ( .I1(n958), .I2(n9359), .O(n9362) );
  NAND3_GATE U10060 ( .I1(n9363), .I2(n9362), .I3(n9361), .O(n9364) );
  NAND_GATE U10061 ( .I1(n9365), .I2(n9364), .O(n10121) );
  NAND_GATE U10062 ( .I1(B[11]), .I2(A[25]), .O(n10201) );
  OR_GATE U10063 ( .I1(n9367), .I2(n9366), .O(n9370) );
  INV_GATE U10064 ( .I1(n9371), .O(n9372) );
  NAND_GATE U10065 ( .I1(n9373), .I2(n9372), .O(n9376) );
  NAND3_GATE U10066 ( .I1(n9376), .I2(n358), .I3(n8913), .O(n9381) );
  NAND_GATE U10067 ( .I1(n8913), .I2(n9376), .O(n9377) );
  NAND_GATE U10068 ( .I1(n9378), .I2(n9377), .O(n9380) );
  NAND3_GATE U10069 ( .I1(n9381), .I2(n9380), .I3(n9379), .O(n9382) );
  NAND_GATE U10070 ( .I1(B[11]), .I2(A[24]), .O(n10217) );
  INV_GATE U10071 ( .I1(n10217), .O(n10101) );
  NAND_GATE U10072 ( .I1(n9384), .I2(n9383), .O(n9388) );
  NAND_GATE U10073 ( .I1(n9388), .I2(n9390), .O(n9387) );
  NAND_GATE U10074 ( .I1(n9395), .I2(n9387), .O(n9392) );
  INV_GATE U10075 ( .I1(n9395), .O(n9389) );
  NAND3_GATE U10076 ( .I1(n9390), .I2(n9389), .I3(n9388), .O(n9391) );
  NAND3_GATE U10077 ( .I1(n9393), .I2(n9392), .I3(n9391), .O(n9400) );
  OR_GATE U10078 ( .I1(n9395), .I2(n9394), .O(n9399) );
  OR_GATE U10079 ( .I1(n9397), .I2(n9396), .O(n9398) );
  NAND3_GATE U10080 ( .I1(n9400), .I2(n9399), .I3(n9398), .O(n10104) );
  NAND_GATE U10081 ( .I1(n10101), .I2(n717), .O(n9699) );
  OR_GATE U10082 ( .I1(n9401), .I2(n9415), .O(n9408) );
  NAND_GATE U10083 ( .I1(n9402), .I2(n9412), .O(n9405) );
  INV_GATE U10084 ( .I1(n9403), .O(n9404) );
  NAND3_GATE U10085 ( .I1(n9406), .I2(n9405), .I3(n9404), .O(n9407) );
  AND_GATE U10086 ( .I1(n9408), .I2(n9407), .O(n9420) );
  NAND_GATE U10087 ( .I1(n9410), .I2(n9409), .O(n9412) );
  INV_GATE U10088 ( .I1(n9415), .O(n9411) );
  NAND3_GATE U10089 ( .I1(n9412), .I2(n9411), .I3(n9413), .O(n9418) );
  NAND_GATE U10090 ( .I1(n9413), .I2(n9412), .O(n9414) );
  NAND_GATE U10091 ( .I1(n9415), .I2(n9414), .O(n9417) );
  NAND3_GATE U10092 ( .I1(n9418), .I2(n9417), .I3(n9416), .O(n9419) );
  NAND_GATE U10093 ( .I1(n9420), .I2(n9419), .O(n10093) );
  NAND_GATE U10094 ( .I1(B[11]), .I2(A[23]), .O(n10091) );
  INV_GATE U10095 ( .I1(n10091), .O(n10089) );
  NAND_GATE U10096 ( .I1(n654), .I2(n10089), .O(n10086) );
  NAND_GATE U10097 ( .I1(B[11]), .I2(A[22]), .O(n10245) );
  INV_GATE U10098 ( .I1(n10245), .O(n10077) );
  NAND_GATE U10099 ( .I1(n9421), .I2(n9201), .O(n9425) );
  INV_GATE U10100 ( .I1(n9422), .O(n9424) );
  NAND3_GATE U10101 ( .I1(n9425), .I2(n9424), .I3(n9423), .O(n9438) );
  OR_GATE U10102 ( .I1(n9432), .I2(n9426), .O(n9437) );
  INV_GATE U10103 ( .I1(n9432), .O(n9429) );
  NAND3_GATE U10104 ( .I1(n9201), .I2(n9429), .I3(n9430), .O(n9435) );
  NAND_GATE U10105 ( .I1(n9430), .I2(n9201), .O(n9431) );
  NAND_GATE U10106 ( .I1(n9432), .I2(n9431), .O(n9434) );
  NAND3_GATE U10107 ( .I1(n9435), .I2(n9434), .I3(n9433), .O(n9436) );
  NAND3_GATE U10108 ( .I1(n9438), .I2(n9437), .I3(n9436), .O(n10079) );
  NAND_GATE U10109 ( .I1(n10077), .I2(n718), .O(n10076) );
  NAND_GATE U10110 ( .I1(B[11]), .I2(A[21]), .O(n9766) );
  INV_GATE U10111 ( .I1(n9766), .O(n9691) );
  NAND_GATE U10112 ( .I1(B[11]), .I2(A[20]), .O(n10070) );
  INV_GATE U10113 ( .I1(n10070), .O(n10062) );
  NAND_GATE U10114 ( .I1(n657), .I2(n9445), .O(n9440) );
  NAND3_GATE U10115 ( .I1(n9441), .I2(n9440), .I3(n9439), .O(n9448) );
  OR_GATE U10116 ( .I1(n9443), .I2(n9442), .O(n9447) );
  OR_GATE U10117 ( .I1(n9445), .I2(n9444), .O(n9446) );
  NAND3_GATE U10118 ( .I1(n9448), .I2(n9447), .I3(n9446), .O(n10060) );
  INV_GATE U10119 ( .I1(n10060), .O(n10064) );
  NAND_GATE U10120 ( .I1(n10062), .I2(n10064), .O(n10058) );
  NAND_GATE U10121 ( .I1(B[11]), .I2(A[19]), .O(n9787) );
  INV_GATE U10122 ( .I1(n9787), .O(n9679) );
  NAND_GATE U10123 ( .I1(B[11]), .I2(A[18]), .O(n10041) );
  INV_GATE U10124 ( .I1(n10041), .O(n10045) );
  OR_GATE U10125 ( .I1(n9449), .I2(n9453), .O(n9452) );
  OR_GATE U10126 ( .I1(n9454), .I2(n9450), .O(n9451) );
  NAND_GATE U10127 ( .I1(n1025), .I2(n9454), .O(n9455) );
  NAND3_GATE U10128 ( .I1(n9457), .I2(n9456), .I3(n9455), .O(n9458) );
  INV_GATE U10129 ( .I1(n10043), .O(n10042) );
  NAND_GATE U10130 ( .I1(n10045), .I2(n10042), .O(n10049) );
  NAND_GATE U10131 ( .I1(B[11]), .I2(A[17]), .O(n9804) );
  INV_GATE U10132 ( .I1(n9804), .O(n9667) );
  NAND_GATE U10133 ( .I1(B[11]), .I2(A[16]), .O(n10031) );
  INV_GATE U10134 ( .I1(n10031), .O(n10025) );
  NAND_GATE U10135 ( .I1(n362), .I2(n9462), .O(n9460) );
  NAND_GATE U10136 ( .I1(n9461), .I2(n9460), .O(n9468) );
  NAND_GATE U10137 ( .I1(n9463), .I2(n9460), .O(n9471) );
  INV_GATE U10138 ( .I1(n9464), .O(n9466) );
  NAND_GATE U10139 ( .I1(n9466), .I2(n9465), .O(n9472) );
  NAND4_GATE U10140 ( .I1(n9470), .I2(n9467), .I3(A[15]), .I4(B[11]), .O(
        n10011) );
  NAND_GATE U10141 ( .I1(n9469), .I2(n9468), .O(n9470) );
  NAND_GATE U10142 ( .I1(B[11]), .I2(A[14]), .O(n9817) );
  INV_GATE U10143 ( .I1(n9817), .O(n9810) );
  NAND_GATE U10144 ( .I1(n9477), .I2(n9476), .O(n9475) );
  NAND_GATE U10145 ( .I1(n9473), .I2(n679), .O(n9474) );
  NAND_GATE U10146 ( .I1(n9475), .I2(n9474), .O(n9988) );
  NAND_GATE U10147 ( .I1(n9478), .I2(n9475), .O(n9991) );
  NAND_GATE U10148 ( .I1(B[11]), .I2(A[13]), .O(n10001) );
  INV_GATE U10149 ( .I1(n10001), .O(n9629) );
  NAND3_GATE U10150 ( .I1(n9990), .I2(n9995), .I3(n9629), .O(n10002) );
  NAND_GATE U10151 ( .I1(B[11]), .I2(A[12]), .O(n9830) );
  INV_GATE U10152 ( .I1(n9830), .O(n9824) );
  NAND_GATE U10153 ( .I1(B[11]), .I2(A[11]), .O(n9979) );
  INV_GATE U10154 ( .I1(n9979), .O(n9615) );
  OR_GATE U10155 ( .I1(n9481), .I2(n9480), .O(n9492) );
  NAND_GATE U10156 ( .I1(n826), .I2(n9481), .O(n9486) );
  NAND_GATE U10157 ( .I1(n9482), .I2(n9486), .O(n9490) );
  NAND_GATE U10158 ( .I1(n9486), .I2(n9485), .O(n9487) );
  NAND_GATE U10159 ( .I1(n9488), .I2(n9487), .O(n9489) );
  NAND_GATE U10160 ( .I1(n9490), .I2(n9489), .O(n9491) );
  NAND_GATE U10161 ( .I1(n9492), .I2(n9491), .O(n9977) );
  NAND_GATE U10162 ( .I1(n9615), .I2(n9977), .O(n9974) );
  NAND_GATE U10163 ( .I1(B[11]), .I2(A[10]), .O(n9844) );
  INV_GATE U10164 ( .I1(n9844), .O(n9838) );
  NAND_GATE U10165 ( .I1(B[11]), .I2(A[9]), .O(n9965) );
  INV_GATE U10166 ( .I1(n9965), .O(n9600) );
  OR_GATE U10167 ( .I1(n9494), .I2(n9493), .O(n9506) );
  NAND_GATE U10168 ( .I1(n9495), .I2(n9494), .O(n9500) );
  NAND_GATE U10169 ( .I1(n9496), .I2(n9500), .O(n9504) );
  NAND_GATE U10170 ( .I1(n9498), .I2(n9497), .O(n9499) );
  NAND_GATE U10171 ( .I1(n9500), .I2(n9499), .O(n9501) );
  NAND_GATE U10172 ( .I1(n9502), .I2(n9501), .O(n9503) );
  NAND_GATE U10173 ( .I1(n9504), .I2(n9503), .O(n9505) );
  NAND_GATE U10174 ( .I1(n9506), .I2(n9505), .O(n9963) );
  NAND_GATE U10175 ( .I1(n9600), .I2(n9963), .O(n9960) );
  NAND_GATE U10176 ( .I1(B[11]), .I2(A[8]), .O(n9858) );
  INV_GATE U10177 ( .I1(n9858), .O(n9852) );
  NAND_GATE U10178 ( .I1(B[11]), .I2(A[7]), .O(n9951) );
  INV_GATE U10179 ( .I1(n9951), .O(n9586) );
  OR_GATE U10180 ( .I1(n9508), .I2(n9507), .O(n9520) );
  NAND_GATE U10181 ( .I1(n9509), .I2(n9508), .O(n9514) );
  NAND_GATE U10182 ( .I1(n9510), .I2(n9514), .O(n9518) );
  NAND_GATE U10183 ( .I1(n9512), .I2(n9511), .O(n9513) );
  NAND_GATE U10184 ( .I1(n9514), .I2(n9513), .O(n9515) );
  NAND_GATE U10185 ( .I1(n9516), .I2(n9515), .O(n9517) );
  NAND_GATE U10186 ( .I1(n9518), .I2(n9517), .O(n9519) );
  NAND_GATE U10187 ( .I1(n9520), .I2(n9519), .O(n9949) );
  NAND_GATE U10188 ( .I1(n9586), .I2(n9949), .O(n9946) );
  NAND_GATE U10189 ( .I1(B[11]), .I2(A[6]), .O(n9872) );
  INV_GATE U10190 ( .I1(n9872), .O(n9866) );
  OR_GATE U10191 ( .I1(n9522), .I2(n9521), .O(n9534) );
  NAND_GATE U10192 ( .I1(n9523), .I2(n9522), .O(n9528) );
  NAND_GATE U10193 ( .I1(n9524), .I2(n9528), .O(n9532) );
  NAND_GATE U10194 ( .I1(n9526), .I2(n9525), .O(n9527) );
  NAND_GATE U10195 ( .I1(n9528), .I2(n9527), .O(n9529) );
  NAND_GATE U10196 ( .I1(n9530), .I2(n9529), .O(n9531) );
  NAND_GATE U10197 ( .I1(n9532), .I2(n9531), .O(n9533) );
  NAND_GATE U10198 ( .I1(n9534), .I2(n9533), .O(n9881) );
  OR_GATE U10199 ( .I1(n9535), .I2(n9539), .O(n9538) );
  OR_GATE U10200 ( .I1(n9536), .I2(n9540), .O(n9537) );
  AND_GATE U10201 ( .I1(n9538), .I2(n9537), .O(n9545) );
  NAND_GATE U10202 ( .I1(n9539), .I2(n1240), .O(n9543) );
  NAND3_GATE U10203 ( .I1(n9543), .I2(n9542), .I3(n9541), .O(n9544) );
  NAND_GATE U10204 ( .I1(n9545), .I2(n9544), .O(n9890) );
  INV_GATE U10205 ( .I1(n9890), .O(n9893) );
  INV_GATE U10206 ( .I1(n9546), .O(n9547) );
  NAND_GATE U10207 ( .I1(n9551), .I2(n9547), .O(n9559) );
  NAND_GATE U10208 ( .I1(n9549), .I2(n9553), .O(n9557) );
  NAND_GATE U10209 ( .I1(n9551), .I2(n9550), .O(n9552) );
  NAND_GATE U10210 ( .I1(n9553), .I2(n9552), .O(n9554) );
  NAND_GATE U10211 ( .I1(n9555), .I2(n9554), .O(n9556) );
  NAND_GATE U10212 ( .I1(n9557), .I2(n9556), .O(n9558) );
  NAND_GATE U10213 ( .I1(n9559), .I2(n9558), .O(n9906) );
  NAND_GATE U10214 ( .I1(n1423), .I2(A[0]), .O(n9560) );
  NAND_GATE U10215 ( .I1(n14241), .I2(n9560), .O(n9561) );
  NAND_GATE U10216 ( .I1(B[13]), .I2(n9561), .O(n9565) );
  NAND_GATE U10217 ( .I1(n1424), .I2(A[1]), .O(n9562) );
  NAND_GATE U10218 ( .I1(n724), .I2(n9562), .O(n9563) );
  NAND_GATE U10219 ( .I1(n1422), .I2(n9563), .O(n9564) );
  NAND_GATE U10220 ( .I1(n9565), .I2(n9564), .O(n9918) );
  NAND_GATE U10221 ( .I1(B[11]), .I2(A[2]), .O(n9922) );
  NAND3_GATE U10222 ( .I1(B[11]), .I2(n1422), .I3(n1254), .O(n9915) );
  NAND_GATE U10223 ( .I1(n9922), .I2(n9915), .O(n9566) );
  NAND_GATE U10224 ( .I1(n9918), .I2(n9566), .O(n9567) );
  INV_GATE U10225 ( .I1(n9922), .O(n9916) );
  INV_GATE U10226 ( .I1(n9915), .O(n9917) );
  NAND_GATE U10227 ( .I1(n9916), .I2(n9917), .O(n9913) );
  NAND_GATE U10228 ( .I1(n9567), .I2(n9913), .O(n9907) );
  NAND_GATE U10229 ( .I1(n9906), .I2(n9907), .O(n9569) );
  NAND_GATE U10230 ( .I1(B[11]), .I2(A[3]), .O(n9908) );
  INV_GATE U10231 ( .I1(n9908), .O(n9568) );
  NAND_GATE U10232 ( .I1(n9906), .I2(n9568), .O(n9903) );
  NAND_GATE U10233 ( .I1(n9907), .I2(n9568), .O(n9902) );
  NAND3_GATE U10234 ( .I1(n9569), .I2(n9903), .I3(n9902), .O(n9892) );
  INV_GATE U10235 ( .I1(n9892), .O(n9889) );
  NAND_GATE U10236 ( .I1(B[11]), .I2(A[4]), .O(n9897) );
  NAND_GATE U10237 ( .I1(n9889), .I2(n9897), .O(n9570) );
  NAND_GATE U10238 ( .I1(n9893), .I2(n9570), .O(n9571) );
  INV_GATE U10239 ( .I1(n9897), .O(n9891) );
  NAND_GATE U10240 ( .I1(n9892), .I2(n9891), .O(n9888) );
  NAND_GATE U10241 ( .I1(n9571), .I2(n9888), .O(n9882) );
  NAND_GATE U10242 ( .I1(n9881), .I2(n9882), .O(n9573) );
  NAND_GATE U10243 ( .I1(B[11]), .I2(A[5]), .O(n9883) );
  INV_GATE U10244 ( .I1(n9883), .O(n9572) );
  NAND_GATE U10245 ( .I1(n9881), .I2(n9572), .O(n9878) );
  NAND_GATE U10246 ( .I1(n9882), .I2(n9572), .O(n9877) );
  NAND3_GATE U10247 ( .I1(n9573), .I2(n9878), .I3(n9877), .O(n9868) );
  NAND_GATE U10248 ( .I1(n9866), .I2(n9868), .O(n9863) );
  OR_GATE U10249 ( .I1(n9574), .I2(n9578), .O(n9577) );
  OR_GATE U10250 ( .I1(n9579), .I2(n9575), .O(n9576) );
  NAND_GATE U10251 ( .I1(n9578), .I2(n1170), .O(n9582) );
  NAND3_GATE U10252 ( .I1(n9582), .I2(n9581), .I3(n9580), .O(n9583) );
  INV_GATE U10253 ( .I1(n9864), .O(n9867) );
  INV_GATE U10254 ( .I1(n9868), .O(n9865) );
  NAND_GATE U10255 ( .I1(n9872), .I2(n9865), .O(n9584) );
  NAND_GATE U10256 ( .I1(n9867), .I2(n9584), .O(n9585) );
  NAND_GATE U10257 ( .I1(n9863), .I2(n9585), .O(n9950) );
  NAND_GATE U10258 ( .I1(n9949), .I2(n9950), .O(n9587) );
  NAND_GATE U10259 ( .I1(n9586), .I2(n9950), .O(n9945) );
  NAND3_GATE U10260 ( .I1(n9946), .I2(n9587), .I3(n9945), .O(n9854) );
  NAND_GATE U10261 ( .I1(n9852), .I2(n9854), .O(n9849) );
  OR_GATE U10262 ( .I1(n9588), .I2(n9592), .O(n9591) );
  OR_GATE U10263 ( .I1(n9593), .I2(n9589), .O(n9590) );
  NAND_GATE U10264 ( .I1(n9592), .I2(n1053), .O(n9596) );
  NAND3_GATE U10265 ( .I1(n9596), .I2(n9595), .I3(n9594), .O(n9597) );
  INV_GATE U10266 ( .I1(n9850), .O(n9853) );
  INV_GATE U10267 ( .I1(n9854), .O(n9851) );
  NAND_GATE U10268 ( .I1(n9858), .I2(n9851), .O(n9598) );
  NAND_GATE U10269 ( .I1(n9853), .I2(n9598), .O(n9599) );
  NAND_GATE U10270 ( .I1(n9849), .I2(n9599), .O(n9964) );
  NAND_GATE U10271 ( .I1(n9963), .I2(n9964), .O(n9601) );
  NAND_GATE U10272 ( .I1(n9600), .I2(n9964), .O(n9959) );
  NAND3_GATE U10273 ( .I1(n9960), .I2(n9601), .I3(n9959), .O(n9840) );
  NAND_GATE U10274 ( .I1(n9838), .I2(n9840), .O(n9835) );
  OR_GATE U10275 ( .I1(n9602), .I2(n9607), .O(n9605) );
  OR_GATE U10276 ( .I1(n9608), .I2(n9603), .O(n9604) );
  INV_GATE U10277 ( .I1(n9608), .O(n9606) );
  NAND_GATE U10278 ( .I1(n9607), .I2(n9606), .O(n9611) );
  NAND_GATE U10279 ( .I1(n1311), .I2(n9608), .O(n9610) );
  NAND3_GATE U10280 ( .I1(n9611), .I2(n9610), .I3(n9609), .O(n9612) );
  INV_GATE U10281 ( .I1(n9836), .O(n9839) );
  INV_GATE U10282 ( .I1(n9840), .O(n9837) );
  NAND_GATE U10283 ( .I1(n9844), .I2(n9837), .O(n9613) );
  NAND_GATE U10284 ( .I1(n9839), .I2(n9613), .O(n9614) );
  NAND_GATE U10285 ( .I1(n9835), .I2(n9614), .O(n9978) );
  NAND_GATE U10286 ( .I1(n9977), .I2(n9978), .O(n9616) );
  NAND_GATE U10287 ( .I1(n9615), .I2(n9978), .O(n9973) );
  NAND3_GATE U10288 ( .I1(n9974), .I2(n9616), .I3(n9973), .O(n9826) );
  NAND_GATE U10289 ( .I1(n9824), .I2(n9826), .O(n9822) );
  OR_GATE U10290 ( .I1(n9617), .I2(n9618), .O(n9626) );
  NAND_GATE U10291 ( .I1(n9618), .I2(n664), .O(n9621) );
  NAND3_GATE U10292 ( .I1(n9621), .I2(n9620), .I3(n9619), .O(n9625) );
  OR_GATE U10293 ( .I1(n9623), .I2(n9622), .O(n9624) );
  NAND3_GATE U10294 ( .I1(n9626), .I2(n9625), .I3(n9624), .O(n9823) );
  INV_GATE U10295 ( .I1(n9823), .O(n9825) );
  NAND_GATE U10296 ( .I1(n9830), .I2(n1310), .O(n9627) );
  NAND_GATE U10297 ( .I1(n9825), .I2(n9627), .O(n9628) );
  NAND_GATE U10298 ( .I1(n9822), .I2(n9628), .O(n10003) );
  NAND3_GATE U10299 ( .I1(n10003), .I2(n9990), .I3(n9995), .O(n9630) );
  NAND_GATE U10300 ( .I1(n9629), .I2(n10003), .O(n9994) );
  NAND3_GATE U10301 ( .I1(n10002), .I2(n9630), .I3(n9994), .O(n9812) );
  NAND_GATE U10302 ( .I1(n9810), .I2(n9812), .O(n9819) );
  NAND_GATE U10303 ( .I1(n9636), .I2(n1029), .O(n9631) );
  NAND3_GATE U10304 ( .I1(n9633), .I2(n9632), .I3(n9631), .O(n9640) );
  OR_GATE U10305 ( .I1(n9635), .I2(n9634), .O(n9639) );
  OR_GATE U10306 ( .I1(n9637), .I2(n9636), .O(n9638) );
  NAND3_GATE U10307 ( .I1(n9640), .I2(n9639), .I3(n9638), .O(n9820) );
  INV_GATE U10308 ( .I1(n9820), .O(n9811) );
  INV_GATE U10309 ( .I1(n9812), .O(n9813) );
  NAND_GATE U10310 ( .I1(n9817), .I2(n9813), .O(n9641) );
  NAND_GATE U10311 ( .I1(n9811), .I2(n9641), .O(n9642) );
  NAND_GATE U10312 ( .I1(n9819), .I2(n9642), .O(n10015) );
  NAND_GATE U10313 ( .I1(n10016), .I2(n10015), .O(n9644) );
  NAND_GATE U10314 ( .I1(B[11]), .I2(A[15]), .O(n10019) );
  INV_GATE U10315 ( .I1(n10019), .O(n9643) );
  NAND_GATE U10316 ( .I1(n10015), .I2(n9643), .O(n10012) );
  NAND3_GATE U10317 ( .I1(n10011), .I2(n9644), .I3(n10012), .O(n10027) );
  NAND_GATE U10318 ( .I1(n10025), .I2(n10027), .O(n10034) );
  OR_GATE U10319 ( .I1(n9645), .I2(n9646), .O(n9654) );
  NAND_GATE U10320 ( .I1(n9646), .I2(n1027), .O(n9647) );
  NAND3_GATE U10321 ( .I1(n9649), .I2(n9648), .I3(n9647), .O(n9653) );
  OR_GATE U10322 ( .I1(n9651), .I2(n9650), .O(n9652) );
  NAND3_GATE U10323 ( .I1(n9654), .I2(n9653), .I3(n9652), .O(n10035) );
  INV_GATE U10324 ( .I1(n10035), .O(n10026) );
  INV_GATE U10325 ( .I1(n10027), .O(n10028) );
  NAND_GATE U10326 ( .I1(n10026), .I2(n9655), .O(n9656) );
  NAND_GATE U10327 ( .I1(n10034), .I2(n9656), .O(n9799) );
  NAND_GATE U10328 ( .I1(n9667), .I2(n9799), .O(n9805) );
  INV_GATE U10329 ( .I1(n9657), .O(n9658) );
  NAND_GATE U10330 ( .I1(n9659), .I2(n640), .O(n9660) );
  NAND_GATE U10331 ( .I1(n9660), .I2(n9663), .O(n9796) );
  NAND_GATE U10332 ( .I1(n9662), .I2(n9661), .O(n9663) );
  NAND_GATE U10333 ( .I1(n9664), .I2(n9663), .O(n9794) );
  NAND_GATE U10334 ( .I1(n9665), .I2(n9794), .O(n9666) );
  NAND_GATE U10335 ( .I1(n9795), .I2(n9666), .O(n9806) );
  NAND_GATE U10336 ( .I1(n9799), .I2(n9806), .O(n9668) );
  NAND_GATE U10337 ( .I1(n9667), .I2(n9806), .O(n9793) );
  NAND_GATE U10338 ( .I1(n10041), .I2(n10043), .O(n9669) );
  NAND_GATE U10339 ( .I1(n10050), .I2(n9669), .O(n9670) );
  NAND_GATE U10340 ( .I1(n10049), .I2(n9670), .O(n9786) );
  NAND_GATE U10341 ( .I1(n9679), .I2(n9786), .O(n9779) );
  INV_GATE U10342 ( .I1(n9676), .O(n9674) );
  NAND_GATE U10343 ( .I1(n9671), .I2(n9678), .O(n9778) );
  INV_GATE U10344 ( .I1(n9778), .O(n9673) );
  NAND_GATE U10345 ( .I1(n9673), .I2(n9780), .O(n9784) );
  NAND_GATE U10346 ( .I1(n9675), .I2(n9674), .O(n9678) );
  NAND_GATE U10347 ( .I1(n394), .I2(n9676), .O(n9677) );
  NAND_GATE U10348 ( .I1(n9678), .I2(n9677), .O(n9775) );
  NAND3_GATE U10349 ( .I1(n9786), .I2(n9784), .I3(n9777), .O(n9680) );
  NAND3_GATE U10350 ( .I1(n9679), .I2(n9784), .I3(n9777), .O(n9774) );
  NAND3_GATE U10351 ( .I1(n9779), .I2(n9680), .I3(n9774), .O(n10063) );
  NAND_GATE U10352 ( .I1(n10070), .I2(n10060), .O(n9681) );
  NAND_GATE U10353 ( .I1(n10063), .I2(n9681), .O(n9682) );
  NAND_GATE U10354 ( .I1(n10058), .I2(n9682), .O(n9767) );
  NAND_GATE U10355 ( .I1(n9691), .I2(n9767), .O(n9769) );
  INV_GATE U10356 ( .I1(n9685), .O(n9686) );
  NAND_GATE U10357 ( .I1(n9684), .I2(n9688), .O(n9758) );
  NAND_GATE U10358 ( .I1(n875), .I2(n9685), .O(n9689) );
  NAND_GATE U10359 ( .I1(n9687), .I2(n9686), .O(n9688) );
  NAND_GATE U10360 ( .I1(n9689), .I2(n9688), .O(n9756) );
  NAND_GATE U10361 ( .I1(n9758), .I2(n9761), .O(n9690) );
  NAND_GATE U10362 ( .I1(n9759), .I2(n9690), .O(n9770) );
  NAND_GATE U10363 ( .I1(n9767), .I2(n9770), .O(n9692) );
  NAND3_GATE U10364 ( .I1(n9769), .I2(n9768), .I3(n9692), .O(n10078) );
  NAND_GATE U10365 ( .I1(n10245), .I2(n10079), .O(n9693) );
  NAND_GATE U10366 ( .I1(n10078), .I2(n9693), .O(n9694) );
  NAND_GATE U10367 ( .I1(n10076), .I2(n9694), .O(n10090) );
  NAND_GATE U10368 ( .I1(n10093), .I2(n10091), .O(n9695) );
  NAND_GATE U10369 ( .I1(n10090), .I2(n9695), .O(n9696) );
  NAND_GATE U10370 ( .I1(n10086), .I2(n9696), .O(n10102) );
  NAND_GATE U10371 ( .I1(n10217), .I2(n10104), .O(n9697) );
  NAND_GATE U10372 ( .I1(n10102), .I2(n9697), .O(n9698) );
  NAND_GATE U10373 ( .I1(n9699), .I2(n9698), .O(n10113) );
  NAND_GATE U10374 ( .I1(n10201), .I2(n10114), .O(n9700) );
  NAND_GATE U10375 ( .I1(n10113), .I2(n9700), .O(n9701) );
  NAND_GATE U10376 ( .I1(n10111), .I2(n9701), .O(n10125) );
  NAND_GATE U10377 ( .I1(n10119), .I2(n10121), .O(n9702) );
  NAND_GATE U10378 ( .I1(n9750), .I2(n9751), .O(n9703) );
  NAND_GATE U10379 ( .I1(n9749), .I2(n9703), .O(n9704) );
  NAND_GATE U10380 ( .I1(n9745), .I2(n9704), .O(n10136) );
  NAND_GATE U10381 ( .I1(n10137), .I2(n10138), .O(n9705) );
  NAND_GATE U10382 ( .I1(n10136), .I2(n9705), .O(n9706) );
  NAND_GATE U10383 ( .I1(n10132), .I2(n9706), .O(n9735) );
  NAND_GATE U10384 ( .I1(n9733), .I2(n9740), .O(n9707) );
  NAND_GATE U10385 ( .I1(n9735), .I2(n9707), .O(n9708) );
  NAND_GATE U10386 ( .I1(n9731), .I2(n9708), .O(n9723) );
  NAND_GATE U10387 ( .I1(n9721), .I2(n9726), .O(n9709) );
  NAND_GATE U10388 ( .I1(n9723), .I2(n9709), .O(n9711) );
  NAND_GATE U10389 ( .I1(n1421), .I2(A[31]), .O(n9710) );
  NAND3_GATE U10390 ( .I1(n9718), .I2(n9711), .I3(n9710), .O(n9715) );
  INV_GATE U10391 ( .I1(n9717), .O(n14816) );
  NAND_GATE U10392 ( .I1(n9712), .I2(n14816), .O(n9713) );
  NAND_GATE U10393 ( .I1(n9714), .I2(n9713), .O(\A1[41] ) );
  NAND_GATE U10394 ( .I1(n9717), .I2(n9716), .O(n10148) );
  INV_GATE U10395 ( .I1(n10148), .O(n14818) );
  INV_GATE U10396 ( .I1(n9718), .O(n9719) );
  NAND_GATE U10397 ( .I1(n9719), .I2(n9723), .O(n9730) );
  INV_GATE U10398 ( .I1(n9723), .O(n9720) );
  NAND_GATE U10399 ( .I1(n9721), .I2(n9720), .O(n9725) );
  NAND_GATE U10400 ( .I1(n9722), .I2(n9725), .O(n9728) );
  NAND_GATE U10401 ( .I1(n1331), .I2(n9723), .O(n9724) );
  NAND_GATE U10402 ( .I1(n9728), .I2(n9727), .O(n9729) );
  NAND_GATE U10403 ( .I1(n9730), .I2(n9729), .O(n10151) );
  NAND_GATE U10404 ( .I1(B[10]), .I2(A[30]), .O(n10156) );
  INV_GATE U10405 ( .I1(n10156), .O(n10145) );
  INV_GATE U10406 ( .I1(n9731), .O(n9732) );
  NAND_GATE U10407 ( .I1(n9732), .I2(n9735), .O(n9744) );
  NAND_GATE U10408 ( .I1(n9734), .I2(n9738), .O(n9742) );
  NAND_GATE U10409 ( .I1(n9736), .I2(n9735), .O(n9737) );
  NAND_GATE U10410 ( .I1(n9738), .I2(n9737), .O(n9739) );
  NAND_GATE U10411 ( .I1(n9740), .I2(n9739), .O(n9741) );
  NAND_GATE U10412 ( .I1(n9742), .I2(n9741), .O(n9743) );
  NAND_GATE U10413 ( .I1(n9744), .I2(n9743), .O(n10162) );
  NAND_GATE U10414 ( .I1(n10145), .I2(n10162), .O(n10160) );
  NAND_GATE U10415 ( .I1(B[10]), .I2(A[29]), .O(n10175) );
  INV_GATE U10416 ( .I1(n10175), .O(n10166) );
  NAND_GATE U10417 ( .I1(B[10]), .I2(A[28]), .O(n10186) );
  INV_GATE U10418 ( .I1(n10186), .O(n10178) );
  INV_GATE U10419 ( .I1(n9745), .O(n9746) );
  NAND_GATE U10420 ( .I1(n9746), .I2(n9749), .O(n9755) );
  NAND_GATE U10421 ( .I1(n9748), .I2(n9747), .O(n9753) );
  NAND_GATE U10422 ( .I1(n9753), .I2(n9752), .O(n9754) );
  NAND_GATE U10423 ( .I1(n9755), .I2(n9754), .O(n10182) );
  NAND_GATE U10424 ( .I1(n10178), .I2(n10182), .O(n10131) );
  NAND_GATE U10425 ( .I1(B[10]), .I2(A[27]), .O(n10196) );
  INV_GATE U10426 ( .I1(n10196), .O(n10189) );
  NAND_GATE U10427 ( .I1(B[10]), .I2(A[26]), .O(n10208) );
  INV_GATE U10428 ( .I1(n10208), .O(n10210) );
  NAND_GATE U10429 ( .I1(B[10]), .I2(A[25]), .O(n10223) );
  INV_GATE U10430 ( .I1(n10223), .O(n10227) );
  NAND_GATE U10431 ( .I1(B[10]), .I2(A[24]), .O(n10239) );
  INV_GATE U10432 ( .I1(n10239), .O(n10099) );
  NAND_GATE U10433 ( .I1(B[10]), .I2(A[23]), .O(n10249) );
  INV_GATE U10434 ( .I1(n10249), .O(n10084) );
  NAND_GATE U10435 ( .I1(B[10]), .I2(A[22]), .O(n10604) );
  INV_GATE U10436 ( .I1(n10604), .O(n10260) );
  NAND_GATE U10437 ( .I1(n9757), .I2(n9756), .O(n9761) );
  NAND_GATE U10438 ( .I1(n9759), .I2(n3), .O(n9763) );
  NAND_GATE U10439 ( .I1(n9761), .I2(n9763), .O(n9760) );
  NAND_GATE U10440 ( .I1(n9767), .I2(n9760), .O(n9765) );
  INV_GATE U10441 ( .I1(n9767), .O(n9762) );
  NAND3_GATE U10442 ( .I1(n9763), .I2(n9762), .I3(n9761), .O(n9764) );
  NAND3_GATE U10443 ( .I1(n9766), .I2(n9765), .I3(n9764), .O(n9773) );
  OR_GATE U10444 ( .I1(n9768), .I2(n9767), .O(n9772) );
  OR_GATE U10445 ( .I1(n9770), .I2(n9769), .O(n9771) );
  NAND3_GATE U10446 ( .I1(n9773), .I2(n9772), .I3(n9771), .O(n10257) );
  NAND_GATE U10447 ( .I1(n10260), .I2(n874), .O(n10075) );
  NAND_GATE U10448 ( .I1(B[10]), .I2(A[21]), .O(n10264) );
  INV_GATE U10449 ( .I1(n10264), .O(n10068) );
  OR_GATE U10450 ( .I1(n9774), .I2(n9786), .O(n9792) );
  NAND_GATE U10451 ( .I1(n9776), .I2(n9775), .O(n9777) );
  NAND_GATE U10452 ( .I1(n9778), .I2(n9777), .O(n9782) );
  INV_GATE U10453 ( .I1(n9779), .O(n9781) );
  NAND3_GATE U10454 ( .I1(n9782), .I2(n9781), .I3(n9780), .O(n9791) );
  INV_GATE U10455 ( .I1(n9786), .O(n9783) );
  NAND3_GATE U10456 ( .I1(n9784), .I2(n9777), .I3(n9783), .O(n9789) );
  NAND_GATE U10457 ( .I1(n9784), .I2(n9777), .O(n9785) );
  NAND_GATE U10458 ( .I1(n9786), .I2(n9785), .O(n9788) );
  NAND3_GATE U10459 ( .I1(n9789), .I2(n9788), .I3(n9787), .O(n9790) );
  NAND3_GATE U10460 ( .I1(n9792), .I2(n9791), .I3(n9790), .O(n10534) );
  NAND_GATE U10461 ( .I1(B[10]), .I2(A[20]), .O(n10531) );
  INV_GATE U10462 ( .I1(n10531), .O(n10536) );
  NAND_GATE U10463 ( .I1(n393), .I2(n10536), .O(n10529) );
  NAND_GATE U10464 ( .I1(B[10]), .I2(A[19]), .O(n10277) );
  INV_GATE U10465 ( .I1(n10277), .O(n10054) );
  OR_GATE U10466 ( .I1(n99), .I2(n72), .O(n9809) );
  NAND_GATE U10467 ( .I1(n9797), .I2(n9796), .O(n9800) );
  NAND_GATE U10468 ( .I1(n9801), .I2(n9800), .O(n9798) );
  NAND_GATE U10469 ( .I1(n9799), .I2(n9798), .O(n9803) );
  NAND3_GATE U10470 ( .I1(n9804), .I2(n9803), .I3(n9802), .O(n9808) );
  OR_GATE U10471 ( .I1(n9806), .I2(n9805), .O(n9807) );
  NAND3_GATE U10472 ( .I1(n9809), .I2(n9808), .I3(n9807), .O(n10291) );
  INV_GATE U10473 ( .I1(n10291), .O(n10287) );
  NAND_GATE U10474 ( .I1(B[10]), .I2(A[18]), .O(n10290) );
  INV_GATE U10475 ( .I1(n10290), .O(n10285) );
  NAND_GATE U10476 ( .I1(n10287), .I2(n10285), .O(n10283) );
  NAND_GATE U10477 ( .I1(B[10]), .I2(A[17]), .O(n10300) );
  INV_GATE U10478 ( .I1(n10300), .O(n10037) );
  NAND_GATE U10479 ( .I1(B[10]), .I2(A[16]), .O(n10507) );
  INV_GATE U10480 ( .I1(n10507), .O(n10512) );
  NAND_GATE U10481 ( .I1(n9810), .I2(n9814), .O(n9818) );
  NAND_GATE U10482 ( .I1(n9812), .I2(n9811), .O(n9815) );
  NAND_GATE U10483 ( .I1(n9813), .I2(n9820), .O(n9814) );
  NAND_GATE U10484 ( .I1(n9815), .I2(n9814), .O(n9816) );
  OR_GATE U10485 ( .I1(n9820), .I2(n9819), .O(n9821) );
  NAND3_GATE U10486 ( .I1(A[15]), .I2(n10497), .I3(B[10]), .O(n10501) );
  NAND_GATE U10487 ( .I1(B[10]), .I2(A[14]), .O(n10311) );
  INV_GATE U10488 ( .I1(n10311), .O(n10304) );
  NAND_GATE U10489 ( .I1(B[10]), .I2(A[13]), .O(n10488) );
  INV_GATE U10490 ( .I1(n10488), .O(n9986) );
  OR_GATE U10491 ( .I1(n9823), .I2(n9822), .O(n9834) );
  NAND_GATE U10492 ( .I1(n1310), .I2(n9823), .O(n9828) );
  NAND_GATE U10493 ( .I1(n9824), .I2(n9828), .O(n9832) );
  NAND_GATE U10494 ( .I1(n9826), .I2(n9825), .O(n9827) );
  NAND_GATE U10495 ( .I1(n9828), .I2(n9827), .O(n9829) );
  NAND_GATE U10496 ( .I1(n9830), .I2(n9829), .O(n9831) );
  NAND_GATE U10497 ( .I1(n9832), .I2(n9831), .O(n9833) );
  NAND_GATE U10498 ( .I1(n9834), .I2(n9833), .O(n10486) );
  NAND_GATE U10499 ( .I1(n9986), .I2(n10486), .O(n10483) );
  NAND_GATE U10500 ( .I1(B[10]), .I2(A[12]), .O(n10324) );
  INV_GATE U10501 ( .I1(n10324), .O(n10319) );
  NAND_GATE U10502 ( .I1(B[10]), .I2(A[11]), .O(n10473) );
  INV_GATE U10503 ( .I1(n10473), .O(n9971) );
  OR_GATE U10504 ( .I1(n9836), .I2(n9835), .O(n9848) );
  NAND_GATE U10505 ( .I1(n9837), .I2(n9836), .O(n9842) );
  NAND_GATE U10506 ( .I1(n9838), .I2(n9842), .O(n9846) );
  NAND_GATE U10507 ( .I1(n9840), .I2(n9839), .O(n9841) );
  NAND_GATE U10508 ( .I1(n9842), .I2(n9841), .O(n9843) );
  NAND_GATE U10509 ( .I1(n9844), .I2(n9843), .O(n9845) );
  NAND_GATE U10510 ( .I1(n9846), .I2(n9845), .O(n9847) );
  NAND_GATE U10511 ( .I1(n9848), .I2(n9847), .O(n10471) );
  NAND_GATE U10512 ( .I1(n9971), .I2(n10471), .O(n10468) );
  NAND_GATE U10513 ( .I1(B[10]), .I2(A[10]), .O(n10338) );
  INV_GATE U10514 ( .I1(n10338), .O(n10332) );
  NAND_GATE U10515 ( .I1(B[10]), .I2(A[9]), .O(n10459) );
  INV_GATE U10516 ( .I1(n10459), .O(n9957) );
  OR_GATE U10517 ( .I1(n9850), .I2(n9849), .O(n9862) );
  NAND_GATE U10518 ( .I1(n9851), .I2(n9850), .O(n9856) );
  NAND_GATE U10519 ( .I1(n9852), .I2(n9856), .O(n9860) );
  NAND_GATE U10520 ( .I1(n9854), .I2(n9853), .O(n9855) );
  NAND_GATE U10521 ( .I1(n9856), .I2(n9855), .O(n9857) );
  NAND_GATE U10522 ( .I1(n9858), .I2(n9857), .O(n9859) );
  NAND_GATE U10523 ( .I1(n9860), .I2(n9859), .O(n9861) );
  NAND_GATE U10524 ( .I1(n9862), .I2(n9861), .O(n10457) );
  NAND_GATE U10525 ( .I1(n9957), .I2(n10457), .O(n10454) );
  NAND_GATE U10526 ( .I1(B[10]), .I2(A[8]), .O(n10352) );
  INV_GATE U10527 ( .I1(n10352), .O(n10346) );
  OR_GATE U10528 ( .I1(n9864), .I2(n9863), .O(n9876) );
  NAND_GATE U10529 ( .I1(n9865), .I2(n9864), .O(n9870) );
  NAND_GATE U10530 ( .I1(n9866), .I2(n9870), .O(n9874) );
  NAND_GATE U10531 ( .I1(n9868), .I2(n9867), .O(n9869) );
  NAND_GATE U10532 ( .I1(n9870), .I2(n9869), .O(n9871) );
  NAND_GATE U10533 ( .I1(n9872), .I2(n9871), .O(n9873) );
  NAND_GATE U10534 ( .I1(n9874), .I2(n9873), .O(n9875) );
  NAND_GATE U10535 ( .I1(n9876), .I2(n9875), .O(n10361) );
  OR_GATE U10536 ( .I1(n9877), .I2(n9881), .O(n9880) );
  OR_GATE U10537 ( .I1(n9878), .I2(n9882), .O(n9879) );
  AND_GATE U10538 ( .I1(n9880), .I2(n9879), .O(n9887) );
  NAND_GATE U10539 ( .I1(n9881), .I2(n1173), .O(n9885) );
  NAND3_GATE U10540 ( .I1(n9885), .I2(n9884), .I3(n9883), .O(n9886) );
  NAND_GATE U10541 ( .I1(n9887), .I2(n9886), .O(n10369) );
  INV_GATE U10542 ( .I1(n10369), .O(n10372) );
  OR_GATE U10543 ( .I1(n9888), .I2(n9890), .O(n9901) );
  NAND_GATE U10544 ( .I1(n9890), .I2(n9889), .O(n9895) );
  NAND_GATE U10545 ( .I1(n9891), .I2(n9895), .O(n9899) );
  NAND_GATE U10546 ( .I1(n9893), .I2(n9892), .O(n9894) );
  NAND_GATE U10547 ( .I1(n9895), .I2(n9894), .O(n9896) );
  NAND_GATE U10548 ( .I1(n9897), .I2(n9896), .O(n9898) );
  NAND_GATE U10549 ( .I1(n9899), .I2(n9898), .O(n9900) );
  NAND_GATE U10550 ( .I1(n9901), .I2(n9900), .O(n10385) );
  OR_GATE U10551 ( .I1(n9902), .I2(n9906), .O(n9905) );
  OR_GATE U10552 ( .I1(n9903), .I2(n9907), .O(n9904) );
  AND_GATE U10553 ( .I1(n9905), .I2(n9904), .O(n9912) );
  NAND_GATE U10554 ( .I1(n9906), .I2(n1241), .O(n9910) );
  NAND3_GATE U10555 ( .I1(n9910), .I2(n9909), .I3(n9908), .O(n9911) );
  NAND_GATE U10556 ( .I1(n9912), .I2(n9911), .O(n10394) );
  INV_GATE U10557 ( .I1(n10394), .O(n10397) );
  INV_GATE U10558 ( .I1(n9913), .O(n9914) );
  NAND_GATE U10559 ( .I1(n9918), .I2(n9914), .O(n9926) );
  NAND_GATE U10560 ( .I1(n9916), .I2(n9920), .O(n9924) );
  NAND_GATE U10561 ( .I1(n9918), .I2(n9917), .O(n9919) );
  NAND_GATE U10562 ( .I1(n9920), .I2(n9919), .O(n9921) );
  NAND_GATE U10563 ( .I1(n9922), .I2(n9921), .O(n9923) );
  NAND_GATE U10564 ( .I1(n9924), .I2(n9923), .O(n9925) );
  NAND_GATE U10565 ( .I1(n9926), .I2(n9925), .O(n10410) );
  NAND_GATE U10566 ( .I1(n1421), .I2(A[0]), .O(n9927) );
  NAND_GATE U10567 ( .I1(n14241), .I2(n9927), .O(n9928) );
  NAND_GATE U10568 ( .I1(n1422), .I2(n9928), .O(n9932) );
  NAND_GATE U10569 ( .I1(n1423), .I2(A[1]), .O(n9929) );
  NAND_GATE U10570 ( .I1(n724), .I2(n9929), .O(n9930) );
  NAND_GATE U10571 ( .I1(B[11]), .I2(n9930), .O(n9931) );
  NAND_GATE U10572 ( .I1(n9932), .I2(n9931), .O(n10422) );
  NAND_GATE U10573 ( .I1(B[10]), .I2(A[2]), .O(n10426) );
  NAND3_GATE U10574 ( .I1(B[10]), .I2(B[11]), .I3(n1254), .O(n10419) );
  NAND_GATE U10575 ( .I1(n10426), .I2(n10419), .O(n9933) );
  NAND_GATE U10576 ( .I1(n10422), .I2(n9933), .O(n9934) );
  INV_GATE U10577 ( .I1(n10426), .O(n10420) );
  INV_GATE U10578 ( .I1(n10419), .O(n10421) );
  NAND_GATE U10579 ( .I1(n10420), .I2(n10421), .O(n10417) );
  NAND_GATE U10580 ( .I1(n9934), .I2(n10417), .O(n10411) );
  NAND_GATE U10581 ( .I1(n10410), .I2(n10411), .O(n9936) );
  NAND_GATE U10582 ( .I1(B[10]), .I2(A[3]), .O(n10412) );
  INV_GATE U10583 ( .I1(n10412), .O(n9935) );
  NAND_GATE U10584 ( .I1(n10410), .I2(n9935), .O(n10407) );
  NAND_GATE U10585 ( .I1(n10411), .I2(n9935), .O(n10406) );
  NAND3_GATE U10586 ( .I1(n9936), .I2(n10407), .I3(n10406), .O(n10396) );
  INV_GATE U10587 ( .I1(n10396), .O(n10393) );
  NAND_GATE U10588 ( .I1(B[10]), .I2(A[4]), .O(n10401) );
  NAND_GATE U10589 ( .I1(n10393), .I2(n10401), .O(n9937) );
  NAND_GATE U10590 ( .I1(n10397), .I2(n9937), .O(n9938) );
  INV_GATE U10591 ( .I1(n10401), .O(n10395) );
  NAND_GATE U10592 ( .I1(n10396), .I2(n10395), .O(n10392) );
  NAND_GATE U10593 ( .I1(n9938), .I2(n10392), .O(n10386) );
  NAND_GATE U10594 ( .I1(n10385), .I2(n10386), .O(n9940) );
  NAND_GATE U10595 ( .I1(B[10]), .I2(A[5]), .O(n10387) );
  INV_GATE U10596 ( .I1(n10387), .O(n9939) );
  NAND_GATE U10597 ( .I1(n10385), .I2(n9939), .O(n10382) );
  NAND_GATE U10598 ( .I1(n10386), .I2(n9939), .O(n10381) );
  NAND3_GATE U10599 ( .I1(n9940), .I2(n10382), .I3(n10381), .O(n10371) );
  INV_GATE U10600 ( .I1(n10371), .O(n10368) );
  NAND_GATE U10601 ( .I1(B[10]), .I2(A[6]), .O(n10376) );
  NAND_GATE U10602 ( .I1(n10368), .I2(n10376), .O(n9941) );
  NAND_GATE U10603 ( .I1(n10372), .I2(n9941), .O(n9942) );
  INV_GATE U10604 ( .I1(n10376), .O(n10370) );
  NAND_GATE U10605 ( .I1(n10371), .I2(n10370), .O(n10367) );
  NAND_GATE U10606 ( .I1(n9942), .I2(n10367), .O(n10362) );
  NAND_GATE U10607 ( .I1(n10361), .I2(n10362), .O(n9944) );
  NAND_GATE U10608 ( .I1(B[10]), .I2(A[7]), .O(n10363) );
  INV_GATE U10609 ( .I1(n10363), .O(n9943) );
  NAND_GATE U10610 ( .I1(n10361), .I2(n9943), .O(n10358) );
  NAND_GATE U10611 ( .I1(n10362), .I2(n9943), .O(n10357) );
  NAND3_GATE U10612 ( .I1(n9944), .I2(n10358), .I3(n10357), .O(n10348) );
  NAND_GATE U10613 ( .I1(n10346), .I2(n10348), .O(n10343) );
  OR_GATE U10614 ( .I1(n9945), .I2(n9949), .O(n9948) );
  OR_GATE U10615 ( .I1(n9950), .I2(n9946), .O(n9947) );
  NAND_GATE U10616 ( .I1(n9949), .I2(n1059), .O(n9953) );
  NAND3_GATE U10617 ( .I1(n9953), .I2(n9952), .I3(n9951), .O(n9954) );
  INV_GATE U10618 ( .I1(n10344), .O(n10347) );
  INV_GATE U10619 ( .I1(n10348), .O(n10345) );
  NAND_GATE U10620 ( .I1(n10352), .I2(n10345), .O(n9955) );
  NAND_GATE U10621 ( .I1(n10347), .I2(n9955), .O(n9956) );
  NAND_GATE U10622 ( .I1(n10343), .I2(n9956), .O(n10458) );
  NAND_GATE U10623 ( .I1(n10457), .I2(n10458), .O(n9958) );
  NAND_GATE U10624 ( .I1(n9957), .I2(n10458), .O(n10453) );
  NAND3_GATE U10625 ( .I1(n10454), .I2(n9958), .I3(n10453), .O(n10334) );
  NAND_GATE U10626 ( .I1(n10332), .I2(n10334), .O(n10329) );
  OR_GATE U10627 ( .I1(n9959), .I2(n9963), .O(n9962) );
  OR_GATE U10628 ( .I1(n9964), .I2(n9960), .O(n9961) );
  NAND_GATE U10629 ( .I1(n9963), .I2(n1038), .O(n9967) );
  NAND3_GATE U10630 ( .I1(n9967), .I2(n9966), .I3(n9965), .O(n9968) );
  INV_GATE U10631 ( .I1(n10330), .O(n10333) );
  INV_GATE U10632 ( .I1(n10334), .O(n10331) );
  NAND_GATE U10633 ( .I1(n10338), .I2(n10331), .O(n9969) );
  NAND_GATE U10634 ( .I1(n10333), .I2(n9969), .O(n9970) );
  NAND_GATE U10635 ( .I1(n10329), .I2(n9970), .O(n10472) );
  NAND_GATE U10636 ( .I1(n10471), .I2(n10472), .O(n9972) );
  NAND_GATE U10637 ( .I1(n9971), .I2(n10472), .O(n10467) );
  NAND3_GATE U10638 ( .I1(n10468), .I2(n9972), .I3(n10467), .O(n10320) );
  NAND_GATE U10639 ( .I1(n10319), .I2(n10320), .O(n10316) );
  OR_GATE U10640 ( .I1(n9973), .I2(n9977), .O(n9976) );
  OR_GATE U10641 ( .I1(n9978), .I2(n9974), .O(n9975) );
  AND_GATE U10642 ( .I1(n9976), .I2(n9975), .O(n9983) );
  NAND_GATE U10643 ( .I1(n9977), .I2(n1300), .O(n9981) );
  NAND3_GATE U10644 ( .I1(n9981), .I2(n9980), .I3(n9979), .O(n9982) );
  INV_GATE U10645 ( .I1(n10320), .O(n10318) );
  NAND_GATE U10646 ( .I1(n10324), .I2(n10318), .O(n9984) );
  NAND_GATE U10647 ( .I1(n749), .I2(n9984), .O(n9985) );
  NAND_GATE U10648 ( .I1(n10316), .I2(n9985), .O(n10487) );
  NAND_GATE U10649 ( .I1(n10486), .I2(n10487), .O(n9987) );
  NAND_GATE U10650 ( .I1(n9986), .I2(n10487), .O(n10482) );
  NAND_GATE U10651 ( .I1(n10304), .I2(n10306), .O(n10303) );
  NAND_GATE U10652 ( .I1(n9989), .I2(n9988), .O(n9990) );
  NAND_GATE U10653 ( .I1(n9991), .I2(n9990), .O(n9992) );
  NAND_GATE U10654 ( .I1(n9993), .I2(n9992), .O(n9997) );
  OR_GATE U10655 ( .I1(n9997), .I2(n9994), .O(n10006) );
  NAND_GATE U10656 ( .I1(n9995), .I2(n9990), .O(n9996) );
  NAND_GATE U10657 ( .I1(n10003), .I2(n9996), .O(n10000) );
  INV_GATE U10658 ( .I1(n10003), .O(n9998) );
  NAND_GATE U10659 ( .I1(n9998), .I2(n9997), .O(n9999) );
  NAND3_GATE U10660 ( .I1(n10001), .I2(n10000), .I3(n9999), .O(n10005) );
  OR_GATE U10661 ( .I1(n10003), .I2(n10002), .O(n10004) );
  NAND3_GATE U10662 ( .I1(n10006), .I2(n10005), .I3(n10004), .O(n10307) );
  INV_GATE U10663 ( .I1(n10307), .O(n10305) );
  NAND_GATE U10664 ( .I1(n10311), .I2(n778), .O(n10007) );
  NAND_GATE U10665 ( .I1(n10305), .I2(n10007), .O(n10008) );
  NAND_GATE U10666 ( .I1(n10303), .I2(n10008), .O(n10502) );
  NAND_GATE U10667 ( .I1(n10497), .I2(n10502), .O(n10010) );
  NAND_GATE U10668 ( .I1(B[10]), .I2(A[15]), .O(n10498) );
  INV_GATE U10669 ( .I1(n10498), .O(n10009) );
  NAND_GATE U10670 ( .I1(n10502), .I2(n10009), .O(n10496) );
  NAND3_GATE U10671 ( .I1(n10501), .I2(n10010), .I3(n10496), .O(n10509) );
  NAND_GATE U10672 ( .I1(n10512), .I2(n10509), .O(n10516) );
  OR_GATE U10673 ( .I1(n10015), .I2(n10011), .O(n10014) );
  OR_GATE U10674 ( .I1(n10012), .I2(n10016), .O(n10013) );
  AND_GATE U10675 ( .I1(n10014), .I2(n10013), .O(n10021) );
  NAND_GATE U10676 ( .I1(n10016), .I2(n1048), .O(n10017) );
  NAND3_GATE U10677 ( .I1(n10019), .I2(n10018), .I3(n10017), .O(n10020) );
  NAND_GATE U10678 ( .I1(n10021), .I2(n10020), .O(n10517) );
  INV_GATE U10679 ( .I1(n10517), .O(n10508) );
  NAND_GATE U10680 ( .I1(n10507), .I2(n10510), .O(n10022) );
  NAND_GATE U10681 ( .I1(n10508), .I2(n10022), .O(n10023) );
  NAND_GATE U10682 ( .I1(n10516), .I2(n10023), .O(n10296) );
  NAND_GATE U10683 ( .I1(n10037), .I2(n10296), .O(n10293) );
  NAND_GATE U10684 ( .I1(n10028), .I2(n10035), .O(n10024) );
  NAND_GATE U10685 ( .I1(n10025), .I2(n10024), .O(n10033) );
  NAND_GATE U10686 ( .I1(n10027), .I2(n10026), .O(n10029) );
  NAND_GATE U10687 ( .I1(n10029), .I2(n10024), .O(n10030) );
  OR_GATE U10688 ( .I1(n10035), .I2(n10034), .O(n10036) );
  NAND_GATE U10689 ( .I1(n10296), .I2(n10297), .O(n10038) );
  NAND_GATE U10690 ( .I1(n10291), .I2(n10290), .O(n10039) );
  NAND_GATE U10691 ( .I1(n10286), .I2(n10039), .O(n10040) );
  NAND_GATE U10692 ( .I1(n10283), .I2(n10040), .O(n10274) );
  NAND_GATE U10693 ( .I1(n10054), .I2(n10274), .O(n10278) );
  NAND3_GATE U10694 ( .I1(n10043), .I2(n886), .I3(n10041), .O(n10048) );
  NAND_GATE U10695 ( .I1(n10042), .I2(n10050), .O(n10047) );
  NAND_GATE U10696 ( .I1(n10043), .I2(n886), .O(n10044) );
  NAND_GATE U10697 ( .I1(n10045), .I2(n10044), .O(n10046) );
  NAND3_GATE U10698 ( .I1(n10048), .I2(n10047), .I3(n10046), .O(n10053) );
  INV_GATE U10699 ( .I1(n10049), .O(n10051) );
  NAND_GATE U10700 ( .I1(n10051), .I2(n10050), .O(n10052) );
  NAND_GATE U10701 ( .I1(n10053), .I2(n10052), .O(n10279) );
  NAND_GATE U10702 ( .I1(n10274), .I2(n10279), .O(n10055) );
  NAND_GATE U10703 ( .I1(n10054), .I2(n10279), .O(n10273) );
  NAND3_GATE U10704 ( .I1(n10278), .I2(n10055), .I3(n10273), .O(n10532) );
  NAND_GATE U10705 ( .I1(n10534), .I2(n10531), .O(n10056) );
  NAND_GATE U10706 ( .I1(n10532), .I2(n10056), .O(n10057) );
  NAND_GATE U10707 ( .I1(n10529), .I2(n10057), .O(n10265) );
  INV_GATE U10708 ( .I1(n10063), .O(n10059) );
  NAND_GATE U10709 ( .I1(n10060), .I2(n10059), .O(n10066) );
  NAND3_GATE U10710 ( .I1(n10062), .I2(n10061), .I3(n10066), .O(n10071) );
  NAND_GATE U10711 ( .I1(n10064), .I2(n10063), .O(n10065) );
  NAND_GATE U10712 ( .I1(n10066), .I2(n10065), .O(n10069) );
  NAND_GATE U10713 ( .I1(n10070), .I2(n10069), .O(n10067) );
  NAND3_GATE U10714 ( .I1(n10068), .I2(n10071), .I3(n10067), .O(n10266) );
  NAND_GATE U10715 ( .I1(n10071), .I2(n10067), .O(n10268) );
  NAND_GATE U10716 ( .I1(n10265), .I2(n646), .O(n10072) );
  NAND3_GATE U10717 ( .I1(n10267), .I2(n10266), .I3(n10072), .O(n10259) );
  NAND_GATE U10718 ( .I1(n10604), .I2(n10257), .O(n10073) );
  NAND_GATE U10719 ( .I1(n10259), .I2(n10073), .O(n10074) );
  NAND_GATE U10720 ( .I1(n10075), .I2(n10074), .O(n10248) );
  NAND_GATE U10721 ( .I1(n10084), .I2(n10248), .O(n10252) );
  NAND_GATE U10722 ( .I1(n10077), .I2(n10080), .O(n10242) );
  NAND_GATE U10723 ( .I1(n718), .I2(n10078), .O(n10081) );
  NAND_GATE U10724 ( .I1(n10079), .I2(n979), .O(n10080) );
  NAND_GATE U10725 ( .I1(n10081), .I2(n10080), .O(n10244) );
  NAND_GATE U10726 ( .I1(n10245), .I2(n10244), .O(n10082) );
  NAND_GATE U10727 ( .I1(n10242), .I2(n10082), .O(n10083) );
  NAND_GATE U10728 ( .I1(n10243), .I2(n10083), .O(n10253) );
  NAND_GATE U10729 ( .I1(n10084), .I2(n10253), .O(n10254) );
  NAND_GATE U10730 ( .I1(n10248), .I2(n10253), .O(n10085) );
  NAND3_GATE U10731 ( .I1(n10252), .I2(n10254), .I3(n10085), .O(n10234) );
  NAND_GATE U10732 ( .I1(n10099), .I2(n10234), .O(n10240) );
  INV_GATE U10733 ( .I1(n10086), .O(n10087) );
  NAND_GATE U10734 ( .I1(n10087), .I2(n10090), .O(n10098) );
  INV_GATE U10735 ( .I1(n10090), .O(n10092) );
  NAND_GATE U10736 ( .I1(n10093), .I2(n10092), .O(n10088) );
  NAND_GATE U10737 ( .I1(n10089), .I2(n10088), .O(n10096) );
  NAND_GATE U10738 ( .I1(n654), .I2(n10090), .O(n10095) );
  NAND3_GATE U10739 ( .I1(n10093), .I2(n10092), .I3(n10091), .O(n10094) );
  NAND3_GATE U10740 ( .I1(n10096), .I2(n10095), .I3(n10094), .O(n10097) );
  NAND_GATE U10741 ( .I1(n10098), .I2(n10097), .O(n10235) );
  NAND_GATE U10742 ( .I1(n10099), .I2(n10235), .O(n10233) );
  NAND_GATE U10743 ( .I1(n10234), .I2(n10235), .O(n10100) );
  NAND3_GATE U10744 ( .I1(n10240), .I2(n10233), .I3(n10100), .O(n10222) );
  NAND_GATE U10745 ( .I1(n10227), .I2(n10222), .O(n10228) );
  NAND3_GATE U10746 ( .I1(n10101), .I2(n10102), .I3(n717), .O(n10219) );
  INV_GATE U10747 ( .I1(n10102), .O(n10103) );
  NAND_GATE U10748 ( .I1(n10101), .I2(n10105), .O(n10218) );
  NAND_GATE U10749 ( .I1(n717), .I2(n10102), .O(n10106) );
  NAND_GATE U10750 ( .I1(n10104), .I2(n10103), .O(n10105) );
  NAND_GATE U10751 ( .I1(n10106), .I2(n10105), .O(n10216) );
  NAND_GATE U10752 ( .I1(n10217), .I2(n10216), .O(n10107) );
  NAND_GATE U10753 ( .I1(n10218), .I2(n10107), .O(n10108) );
  NAND_GATE U10754 ( .I1(n10219), .I2(n10108), .O(n10229) );
  NAND_GATE U10755 ( .I1(n10227), .I2(n10229), .O(n10110) );
  NAND_GATE U10756 ( .I1(n10222), .I2(n10229), .O(n10109) );
  NAND3_GATE U10757 ( .I1(n10228), .I2(n10110), .I3(n10109), .O(n10205) );
  NAND_GATE U10758 ( .I1(n10210), .I2(n10205), .O(n10211) );
  NAND_GATE U10759 ( .I1(n10114), .I2(n991), .O(n10112) );
  NAND_GATE U10760 ( .I1(n571), .I2(n10112), .O(n10199) );
  NAND_GATE U10761 ( .I1(n10199), .I2(n10115), .O(n10116) );
  NAND_GATE U10762 ( .I1(n10200), .I2(n10116), .O(n10212) );
  NAND_GATE U10763 ( .I1(n10210), .I2(n10212), .O(n10118) );
  NAND_GATE U10764 ( .I1(n10205), .I2(n10212), .O(n10117) );
  NAND3_GATE U10765 ( .I1(n10211), .I2(n10118), .I3(n10117), .O(n10195) );
  NAND_GATE U10766 ( .I1(n10189), .I2(n10195), .O(n10190) );
  INV_GATE U10767 ( .I1(n10125), .O(n10120) );
  NAND3_GATE U10768 ( .I1(n10121), .I2(n10120), .I3(n10119), .O(n10123) );
  NAND3_GATE U10769 ( .I1(n10124), .I2(n10123), .I3(n10122), .O(n10127) );
  NAND_GATE U10770 ( .I1(n1284), .I2(n10125), .O(n10126) );
  NAND_GATE U10771 ( .I1(n10127), .I2(n10126), .O(n10194) );
  NAND_GATE U10772 ( .I1(n10189), .I2(n10194), .O(n10129) );
  NAND_GATE U10773 ( .I1(n10195), .I2(n10194), .O(n10128) );
  NAND3_GATE U10774 ( .I1(n10190), .I2(n10129), .I3(n10128), .O(n10183) );
  NAND_GATE U10775 ( .I1(n10183), .I2(n10182), .O(n10130) );
  NAND_GATE U10776 ( .I1(n10178), .I2(n10183), .O(n10179) );
  NAND3_GATE U10777 ( .I1(n10131), .I2(n10130), .I3(n10179), .O(n10172) );
  NAND_GATE U10778 ( .I1(n10166), .I2(n10172), .O(n10167) );
  INV_GATE U10779 ( .I1(n10132), .O(n10133) );
  NAND_GATE U10780 ( .I1(n10133), .I2(n10136), .O(n10142) );
  NAND_GATE U10781 ( .I1(n10135), .I2(n10134), .O(n10140) );
  NAND_GATE U10782 ( .I1(n10140), .I2(n10139), .O(n10141) );
  NAND_GATE U10783 ( .I1(n10142), .I2(n10141), .O(n10171) );
  NAND_GATE U10784 ( .I1(n10166), .I2(n10171), .O(n10144) );
  NAND_GATE U10785 ( .I1(n10172), .I2(n10171), .O(n10143) );
  NAND3_GATE U10786 ( .I1(n10167), .I2(n10144), .I3(n10143), .O(n10159) );
  NAND_GATE U10787 ( .I1(n10159), .I2(n10162), .O(n10146) );
  NAND_GATE U10788 ( .I1(n10145), .I2(n10159), .O(n10161) );
  AND3_GATE U10789 ( .I1(n10160), .I2(n10146), .I3(n10161), .O(n10153) );
  NAND_GATE U10790 ( .I1(n1420), .I2(A[31]), .O(n10152) );
  NAND_GATE U10791 ( .I1(n10153), .I2(n10152), .O(n10147) );
  NAND_GATE U10792 ( .I1(n10151), .I2(n10147), .O(n10155) );
  NAND_GATE U10793 ( .I1(n14818), .I2(n10155), .O(n10150) );
  NAND_GATE U10794 ( .I1(n10148), .I2(n830), .O(n10149) );
  NAND_GATE U10795 ( .I1(n10150), .I2(n10149), .O(\A1[40] ) );
  NAND_GATE U10796 ( .I1(n10155), .I2(n10154), .O(n10571) );
  NAND_GATE U10797 ( .I1(n950), .I2(n10162), .O(n10158) );
  NAND3_GATE U10798 ( .I1(n10158), .I2(n10157), .I3(n10156), .O(n10165) );
  OR_GATE U10799 ( .I1(n10160), .I2(n10159), .O(n10164) );
  OR_GATE U10800 ( .I1(n10162), .I2(n10161), .O(n10163) );
  NAND3_GATE U10801 ( .I1(n10165), .I2(n10164), .I3(n10163), .O(n10574) );
  INV_GATE U10802 ( .I1(n10172), .O(n10170) );
  NAND3_GATE U10803 ( .I1(n10170), .I2(n10166), .I3(n10171), .O(n10169) );
  OR_GATE U10804 ( .I1(n10171), .I2(n10167), .O(n10168) );
  AND_GATE U10805 ( .I1(n10169), .I2(n10168), .O(n10177) );
  NAND_GATE U10806 ( .I1(n10170), .I2(n10171), .O(n10174) );
  NAND3_GATE U10807 ( .I1(n10175), .I2(n10174), .I3(n10173), .O(n10176) );
  NAND_GATE U10808 ( .I1(n10177), .I2(n10176), .O(n10579) );
  NAND_GATE U10809 ( .I1(n1418), .I2(A[30]), .O(n10577) );
  INV_GATE U10810 ( .I1(n10577), .O(n10580) );
  NAND_GATE U10811 ( .I1(n719), .I2(n10580), .O(n10575) );
  NAND_GATE U10812 ( .I1(n1418), .I2(A[29]), .O(n10964) );
  INV_GATE U10813 ( .I1(n10964), .O(n10959) );
  NAND3_GATE U10814 ( .I1(n10178), .I2(n169), .I3(n10182), .O(n10181) );
  OR_GATE U10815 ( .I1(n10182), .I2(n10179), .O(n10180) );
  AND_GATE U10816 ( .I1(n10181), .I2(n10180), .O(n10188) );
  NAND_GATE U10817 ( .I1(n169), .I2(n10182), .O(n10185) );
  NAND3_GATE U10818 ( .I1(n10186), .I2(n10185), .I3(n10184), .O(n10187) );
  NAND_GATE U10819 ( .I1(n10188), .I2(n10187), .O(n10961) );
  INV_GATE U10820 ( .I1(n10961), .O(n10963) );
  NAND_GATE U10821 ( .I1(n1418), .I2(A[28]), .O(n10989) );
  INV_GATE U10822 ( .I1(n10989), .O(n10951) );
  INV_GATE U10823 ( .I1(n10195), .O(n10193) );
  NAND3_GATE U10824 ( .I1(n10189), .I2(n10193), .I3(n10194), .O(n10192) );
  OR_GATE U10825 ( .I1(n10194), .I2(n10190), .O(n10191) );
  AND_GATE U10826 ( .I1(n10192), .I2(n10191), .O(n10586) );
  NAND_GATE U10827 ( .I1(n10193), .I2(n10194), .O(n10198) );
  NAND3_GATE U10828 ( .I1(n10198), .I2(n10197), .I3(n10196), .O(n10587) );
  NAND_GATE U10829 ( .I1(n10586), .I2(n10587), .O(n10949) );
  NAND_GATE U10830 ( .I1(n10951), .I2(n10591), .O(n10565) );
  NAND_GATE U10831 ( .I1(n1418), .I2(A[27]), .O(n11009) );
  INV_GATE U10832 ( .I1(n11009), .O(n10597) );
  INV_GATE U10833 ( .I1(n10205), .O(n10209) );
  NAND_GATE U10834 ( .I1(n10203), .I2(n10202), .O(n10204) );
  NAND_GATE U10835 ( .I1(n10205), .I2(n10204), .O(n10206) );
  NAND3_GATE U10836 ( .I1(n10208), .I2(n10207), .I3(n10206), .O(n10215) );
  NAND3_GATE U10837 ( .I1(n10210), .I2(n10209), .I3(n10212), .O(n10214) );
  OR_GATE U10838 ( .I1(n10212), .I2(n10211), .O(n10213) );
  NAND3_GATE U10839 ( .I1(n10215), .I2(n10214), .I3(n10213), .O(n10595) );
  NAND_GATE U10840 ( .I1(n10597), .I2(n621), .O(n10562) );
  NAND_GATE U10841 ( .I1(n1418), .I2(A[26]), .O(n11022) );
  INV_GATE U10842 ( .I1(n11022), .O(n10935) );
  INV_GATE U10843 ( .I1(n10222), .O(n10226) );
  NAND3_GATE U10844 ( .I1(n10107), .I2(n10226), .I3(n10220), .O(n10225) );
  NAND_GATE U10845 ( .I1(n10220), .I2(n10107), .O(n10221) );
  NAND_GATE U10846 ( .I1(n10222), .I2(n10221), .O(n10224) );
  NAND3_GATE U10847 ( .I1(n10225), .I2(n10224), .I3(n10223), .O(n10232) );
  NAND3_GATE U10848 ( .I1(n10227), .I2(n10226), .I3(n10229), .O(n10231) );
  OR_GATE U10849 ( .I1(n10229), .I2(n10228), .O(n10230) );
  NAND3_GATE U10850 ( .I1(n10232), .I2(n10231), .I3(n10230), .O(n10937) );
  NAND_GATE U10851 ( .I1(n10935), .I2(n677), .O(n10559) );
  INV_GATE U10852 ( .I1(n10234), .O(n10236) );
  NAND_GATE U10853 ( .I1(n10234), .I2(n678), .O(n10238) );
  NAND_GATE U10854 ( .I1(n10236), .I2(n10235), .O(n10237) );
  NAND3_GATE U10855 ( .I1(n10239), .I2(n10238), .I3(n10237), .O(n10551) );
  INV_GATE U10856 ( .I1(n10240), .O(n10241) );
  NAND_GATE U10857 ( .I1(n10241), .I2(n678), .O(n10553) );
  INV_GATE U10858 ( .I1(n10248), .O(n10255) );
  NAND3_GATE U10859 ( .I1(n10246), .I2(n10082), .I3(n10255), .O(n10251) );
  NAND_GATE U10860 ( .I1(n10246), .I2(n10082), .O(n10247) );
  NAND_GATE U10861 ( .I1(n10248), .I2(n10247), .O(n10250) );
  NAND3_GATE U10862 ( .I1(n10251), .I2(n10250), .I3(n10249), .O(n10924) );
  NAND_GATE U10863 ( .I1(n1418), .I2(A[24]), .O(n11044) );
  INV_GATE U10864 ( .I1(n11044), .O(n10919) );
  NAND3_GATE U10865 ( .I1(n10924), .I2(n968), .I3(n10919), .O(n10920) );
  NAND_GATE U10866 ( .I1(n1418), .I2(A[23]), .O(n10611) );
  INV_GATE U10867 ( .I1(n10611), .O(n10614) );
  NAND_GATE U10868 ( .I1(n874), .I2(n10259), .O(n10256) );
  NAND_GATE U10869 ( .I1(n10256), .I2(n10258), .O(n10603) );
  NAND_GATE U10870 ( .I1(n10257), .I2(n6), .O(n10258) );
  NAND_GATE U10871 ( .I1(n10260), .I2(n10258), .O(n10605) );
  NAND_GATE U10872 ( .I1(n10607), .I2(n10605), .O(n10261) );
  NAND3_GATE U10873 ( .I1(n10260), .I2(n10259), .I3(n874), .O(n10606) );
  NAND_GATE U10874 ( .I1(n10261), .I2(n10606), .O(n10615) );
  NAND_GATE U10875 ( .I1(n1418), .I2(A[22]), .O(n11056) );
  INV_GATE U10876 ( .I1(n11056), .O(n10626) );
  NAND_GATE U10877 ( .I1(n10265), .I2(n10268), .O(n10263) );
  NAND_GATE U10878 ( .I1(n397), .I2(n646), .O(n10262) );
  NAND3_GATE U10879 ( .I1(n10264), .I2(n10263), .I3(n10262), .O(n10272) );
  OR_GATE U10880 ( .I1(n10266), .I2(n10265), .O(n10271) );
  INV_GATE U10881 ( .I1(n10267), .O(n10269) );
  NAND_GATE U10882 ( .I1(n10269), .I2(n10268), .O(n10270) );
  NAND3_GATE U10883 ( .I1(n10272), .I2(n10271), .I3(n10270), .O(n10622) );
  NAND_GATE U10884 ( .I1(n10626), .I2(n10624), .O(n10546) );
  NAND_GATE U10885 ( .I1(n1418), .I2(A[21]), .O(n10633) );
  INV_GATE U10886 ( .I1(n10633), .O(n10542) );
  NAND_GATE U10887 ( .I1(n1418), .I2(A[20]), .O(n10899) );
  OR_GATE U10888 ( .I1(n10273), .I2(n10274), .O(n10282) );
  NAND_GATE U10889 ( .I1(n1299), .I2(n10279), .O(n10275) );
  NAND3_GATE U10890 ( .I1(n10277), .I2(n10276), .I3(n10275), .O(n10281) );
  OR_GATE U10891 ( .I1(n10279), .I2(n10278), .O(n10280) );
  NAND3_GATE U10892 ( .I1(n10282), .I2(n10281), .I3(n10280), .O(n10898) );
  NAND_GATE U10893 ( .I1(n10291), .I2(n1393), .O(n10284) );
  NAND_GATE U10894 ( .I1(n10285), .I2(n10284), .O(n10289) );
  NAND_GATE U10895 ( .I1(n10287), .I2(n10286), .O(n10288) );
  NAND_GATE U10896 ( .I1(n10289), .I2(n10288), .O(n10637) );
  NAND_GATE U10897 ( .I1(n10640), .I2(n10637), .O(n10524) );
  NAND3_GATE U10898 ( .I1(n10291), .I2(n1393), .I3(n10290), .O(n10638) );
  NAND_GATE U10899 ( .I1(n1418), .I2(A[19]), .O(n10647) );
  INV_GATE U10900 ( .I1(n10647), .O(n10525) );
  NAND3_GATE U10901 ( .I1(n10524), .I2(n10638), .I3(n10525), .O(n10642) );
  OR_GATE U10902 ( .I1(n10292), .I2(n10296), .O(n10295) );
  OR_GATE U10903 ( .I1(n10297), .I2(n10293), .O(n10294) );
  AND_GATE U10904 ( .I1(n10295), .I2(n10294), .O(n10302) );
  NAND_GATE U10905 ( .I1(n1022), .I2(n10297), .O(n10298) );
  NAND3_GATE U10906 ( .I1(n10300), .I2(n10299), .I3(n10298), .O(n10301) );
  NAND_GATE U10907 ( .I1(n10302), .I2(n10301), .O(n10887) );
  NAND_GATE U10908 ( .I1(n1418), .I2(A[18]), .O(n11324) );
  INV_GATE U10909 ( .I1(n11324), .O(n10882) );
  NAND_GATE U10910 ( .I1(n10885), .I2(n10882), .O(n10883) );
  NAND_GATE U10911 ( .I1(n1418), .I2(A[17]), .O(n10876) );
  INV_GATE U10912 ( .I1(n10876), .O(n10520) );
  NAND_GATE U10913 ( .I1(n1418), .I2(A[16]), .O(n10861) );
  INV_GATE U10914 ( .I1(n10861), .O(n10856) );
  NAND_GATE U10915 ( .I1(n1418), .I2(A[15]), .O(n10848) );
  INV_GATE U10916 ( .I1(n10848), .O(n10494) );
  OR_GATE U10917 ( .I1(n10307), .I2(n10303), .O(n10315) );
  NAND_GATE U10918 ( .I1(n10304), .I2(n10308), .O(n10313) );
  NAND_GATE U10919 ( .I1(n778), .I2(n10307), .O(n10308) );
  NAND_GATE U10920 ( .I1(n10309), .I2(n10308), .O(n10310) );
  NAND_GATE U10921 ( .I1(n10311), .I2(n10310), .O(n10312) );
  NAND_GATE U10922 ( .I1(n10313), .I2(n10312), .O(n10314) );
  NAND_GATE U10923 ( .I1(n10315), .I2(n10314), .O(n10846) );
  NAND_GATE U10924 ( .I1(n1418), .I2(A[14]), .O(n10659) );
  INV_GATE U10925 ( .I1(n10659), .O(n10654) );
  NAND_GATE U10926 ( .I1(n1418), .I2(A[13]), .O(n10833) );
  INV_GATE U10927 ( .I1(n10833), .O(n10480) );
  OR_GATE U10928 ( .I1(n10317), .I2(n10316), .O(n10328) );
  NAND_GATE U10929 ( .I1(n10319), .I2(n10322), .O(n10326) );
  NAND_GATE U10930 ( .I1(n10320), .I2(n749), .O(n10321) );
  NAND_GATE U10931 ( .I1(n10322), .I2(n10321), .O(n10323) );
  NAND_GATE U10932 ( .I1(n10324), .I2(n10323), .O(n10325) );
  NAND_GATE U10933 ( .I1(n10326), .I2(n10325), .O(n10327) );
  NAND_GATE U10934 ( .I1(n10328), .I2(n10327), .O(n10831) );
  NAND_GATE U10935 ( .I1(n10480), .I2(n10831), .O(n10828) );
  NAND_GATE U10936 ( .I1(n1418), .I2(A[12]), .O(n10671) );
  INV_GATE U10937 ( .I1(n10671), .O(n10666) );
  NAND_GATE U10938 ( .I1(n1418), .I2(A[11]), .O(n10819) );
  INV_GATE U10939 ( .I1(n10819), .O(n10465) );
  OR_GATE U10940 ( .I1(n10330), .I2(n10329), .O(n10342) );
  NAND_GATE U10941 ( .I1(n10331), .I2(n10330), .O(n10336) );
  NAND_GATE U10942 ( .I1(n10332), .I2(n10336), .O(n10340) );
  NAND_GATE U10943 ( .I1(n10334), .I2(n10333), .O(n10335) );
  NAND_GATE U10944 ( .I1(n10336), .I2(n10335), .O(n10337) );
  NAND_GATE U10945 ( .I1(n10338), .I2(n10337), .O(n10339) );
  NAND_GATE U10946 ( .I1(n10340), .I2(n10339), .O(n10341) );
  NAND_GATE U10947 ( .I1(n10342), .I2(n10341), .O(n10817) );
  NAND_GATE U10948 ( .I1(n10465), .I2(n10817), .O(n10814) );
  NAND_GATE U10949 ( .I1(n1418), .I2(A[10]), .O(n10683) );
  INV_GATE U10950 ( .I1(n10683), .O(n10677) );
  OR_GATE U10951 ( .I1(n10344), .I2(n10343), .O(n10356) );
  NAND_GATE U10952 ( .I1(n10345), .I2(n10344), .O(n10350) );
  NAND_GATE U10953 ( .I1(n10346), .I2(n10350), .O(n10354) );
  NAND_GATE U10954 ( .I1(n10348), .I2(n10347), .O(n10349) );
  NAND_GATE U10955 ( .I1(n10350), .I2(n10349), .O(n10351) );
  NAND_GATE U10956 ( .I1(n10352), .I2(n10351), .O(n10353) );
  NAND_GATE U10957 ( .I1(n10354), .I2(n10353), .O(n10355) );
  NAND_GATE U10958 ( .I1(n10356), .I2(n10355), .O(n10692) );
  OR_GATE U10959 ( .I1(n10357), .I2(n10361), .O(n10360) );
  OR_GATE U10960 ( .I1(n10358), .I2(n10362), .O(n10359) );
  NAND_GATE U10961 ( .I1(n10361), .I2(n1064), .O(n10365) );
  NAND3_GATE U10962 ( .I1(n10365), .I2(n10364), .I3(n10363), .O(n10366) );
  INV_GATE U10963 ( .I1(n10700), .O(n10703) );
  OR_GATE U10964 ( .I1(n10367), .I2(n10369), .O(n10380) );
  NAND_GATE U10965 ( .I1(n10369), .I2(n10368), .O(n10374) );
  NAND_GATE U10966 ( .I1(n10370), .I2(n10374), .O(n10378) );
  NAND_GATE U10967 ( .I1(n10372), .I2(n10371), .O(n10373) );
  NAND_GATE U10968 ( .I1(n10374), .I2(n10373), .O(n10375) );
  NAND_GATE U10969 ( .I1(n10376), .I2(n10375), .O(n10377) );
  NAND_GATE U10970 ( .I1(n10378), .I2(n10377), .O(n10379) );
  NAND_GATE U10971 ( .I1(n10380), .I2(n10379), .O(n10716) );
  OR_GATE U10972 ( .I1(n10381), .I2(n10385), .O(n10384) );
  OR_GATE U10973 ( .I1(n10382), .I2(n10386), .O(n10383) );
  AND_GATE U10974 ( .I1(n10384), .I2(n10383), .O(n10391) );
  NAND_GATE U10975 ( .I1(n10385), .I2(n1176), .O(n10389) );
  NAND3_GATE U10976 ( .I1(n10389), .I2(n10388), .I3(n10387), .O(n10390) );
  NAND_GATE U10977 ( .I1(n10391), .I2(n10390), .O(n10725) );
  INV_GATE U10978 ( .I1(n10725), .O(n10728) );
  OR_GATE U10979 ( .I1(n10392), .I2(n10394), .O(n10405) );
  NAND_GATE U10980 ( .I1(n10394), .I2(n10393), .O(n10399) );
  NAND_GATE U10981 ( .I1(n10395), .I2(n10399), .O(n10403) );
  NAND_GATE U10982 ( .I1(n10397), .I2(n10396), .O(n10398) );
  NAND_GATE U10983 ( .I1(n10399), .I2(n10398), .O(n10400) );
  NAND_GATE U10984 ( .I1(n10401), .I2(n10400), .O(n10402) );
  NAND_GATE U10985 ( .I1(n10403), .I2(n10402), .O(n10404) );
  NAND_GATE U10986 ( .I1(n10405), .I2(n10404), .O(n10741) );
  OR_GATE U10987 ( .I1(n10406), .I2(n10410), .O(n10409) );
  OR_GATE U10988 ( .I1(n10407), .I2(n10411), .O(n10408) );
  AND_GATE U10989 ( .I1(n10409), .I2(n10408), .O(n10416) );
  NAND_GATE U10990 ( .I1(n10410), .I2(n1242), .O(n10414) );
  NAND3_GATE U10991 ( .I1(n10414), .I2(n10413), .I3(n10412), .O(n10415) );
  NAND_GATE U10992 ( .I1(n10416), .I2(n10415), .O(n10750) );
  INV_GATE U10993 ( .I1(n10750), .O(n10753) );
  INV_GATE U10994 ( .I1(n10417), .O(n10418) );
  NAND_GATE U10995 ( .I1(n10422), .I2(n10418), .O(n10430) );
  NAND_GATE U10996 ( .I1(n10420), .I2(n10424), .O(n10428) );
  NAND_GATE U10997 ( .I1(n10422), .I2(n10421), .O(n10423) );
  NAND_GATE U10998 ( .I1(n10424), .I2(n10423), .O(n10425) );
  NAND_GATE U10999 ( .I1(n10426), .I2(n10425), .O(n10427) );
  NAND_GATE U11000 ( .I1(n10428), .I2(n10427), .O(n10429) );
  NAND_GATE U11001 ( .I1(n10430), .I2(n10429), .O(n10766) );
  NAND_GATE U11002 ( .I1(n1420), .I2(A[0]), .O(n10431) );
  NAND_GATE U11003 ( .I1(n14241), .I2(n10431), .O(n10432) );
  NAND_GATE U11004 ( .I1(B[11]), .I2(n10432), .O(n10436) );
  NAND_GATE U11005 ( .I1(n1421), .I2(A[1]), .O(n10433) );
  NAND_GATE U11006 ( .I1(n724), .I2(n10433), .O(n10434) );
  NAND_GATE U11007 ( .I1(B[10]), .I2(n10434), .O(n10435) );
  NAND_GATE U11008 ( .I1(n10436), .I2(n10435), .O(n10778) );
  NAND_GATE U11009 ( .I1(n1418), .I2(A[2]), .O(n10782) );
  NAND3_GATE U11010 ( .I1(n1418), .I2(B[10]), .I3(n1254), .O(n10775) );
  NAND_GATE U11011 ( .I1(n10782), .I2(n10775), .O(n10437) );
  NAND_GATE U11012 ( .I1(n10778), .I2(n10437), .O(n10438) );
  INV_GATE U11013 ( .I1(n10782), .O(n10776) );
  INV_GATE U11014 ( .I1(n10775), .O(n10777) );
  NAND_GATE U11015 ( .I1(n10776), .I2(n10777), .O(n10773) );
  NAND_GATE U11016 ( .I1(n10438), .I2(n10773), .O(n10767) );
  NAND_GATE U11017 ( .I1(n10766), .I2(n10767), .O(n10440) );
  NAND_GATE U11018 ( .I1(n1418), .I2(A[3]), .O(n10768) );
  INV_GATE U11019 ( .I1(n10768), .O(n10439) );
  NAND_GATE U11020 ( .I1(n10766), .I2(n10439), .O(n10763) );
  NAND_GATE U11021 ( .I1(n10767), .I2(n10439), .O(n10762) );
  NAND3_GATE U11022 ( .I1(n10440), .I2(n10763), .I3(n10762), .O(n10752) );
  INV_GATE U11023 ( .I1(n10752), .O(n10749) );
  NAND_GATE U11024 ( .I1(n1418), .I2(A[4]), .O(n10757) );
  NAND_GATE U11025 ( .I1(n10749), .I2(n10757), .O(n10441) );
  NAND_GATE U11026 ( .I1(n10753), .I2(n10441), .O(n10442) );
  INV_GATE U11027 ( .I1(n10757), .O(n10751) );
  NAND_GATE U11028 ( .I1(n10752), .I2(n10751), .O(n10748) );
  NAND_GATE U11029 ( .I1(n10442), .I2(n10748), .O(n10742) );
  NAND_GATE U11030 ( .I1(n10741), .I2(n10742), .O(n10444) );
  NAND_GATE U11031 ( .I1(n1418), .I2(A[5]), .O(n10743) );
  INV_GATE U11032 ( .I1(n10743), .O(n10443) );
  NAND_GATE U11033 ( .I1(n10741), .I2(n10443), .O(n10738) );
  NAND_GATE U11034 ( .I1(n10742), .I2(n10443), .O(n10737) );
  NAND3_GATE U11035 ( .I1(n10444), .I2(n10738), .I3(n10737), .O(n10727) );
  INV_GATE U11036 ( .I1(n10727), .O(n10724) );
  NAND_GATE U11037 ( .I1(n1418), .I2(A[6]), .O(n10732) );
  NAND_GATE U11038 ( .I1(n10724), .I2(n10732), .O(n10445) );
  NAND_GATE U11039 ( .I1(n10728), .I2(n10445), .O(n10446) );
  INV_GATE U11040 ( .I1(n10732), .O(n10726) );
  NAND_GATE U11041 ( .I1(n10727), .I2(n10726), .O(n10723) );
  NAND_GATE U11042 ( .I1(n10446), .I2(n10723), .O(n10717) );
  NAND_GATE U11043 ( .I1(n10716), .I2(n10717), .O(n10448) );
  NAND_GATE U11044 ( .I1(n1418), .I2(A[7]), .O(n10718) );
  INV_GATE U11045 ( .I1(n10718), .O(n10447) );
  NAND_GATE U11046 ( .I1(n10716), .I2(n10447), .O(n10713) );
  NAND_GATE U11047 ( .I1(n10717), .I2(n10447), .O(n10712) );
  NAND3_GATE U11048 ( .I1(n10448), .I2(n10713), .I3(n10712), .O(n10702) );
  INV_GATE U11049 ( .I1(n10702), .O(n10699) );
  NAND_GATE U11050 ( .I1(n1418), .I2(A[8]), .O(n10707) );
  NAND_GATE U11051 ( .I1(n10699), .I2(n10707), .O(n10449) );
  NAND_GATE U11052 ( .I1(n10703), .I2(n10449), .O(n10450) );
  INV_GATE U11053 ( .I1(n10707), .O(n10701) );
  NAND_GATE U11054 ( .I1(n10702), .I2(n10701), .O(n10698) );
  NAND_GATE U11055 ( .I1(n10450), .I2(n10698), .O(n10693) );
  NAND_GATE U11056 ( .I1(n10692), .I2(n10693), .O(n10452) );
  NAND_GATE U11057 ( .I1(n1418), .I2(A[9]), .O(n10694) );
  INV_GATE U11058 ( .I1(n10694), .O(n10451) );
  NAND_GATE U11059 ( .I1(n10692), .I2(n10451), .O(n10689) );
  NAND_GATE U11060 ( .I1(n10693), .I2(n10451), .O(n10688) );
  NAND3_GATE U11061 ( .I1(n10452), .I2(n10689), .I3(n10688), .O(n10679) );
  NAND_GATE U11062 ( .I1(n10677), .I2(n10679), .O(n10674) );
  OR_GATE U11063 ( .I1(n10453), .I2(n10457), .O(n10456) );
  OR_GATE U11064 ( .I1(n10458), .I2(n10454), .O(n10455) );
  NAND_GATE U11065 ( .I1(n10457), .I2(n1051), .O(n10461) );
  NAND3_GATE U11066 ( .I1(n10461), .I2(n10460), .I3(n10459), .O(n10462) );
  INV_GATE U11067 ( .I1(n10675), .O(n10678) );
  INV_GATE U11068 ( .I1(n10679), .O(n10676) );
  NAND_GATE U11069 ( .I1(n10683), .I2(n10676), .O(n10463) );
  NAND_GATE U11070 ( .I1(n10678), .I2(n10463), .O(n10464) );
  NAND_GATE U11071 ( .I1(n10674), .I2(n10464), .O(n10818) );
  NAND_GATE U11072 ( .I1(n10817), .I2(n10818), .O(n10466) );
  NAND_GATE U11073 ( .I1(n10465), .I2(n10818), .O(n10813) );
  NAND3_GATE U11074 ( .I1(n10814), .I2(n10466), .I3(n10813), .O(n10667) );
  NAND_GATE U11075 ( .I1(n10666), .I2(n10667), .O(n10663) );
  OR_GATE U11076 ( .I1(n10467), .I2(n10471), .O(n10470) );
  OR_GATE U11077 ( .I1(n10472), .I2(n10468), .O(n10469) );
  AND_GATE U11078 ( .I1(n10470), .I2(n10469), .O(n10477) );
  NAND_GATE U11079 ( .I1(n10471), .I2(n1008), .O(n10475) );
  NAND3_GATE U11080 ( .I1(n10475), .I2(n10474), .I3(n10473), .O(n10476) );
  NAND_GATE U11081 ( .I1(n10477), .I2(n10476), .O(n10664) );
  INV_GATE U11082 ( .I1(n10667), .O(n10665) );
  NAND_GATE U11083 ( .I1(n10671), .I2(n10665), .O(n10478) );
  NAND_GATE U11084 ( .I1(n656), .I2(n10478), .O(n10479) );
  NAND_GATE U11085 ( .I1(n10663), .I2(n10479), .O(n10832) );
  NAND_GATE U11086 ( .I1(n10831), .I2(n10832), .O(n10481) );
  NAND_GATE U11087 ( .I1(n10480), .I2(n10832), .O(n10827) );
  NAND3_GATE U11088 ( .I1(n10828), .I2(n10481), .I3(n10827), .O(n10655) );
  NAND_GATE U11089 ( .I1(n10654), .I2(n10655), .O(n10652) );
  OR_GATE U11090 ( .I1(n10482), .I2(n10486), .O(n10485) );
  OR_GATE U11091 ( .I1(n10487), .I2(n10483), .O(n10484) );
  NAND_GATE U11092 ( .I1(n10486), .I2(n1000), .O(n10490) );
  NAND3_GATE U11093 ( .I1(n10490), .I2(n10489), .I3(n10488), .O(n10491) );
  INV_GATE U11094 ( .I1(n10655), .O(n10653) );
  NAND_GATE U11095 ( .I1(n10659), .I2(n10653), .O(n10492) );
  NAND_GATE U11096 ( .I1(n779), .I2(n10492), .O(n10493) );
  NAND_GATE U11097 ( .I1(n10652), .I2(n10493), .O(n10847) );
  NAND_GATE U11098 ( .I1(n10846), .I2(n10847), .O(n10495) );
  NAND_GATE U11099 ( .I1(n10494), .I2(n10847), .O(n10842) );
  NAND3_GATE U11100 ( .I1(n10843), .I2(n10495), .I3(n10842), .O(n10857) );
  NAND_GATE U11101 ( .I1(n10856), .I2(n10857), .O(n10855) );
  OR_GATE U11102 ( .I1(n10496), .I2(n10497), .O(n10505) );
  NAND_GATE U11103 ( .I1(n10497), .I2(n1026), .O(n10500) );
  NAND3_GATE U11104 ( .I1(n10500), .I2(n10499), .I3(n10498), .O(n10504) );
  OR_GATE U11105 ( .I1(n10502), .I2(n10501), .O(n10503) );
  NAND3_GATE U11106 ( .I1(n10505), .I2(n10504), .I3(n10503), .O(n10858) );
  INV_GATE U11107 ( .I1(n10857), .O(n10859) );
  NAND_GATE U11108 ( .I1(n10855), .I2(n10506), .O(n10872) );
  NAND3_GATE U11109 ( .I1(n10517), .I2(n10507), .I3(n10510), .O(n10515) );
  NAND_GATE U11110 ( .I1(n10509), .I2(n10508), .O(n10514) );
  NAND_GATE U11111 ( .I1(n10510), .I2(n10517), .O(n10511) );
  NAND_GATE U11112 ( .I1(n10512), .I2(n10511), .O(n10513) );
  NAND3_GATE U11113 ( .I1(n10515), .I2(n10514), .I3(n10513), .O(n10519) );
  OR_GATE U11114 ( .I1(n10517), .I2(n10516), .O(n10518) );
  NAND_GATE U11115 ( .I1(n10519), .I2(n10518), .O(n10873) );
  NAND_GATE U11116 ( .I1(n10872), .I2(n10873), .O(n10521) );
  NAND_GATE U11117 ( .I1(n10520), .I2(n10873), .O(n10868) );
  NAND3_GATE U11118 ( .I1(n10869), .I2(n10521), .I3(n10868), .O(n10884) );
  NAND_GATE U11119 ( .I1(n10887), .I2(n11324), .O(n10522) );
  NAND_GATE U11120 ( .I1(n10884), .I2(n10522), .O(n10523) );
  NAND_GATE U11121 ( .I1(n10883), .I2(n10523), .O(n10646) );
  NAND3_GATE U11122 ( .I1(n10646), .I2(n10524), .I3(n10638), .O(n10526) );
  NAND_GATE U11123 ( .I1(n10525), .I2(n10646), .O(n10641) );
  NAND3_GATE U11124 ( .I1(n10642), .I2(n10526), .I3(n10641), .O(n10903) );
  NAND_GATE U11125 ( .I1(n10899), .I2(n10898), .O(n10527) );
  NAND_GATE U11126 ( .I1(n10903), .I2(n10527), .O(n10528) );
  NAND_GATE U11127 ( .I1(n10902), .I2(n10528), .O(n10632) );
  NAND_GATE U11128 ( .I1(n10542), .I2(n10632), .O(n10628) );
  INV_GATE U11129 ( .I1(n10529), .O(n10530) );
  NAND_GATE U11130 ( .I1(n10530), .I2(n10532), .O(n10541) );
  INV_GATE U11131 ( .I1(n10532), .O(n10533) );
  NAND3_GATE U11132 ( .I1(n10534), .I2(n10533), .I3(n10531), .O(n10539) );
  NAND_GATE U11133 ( .I1(n393), .I2(n10532), .O(n10538) );
  NAND_GATE U11134 ( .I1(n10534), .I2(n10533), .O(n10535) );
  NAND_GATE U11135 ( .I1(n10536), .I2(n10535), .O(n10537) );
  NAND3_GATE U11136 ( .I1(n10539), .I2(n10538), .I3(n10537), .O(n10540) );
  NAND_GATE U11137 ( .I1(n10541), .I2(n10540), .O(n10631) );
  NAND_GATE U11138 ( .I1(n10632), .I2(n10631), .O(n10543) );
  NAND_GATE U11139 ( .I1(n10542), .I2(n10631), .O(n10627) );
  NAND3_GATE U11140 ( .I1(n10628), .I2(n10543), .I3(n10627), .O(n10625) );
  NAND_GATE U11141 ( .I1(n11056), .I2(n10622), .O(n10544) );
  NAND_GATE U11142 ( .I1(n10625), .I2(n10544), .O(n10545) );
  NAND_GATE U11143 ( .I1(n10546), .I2(n10545), .O(n10610) );
  NAND_GATE U11144 ( .I1(n10615), .I2(n10610), .O(n10547) );
  NAND_GATE U11145 ( .I1(n10614), .I2(n10610), .O(n10616) );
  NAND3_GATE U11146 ( .I1(n10548), .I2(n10547), .I3(n10616), .O(n10926) );
  NAND_GATE U11147 ( .I1(n10919), .I2(n10926), .O(n10550) );
  NAND4_GATE U11148 ( .I1(n10925), .I2(n10923), .I3(n10926), .I4(n10924), .O(
        n10549) );
  NAND3_GATE U11149 ( .I1(n10920), .I2(n10550), .I3(n10549), .O(n10600) );
  NAND4_GATE U11150 ( .I1(n10552), .I2(n10551), .I3(n10553), .I4(n10600), .O(
        n10556) );
  NAND_GATE U11151 ( .I1(n1418), .I2(A[25]), .O(n11385) );
  NAND_GATE U11152 ( .I1(n532), .I2(n10600), .O(n10555) );
  NAND3_GATE U11153 ( .I1(n10553), .I2(n10552), .I3(n10551), .O(n10602) );
  NAND_GATE U11154 ( .I1(n681), .I2(n532), .O(n10554) );
  NAND3_GATE U11155 ( .I1(n10556), .I2(n10555), .I3(n10554), .O(n10938) );
  NAND_GATE U11156 ( .I1(n11022), .I2(n10937), .O(n10557) );
  NAND_GATE U11157 ( .I1(n10938), .I2(n10557), .O(n10558) );
  NAND_GATE U11158 ( .I1(n10559), .I2(n10558), .O(n10598) );
  NAND_GATE U11159 ( .I1(n11009), .I2(n10595), .O(n10560) );
  NAND_GATE U11160 ( .I1(n10598), .I2(n10560), .O(n10561) );
  NAND_GATE U11161 ( .I1(n10562), .I2(n10561), .O(n10592) );
  NAND_GATE U11162 ( .I1(n10989), .I2(n10949), .O(n10563) );
  NAND_GATE U11163 ( .I1(n10592), .I2(n10563), .O(n10564) );
  NAND_GATE U11164 ( .I1(n10565), .I2(n10564), .O(n10962) );
  NAND_GATE U11165 ( .I1(n10964), .I2(n10961), .O(n10566) );
  NAND_GATE U11166 ( .I1(n10962), .I2(n10566), .O(n10567) );
  NAND_GATE U11167 ( .I1(n10579), .I2(n10577), .O(n10568) );
  NAND_GATE U11168 ( .I1(n10578), .I2(n10568), .O(n10570) );
  NAND_GATE U11169 ( .I1(n1419), .I2(A[31]), .O(n10569) );
  NAND_GATE U11170 ( .I1(n10571), .I2(n1323), .O(n10572) );
  NAND_GATE U11171 ( .I1(n10573), .I2(n10572), .O(\A1[39] ) );
  INV_GATE U11172 ( .I1(n10575), .O(n10576) );
  NAND_GATE U11173 ( .I1(n10576), .I2(n10578), .O(n10585) );
  NAND3_GATE U11174 ( .I1(n10577), .I2(n926), .I3(n10579), .O(n10583) );
  NAND_GATE U11175 ( .I1(n719), .I2(n10578), .O(n10582) );
  NAND3_GATE U11176 ( .I1(n10583), .I2(n10582), .I3(n10581), .O(n10584) );
  NAND_GATE U11177 ( .I1(n10585), .I2(n10584), .O(n10973) );
  NAND_GATE U11178 ( .I1(n1417), .I2(A[31]), .O(n10971) );
  NAND3_GATE U11179 ( .I1(n10592), .I2(n10591), .I3(n10951), .O(n10996) );
  NAND_GATE U11180 ( .I1(n10951), .I2(n10592), .O(n10589) );
  NAND3_GATE U11181 ( .I1(n10587), .I2(n10586), .I3(n10951), .O(n10588) );
  NAND_GATE U11182 ( .I1(n10589), .I2(n10588), .O(n10590) );
  NAND_GATE U11183 ( .I1(n10996), .I2(n10590), .O(n10998) );
  NAND_GATE U11184 ( .I1(n10591), .I2(n10592), .O(n10593) );
  INV_GATE U11185 ( .I1(n10592), .O(n10948) );
  NAND_GATE U11186 ( .I1(n10593), .I2(n10950), .O(n10988) );
  NAND_GATE U11187 ( .I1(n1415), .I2(A[29]), .O(n10991) );
  INV_GATE U11188 ( .I1(n10991), .O(n10999) );
  NAND3_GATE U11189 ( .I1(n10998), .I2(n10992), .I3(n10999), .O(n10955) );
  NAND_GATE U11190 ( .I1(n10594), .I2(n10596), .O(n11008) );
  NAND_GATE U11191 ( .I1(n11009), .I2(n11008), .O(n10945) );
  NAND_GATE U11192 ( .I1(n10595), .I2(n569), .O(n10596) );
  NAND3_GATE U11193 ( .I1(n10598), .I2(n621), .I3(n10597), .O(n11011) );
  NAND_GATE U11194 ( .I1(n1271), .I2(n11011), .O(n10944) );
  NAND_GATE U11195 ( .I1(n1415), .I2(A[28]), .O(n11005) );
  INV_GATE U11196 ( .I1(n11005), .O(n11013) );
  NAND3_GATE U11197 ( .I1(n10945), .I2(n10944), .I3(n11013), .O(n10947) );
  NAND_GATE U11198 ( .I1(n1415), .I2(A[27]), .O(n11029) );
  INV_GATE U11199 ( .I1(n11029), .O(n11033) );
  NAND_GATE U11200 ( .I1(n1415), .I2(A[26]), .O(n11397) );
  INV_GATE U11201 ( .I1(n11397), .O(n11390) );
  INV_GATE U11202 ( .I1(n10600), .O(n10601) );
  NAND_GATE U11203 ( .I1(n10602), .I2(n10601), .O(n10599) );
  NAND_GATE U11204 ( .I1(n532), .I2(n10599), .O(n11387) );
  NAND3_GATE U11205 ( .I1(n532), .I2(n10600), .I3(n681), .O(n11384) );
  NAND3_GATE U11206 ( .I1(n11390), .I2(n11392), .I3(n11386), .O(n10934) );
  NAND_GATE U11207 ( .I1(n1415), .I2(A[25]), .O(n11049) );
  INV_GATE U11208 ( .I1(n11049), .O(n10921) );
  NAND_GATE U11209 ( .I1(n1415), .I2(A[24]), .O(n11374) );
  INV_GATE U11210 ( .I1(n11374), .O(n11371) );
  NAND_GATE U11211 ( .I1(n10604), .I2(n10603), .O(n10607) );
  NAND3_GATE U11212 ( .I1(n10607), .I2(n391), .I3(n10608), .O(n10613) );
  NAND_GATE U11213 ( .I1(n10608), .I2(n10607), .O(n10609) );
  NAND_GATE U11214 ( .I1(n10610), .I2(n10609), .O(n10612) );
  NAND3_GATE U11215 ( .I1(n10613), .I2(n10612), .I3(n10611), .O(n10619) );
  NAND3_GATE U11216 ( .I1(n391), .I2(n10614), .I3(n10615), .O(n10618) );
  OR_GATE U11217 ( .I1(n10616), .I2(n10615), .O(n10617) );
  NAND3_GATE U11218 ( .I1(n10619), .I2(n10618), .I3(n10617), .O(n11375) );
  NAND_GATE U11219 ( .I1(n11371), .I2(n392), .O(n11372) );
  NAND_GATE U11220 ( .I1(n1415), .I2(A[23]), .O(n11060) );
  INV_GATE U11221 ( .I1(n11060), .O(n10909) );
  NAND_GATE U11222 ( .I1(n10624), .I2(n10625), .O(n10620) );
  NAND_GATE U11223 ( .I1(n10623), .I2(n10620), .O(n11055) );
  NAND_GATE U11224 ( .I1(n10622), .I2(n10621), .O(n10623) );
  NAND_GATE U11225 ( .I1(n10626), .I2(n10623), .O(n10910) );
  NAND3_GATE U11226 ( .I1(n10626), .I2(n10625), .I3(n10624), .O(n10912) );
  NAND3_GATE U11227 ( .I1(n10909), .I2(n11057), .I3(n11058), .O(n11065) );
  NAND_GATE U11228 ( .I1(n1415), .I2(A[22]), .O(n11355) );
  OR_GATE U11229 ( .I1(n10627), .I2(n10632), .O(n10630) );
  OR_GATE U11230 ( .I1(n10631), .I2(n10628), .O(n10629) );
  NAND_GATE U11231 ( .I1(n1047), .I2(n10631), .O(n10635) );
  NAND3_GATE U11232 ( .I1(n10635), .I2(n10634), .I3(n10633), .O(n10636) );
  INV_GATE U11233 ( .I1(n11357), .O(n11358) );
  NAND_GATE U11234 ( .I1(n10640), .I2(n10639), .O(n10645) );
  OR_GATE U11235 ( .I1(n10645), .I2(n10641), .O(n10644) );
  OR_GATE U11236 ( .I1(n10646), .I2(n10642), .O(n10643) );
  AND_GATE U11237 ( .I1(n10644), .I2(n10643), .O(n10651) );
  NAND_GATE U11238 ( .I1(n695), .I2(n10645), .O(n10649) );
  NAND3_GATE U11239 ( .I1(n10649), .I2(n10648), .I3(n10647), .O(n10650) );
  NAND_GATE U11240 ( .I1(n10651), .I2(n10650), .O(n11342) );
  NAND_GATE U11241 ( .I1(n1415), .I2(A[20]), .O(n11343) );
  INV_GATE U11242 ( .I1(n11343), .O(n11340) );
  NAND_GATE U11243 ( .I1(n638), .I2(n11340), .O(n11346) );
  NAND_GATE U11244 ( .I1(n1416), .I2(A[19]), .O(n11330) );
  INV_GATE U11245 ( .I1(n11330), .O(n10892) );
  NAND_GATE U11246 ( .I1(n1416), .I2(A[17]), .O(n11086) );
  INV_GATE U11247 ( .I1(n11086), .O(n10866) );
  NAND_GATE U11248 ( .I1(n1416), .I2(A[16]), .O(n11303) );
  INV_GATE U11249 ( .I1(n11303), .O(n11296) );
  NAND_GATE U11250 ( .I1(n1416), .I2(A[15]), .O(n11289) );
  INV_GATE U11251 ( .I1(n11289), .O(n10840) );
  OR_GATE U11252 ( .I1(n26), .I2(n10652), .O(n10662) );
  NAND_GATE U11253 ( .I1(n10654), .I2(n10657), .O(n10661) );
  NAND_GATE U11254 ( .I1(n10655), .I2(n779), .O(n10656) );
  NAND_GATE U11255 ( .I1(n10657), .I2(n10656), .O(n10658) );
  NAND_GATE U11256 ( .I1(n10659), .I2(n10658), .O(n10660) );
  NAND_GATE U11257 ( .I1(n1416), .I2(A[14]), .O(n11099) );
  INV_GATE U11258 ( .I1(n11099), .O(n11093) );
  NAND_GATE U11259 ( .I1(n1416), .I2(A[13]), .O(n11275) );
  INV_GATE U11260 ( .I1(n11275), .O(n10825) );
  OR_GATE U11261 ( .I1(n10664), .I2(n10663), .O(n10673) );
  NAND_GATE U11262 ( .I1(n10665), .I2(n10664), .O(n10669) );
  NAND_GATE U11263 ( .I1(n10666), .I2(n10669), .O(n10672) );
  NAND_GATE U11264 ( .I1(n10667), .I2(n656), .O(n10668) );
  NAND_GATE U11265 ( .I1(n10669), .I2(n10668), .O(n10670) );
  NAND_GATE U11266 ( .I1(n10825), .I2(n11273), .O(n11270) );
  NAND_GATE U11267 ( .I1(n1416), .I2(A[12]), .O(n11111) );
  INV_GATE U11268 ( .I1(n11111), .O(n11105) );
  OR_GATE U11269 ( .I1(n10675), .I2(n10674), .O(n10687) );
  NAND_GATE U11270 ( .I1(n10676), .I2(n10675), .O(n10681) );
  NAND_GATE U11271 ( .I1(n10677), .I2(n10681), .O(n10685) );
  NAND_GATE U11272 ( .I1(n10679), .I2(n10678), .O(n10680) );
  NAND_GATE U11273 ( .I1(n10681), .I2(n10680), .O(n10682) );
  NAND_GATE U11274 ( .I1(n10683), .I2(n10682), .O(n10684) );
  NAND_GATE U11275 ( .I1(n10685), .I2(n10684), .O(n10686) );
  NAND_GATE U11276 ( .I1(n10687), .I2(n10686), .O(n11120) );
  OR_GATE U11277 ( .I1(n10688), .I2(n10692), .O(n10691) );
  OR_GATE U11278 ( .I1(n10689), .I2(n10693), .O(n10690) );
  NAND_GATE U11279 ( .I1(n10692), .I2(n1058), .O(n10696) );
  NAND3_GATE U11280 ( .I1(n10696), .I2(n10695), .I3(n10694), .O(n10697) );
  INV_GATE U11281 ( .I1(n11128), .O(n11131) );
  OR_GATE U11282 ( .I1(n10698), .I2(n10700), .O(n10711) );
  NAND_GATE U11283 ( .I1(n10700), .I2(n10699), .O(n10705) );
  NAND_GATE U11284 ( .I1(n10701), .I2(n10705), .O(n10709) );
  NAND_GATE U11285 ( .I1(n10703), .I2(n10702), .O(n10704) );
  NAND_GATE U11286 ( .I1(n10705), .I2(n10704), .O(n10706) );
  NAND_GATE U11287 ( .I1(n10707), .I2(n10706), .O(n10708) );
  NAND_GATE U11288 ( .I1(n10709), .I2(n10708), .O(n10710) );
  NAND_GATE U11289 ( .I1(n10711), .I2(n10710), .O(n11144) );
  OR_GATE U11290 ( .I1(n10712), .I2(n10716), .O(n10715) );
  OR_GATE U11291 ( .I1(n10713), .I2(n10717), .O(n10714) );
  AND_GATE U11292 ( .I1(n10715), .I2(n10714), .O(n10722) );
  NAND_GATE U11293 ( .I1(n10716), .I2(n1069), .O(n10720) );
  NAND3_GATE U11294 ( .I1(n10720), .I2(n10719), .I3(n10718), .O(n10721) );
  NAND_GATE U11295 ( .I1(n10722), .I2(n10721), .O(n11152) );
  INV_GATE U11296 ( .I1(n11152), .O(n11155) );
  OR_GATE U11297 ( .I1(n10723), .I2(n10725), .O(n10736) );
  NAND_GATE U11298 ( .I1(n10725), .I2(n10724), .O(n10730) );
  NAND_GATE U11299 ( .I1(n10726), .I2(n10730), .O(n10734) );
  NAND_GATE U11300 ( .I1(n10728), .I2(n10727), .O(n10729) );
  NAND_GATE U11301 ( .I1(n10730), .I2(n10729), .O(n10731) );
  NAND_GATE U11302 ( .I1(n10732), .I2(n10731), .O(n10733) );
  NAND_GATE U11303 ( .I1(n10734), .I2(n10733), .O(n10735) );
  NAND_GATE U11304 ( .I1(n10736), .I2(n10735), .O(n11168) );
  OR_GATE U11305 ( .I1(n10737), .I2(n10741), .O(n10740) );
  OR_GATE U11306 ( .I1(n10738), .I2(n10742), .O(n10739) );
  AND_GATE U11307 ( .I1(n10740), .I2(n10739), .O(n10747) );
  NAND_GATE U11308 ( .I1(n10741), .I2(n1179), .O(n10745) );
  NAND3_GATE U11309 ( .I1(n10745), .I2(n10744), .I3(n10743), .O(n10746) );
  NAND_GATE U11310 ( .I1(n10747), .I2(n10746), .O(n11177) );
  INV_GATE U11311 ( .I1(n11177), .O(n11180) );
  OR_GATE U11312 ( .I1(n10748), .I2(n10750), .O(n10761) );
  NAND_GATE U11313 ( .I1(n10750), .I2(n10749), .O(n10755) );
  NAND_GATE U11314 ( .I1(n10751), .I2(n10755), .O(n10759) );
  NAND_GATE U11315 ( .I1(n10753), .I2(n10752), .O(n10754) );
  NAND_GATE U11316 ( .I1(n10755), .I2(n10754), .O(n10756) );
  NAND_GATE U11317 ( .I1(n10757), .I2(n10756), .O(n10758) );
  NAND_GATE U11318 ( .I1(n10759), .I2(n10758), .O(n10760) );
  NAND_GATE U11319 ( .I1(n10761), .I2(n10760), .O(n11193) );
  OR_GATE U11320 ( .I1(n10762), .I2(n10766), .O(n10765) );
  OR_GATE U11321 ( .I1(n10763), .I2(n10767), .O(n10764) );
  AND_GATE U11322 ( .I1(n10765), .I2(n10764), .O(n10772) );
  NAND_GATE U11323 ( .I1(n10766), .I2(n1243), .O(n10770) );
  NAND3_GATE U11324 ( .I1(n10770), .I2(n10769), .I3(n10768), .O(n10771) );
  NAND_GATE U11325 ( .I1(n10772), .I2(n10771), .O(n11202) );
  INV_GATE U11326 ( .I1(n11202), .O(n11205) );
  INV_GATE U11327 ( .I1(n10773), .O(n10774) );
  NAND_GATE U11328 ( .I1(n10778), .I2(n10774), .O(n10786) );
  NAND_GATE U11329 ( .I1(n10776), .I2(n10780), .O(n10784) );
  NAND_GATE U11330 ( .I1(n10778), .I2(n10777), .O(n10779) );
  NAND_GATE U11331 ( .I1(n10780), .I2(n10779), .O(n10781) );
  NAND_GATE U11332 ( .I1(n10782), .I2(n10781), .O(n10783) );
  NAND_GATE U11333 ( .I1(n10784), .I2(n10783), .O(n10785) );
  NAND_GATE U11334 ( .I1(n10786), .I2(n10785), .O(n11218) );
  NAND_GATE U11335 ( .I1(n1419), .I2(A[0]), .O(n10787) );
  NAND_GATE U11336 ( .I1(n14241), .I2(n10787), .O(n10788) );
  NAND_GATE U11337 ( .I1(B[10]), .I2(n10788), .O(n10792) );
  NAND_GATE U11338 ( .I1(n1420), .I2(A[1]), .O(n10789) );
  NAND_GATE U11339 ( .I1(n724), .I2(n10789), .O(n10790) );
  NAND_GATE U11340 ( .I1(n1418), .I2(n10790), .O(n10791) );
  NAND_GATE U11341 ( .I1(n10792), .I2(n10791), .O(n11230) );
  NAND_GATE U11342 ( .I1(n1416), .I2(A[2]), .O(n11234) );
  NAND3_GATE U11343 ( .I1(n1416), .I2(n1418), .I3(n1254), .O(n11227) );
  NAND_GATE U11344 ( .I1(n11234), .I2(n11227), .O(n10793) );
  NAND_GATE U11345 ( .I1(n11230), .I2(n10793), .O(n10794) );
  INV_GATE U11346 ( .I1(n11234), .O(n11228) );
  INV_GATE U11347 ( .I1(n11227), .O(n11229) );
  NAND_GATE U11348 ( .I1(n11228), .I2(n11229), .O(n11225) );
  NAND_GATE U11349 ( .I1(n10794), .I2(n11225), .O(n11219) );
  NAND_GATE U11350 ( .I1(n11218), .I2(n11219), .O(n10796) );
  NAND_GATE U11351 ( .I1(n1415), .I2(A[3]), .O(n11220) );
  INV_GATE U11352 ( .I1(n11220), .O(n10795) );
  NAND_GATE U11353 ( .I1(n11218), .I2(n10795), .O(n11215) );
  NAND_GATE U11354 ( .I1(n11219), .I2(n10795), .O(n11214) );
  NAND3_GATE U11355 ( .I1(n10796), .I2(n11215), .I3(n11214), .O(n11204) );
  INV_GATE U11356 ( .I1(n11204), .O(n11201) );
  NAND_GATE U11357 ( .I1(n1415), .I2(A[4]), .O(n11209) );
  NAND_GATE U11358 ( .I1(n11201), .I2(n11209), .O(n10797) );
  NAND_GATE U11359 ( .I1(n11205), .I2(n10797), .O(n10798) );
  INV_GATE U11360 ( .I1(n11209), .O(n11203) );
  NAND_GATE U11361 ( .I1(n11204), .I2(n11203), .O(n11200) );
  NAND_GATE U11362 ( .I1(n10798), .I2(n11200), .O(n11194) );
  NAND_GATE U11363 ( .I1(n11193), .I2(n11194), .O(n10800) );
  NAND_GATE U11364 ( .I1(n1415), .I2(A[5]), .O(n11195) );
  INV_GATE U11365 ( .I1(n11195), .O(n10799) );
  NAND_GATE U11366 ( .I1(n11193), .I2(n10799), .O(n11190) );
  NAND_GATE U11367 ( .I1(n11194), .I2(n10799), .O(n11189) );
  NAND3_GATE U11368 ( .I1(n10800), .I2(n11190), .I3(n11189), .O(n11179) );
  INV_GATE U11369 ( .I1(n11179), .O(n11176) );
  NAND_GATE U11370 ( .I1(n1415), .I2(A[6]), .O(n11184) );
  NAND_GATE U11371 ( .I1(n11176), .I2(n11184), .O(n10801) );
  NAND_GATE U11372 ( .I1(n11180), .I2(n10801), .O(n10802) );
  INV_GATE U11373 ( .I1(n11184), .O(n11178) );
  NAND_GATE U11374 ( .I1(n11179), .I2(n11178), .O(n11175) );
  NAND_GATE U11375 ( .I1(n10802), .I2(n11175), .O(n11169) );
  NAND_GATE U11376 ( .I1(n11168), .I2(n11169), .O(n10804) );
  NAND_GATE U11377 ( .I1(n1415), .I2(A[7]), .O(n11170) );
  INV_GATE U11378 ( .I1(n11170), .O(n10803) );
  NAND_GATE U11379 ( .I1(n11168), .I2(n10803), .O(n11165) );
  NAND_GATE U11380 ( .I1(n11169), .I2(n10803), .O(n11164) );
  NAND3_GATE U11381 ( .I1(n10804), .I2(n11165), .I3(n11164), .O(n11154) );
  INV_GATE U11382 ( .I1(n11154), .O(n11151) );
  NAND_GATE U11383 ( .I1(n1415), .I2(A[8]), .O(n11159) );
  NAND_GATE U11384 ( .I1(n11151), .I2(n11159), .O(n10805) );
  NAND_GATE U11385 ( .I1(n11155), .I2(n10805), .O(n10806) );
  INV_GATE U11386 ( .I1(n11159), .O(n11153) );
  NAND_GATE U11387 ( .I1(n11154), .I2(n11153), .O(n11150) );
  NAND_GATE U11388 ( .I1(n10806), .I2(n11150), .O(n11145) );
  NAND_GATE U11389 ( .I1(n11144), .I2(n11145), .O(n10808) );
  NAND_GATE U11390 ( .I1(n1415), .I2(A[9]), .O(n11146) );
  INV_GATE U11391 ( .I1(n11146), .O(n10807) );
  NAND_GATE U11392 ( .I1(n11144), .I2(n10807), .O(n11141) );
  NAND_GATE U11393 ( .I1(n11145), .I2(n10807), .O(n11140) );
  NAND3_GATE U11394 ( .I1(n10808), .I2(n11141), .I3(n11140), .O(n11130) );
  INV_GATE U11395 ( .I1(n11130), .O(n11127) );
  NAND_GATE U11396 ( .I1(n1415), .I2(A[10]), .O(n11135) );
  NAND_GATE U11397 ( .I1(n11127), .I2(n11135), .O(n10809) );
  NAND_GATE U11398 ( .I1(n11131), .I2(n10809), .O(n10810) );
  INV_GATE U11399 ( .I1(n11135), .O(n11129) );
  NAND_GATE U11400 ( .I1(n11130), .I2(n11129), .O(n11126) );
  NAND_GATE U11401 ( .I1(n10810), .I2(n11126), .O(n11121) );
  NAND_GATE U11402 ( .I1(n11120), .I2(n11121), .O(n10812) );
  NAND_GATE U11403 ( .I1(n1415), .I2(A[11]), .O(n11122) );
  INV_GATE U11404 ( .I1(n11122), .O(n10811) );
  NAND_GATE U11405 ( .I1(n11120), .I2(n10811), .O(n11117) );
  NAND_GATE U11406 ( .I1(n11121), .I2(n10811), .O(n11116) );
  NAND3_GATE U11407 ( .I1(n10812), .I2(n11117), .I3(n11116), .O(n11107) );
  NAND_GATE U11408 ( .I1(n11105), .I2(n11107), .O(n11102) );
  OR_GATE U11409 ( .I1(n10813), .I2(n10817), .O(n10816) );
  OR_GATE U11410 ( .I1(n10818), .I2(n10814), .O(n10815) );
  NAND_GATE U11411 ( .I1(n10817), .I2(n1035), .O(n10821) );
  NAND3_GATE U11412 ( .I1(n10821), .I2(n10820), .I3(n10819), .O(n10822) );
  INV_GATE U11413 ( .I1(n11103), .O(n11106) );
  INV_GATE U11414 ( .I1(n11107), .O(n11104) );
  NAND_GATE U11415 ( .I1(n11111), .I2(n11104), .O(n10823) );
  NAND_GATE U11416 ( .I1(n11106), .I2(n10823), .O(n10824) );
  NAND_GATE U11417 ( .I1(n11102), .I2(n10824), .O(n11274) );
  NAND_GATE U11418 ( .I1(n11273), .I2(n11274), .O(n10826) );
  NAND_GATE U11419 ( .I1(n10825), .I2(n11274), .O(n11269) );
  NAND3_GATE U11420 ( .I1(n11270), .I2(n10826), .I3(n11269), .O(n11095) );
  NAND_GATE U11421 ( .I1(n11093), .I2(n11095), .O(n11090) );
  OR_GATE U11422 ( .I1(n10827), .I2(n10831), .O(n10830) );
  OR_GATE U11423 ( .I1(n10832), .I2(n10828), .O(n10829) );
  AND_GATE U11424 ( .I1(n10830), .I2(n10829), .O(n10837) );
  NAND_GATE U11425 ( .I1(n10831), .I2(n1003), .O(n10835) );
  NAND3_GATE U11426 ( .I1(n10835), .I2(n10834), .I3(n10833), .O(n10836) );
  NAND_GATE U11427 ( .I1(n10837), .I2(n10836), .O(n11091) );
  INV_GATE U11428 ( .I1(n11091), .O(n11094) );
  INV_GATE U11429 ( .I1(n11095), .O(n11092) );
  NAND_GATE U11430 ( .I1(n11094), .I2(n10838), .O(n10839) );
  NAND_GATE U11431 ( .I1(n11090), .I2(n10839), .O(n11288) );
  NAND_GATE U11432 ( .I1(n11287), .I2(n11288), .O(n10841) );
  NAND_GATE U11433 ( .I1(n10840), .I2(n11288), .O(n11283) );
  NAND3_GATE U11434 ( .I1(n11284), .I2(n10841), .I3(n11283), .O(n11298) );
  NAND_GATE U11435 ( .I1(n11296), .I2(n11298), .O(n11295) );
  OR_GATE U11436 ( .I1(n10842), .I2(n10846), .O(n10845) );
  OR_GATE U11437 ( .I1(n10847), .I2(n10843), .O(n10844) );
  AND_GATE U11438 ( .I1(n10845), .I2(n10844), .O(n10852) );
  NAND_GATE U11439 ( .I1(n998), .I2(n10847), .O(n10849) );
  NAND3_GATE U11440 ( .I1(n10850), .I2(n10849), .I3(n10848), .O(n10851) );
  NAND_GATE U11441 ( .I1(n10852), .I2(n10851), .O(n11299) );
  NAND_GATE U11442 ( .I1(n11303), .I2(n35), .O(n10853) );
  NAND_GATE U11443 ( .I1(n11297), .I2(n10853), .O(n10854) );
  NAND_GATE U11444 ( .I1(n11295), .I2(n10854), .O(n11085) );
  NAND_GATE U11445 ( .I1(n10866), .I2(n11085), .O(n11081) );
  OR_GATE U11446 ( .I1(n10858), .I2(n10855), .O(n10865) );
  NAND_GATE U11447 ( .I1(n10856), .I2(n10860), .O(n10863) );
  NAND_GATE U11448 ( .I1(n10859), .I2(n10858), .O(n10860) );
  NAND_GATE U11449 ( .I1(n10863), .I2(n10862), .O(n10864) );
  NAND_GATE U11450 ( .I1(n10865), .I2(n10864), .O(n11084) );
  NAND_GATE U11451 ( .I1(n11085), .I2(n11084), .O(n10867) );
  NAND_GATE U11452 ( .I1(n10866), .I2(n11084), .O(n11080) );
  NAND3_GATE U11453 ( .I1(n11081), .I2(n10867), .I3(n11080), .O(n11314) );
  NAND_GATE U11454 ( .I1(n1415), .I2(A[18]), .O(n11317) );
  OR_GATE U11455 ( .I1(n10868), .I2(n10872), .O(n10871) );
  OR_GATE U11456 ( .I1(n10873), .I2(n10869), .O(n10870) );
  AND_GATE U11457 ( .I1(n10871), .I2(n10870), .O(n10878) );
  NAND_GATE U11458 ( .I1(n58), .I2(n10873), .O(n10874) );
  NAND3_GATE U11459 ( .I1(n10876), .I2(n10875), .I3(n10874), .O(n10877) );
  NAND_GATE U11460 ( .I1(n10878), .I2(n10877), .O(n11310) );
  NAND_GATE U11461 ( .I1(n11317), .I2(n11310), .O(n10879) );
  NAND_GATE U11462 ( .I1(n11314), .I2(n10879), .O(n10881) );
  INV_GATE U11463 ( .I1(n11317), .O(n11312) );
  INV_GATE U11464 ( .I1(n11310), .O(n11313) );
  NAND_GATE U11465 ( .I1(n11312), .I2(n11313), .O(n10880) );
  NAND_GATE U11466 ( .I1(n10881), .I2(n10880), .O(n11327) );
  NAND_GATE U11467 ( .I1(n10892), .I2(n11327), .O(n11331) );
  INV_GATE U11468 ( .I1(n10884), .O(n10886) );
  NAND_GATE U11469 ( .I1(n10882), .I2(n10888), .O(n11325) );
  NAND_GATE U11470 ( .I1(n10885), .I2(n10884), .O(n10889) );
  NAND_GATE U11471 ( .I1(n10887), .I2(n10886), .O(n10888) );
  NAND_GATE U11472 ( .I1(n10889), .I2(n10888), .O(n11323) );
  NAND_GATE U11473 ( .I1(n11324), .I2(n11323), .O(n10890) );
  NAND3_GATE U11474 ( .I1(n11327), .I2(n10891), .I3(n10890), .O(n10893) );
  NAND3_GATE U11475 ( .I1(n10892), .I2(n10891), .I3(n10890), .O(n11322) );
  NAND3_GATE U11476 ( .I1(n11331), .I2(n10893), .I3(n11322), .O(n11347) );
  NAND_GATE U11477 ( .I1(n11342), .I2(n11343), .O(n10894) );
  NAND_GATE U11478 ( .I1(n11347), .I2(n10894), .O(n10895) );
  NAND_GATE U11479 ( .I1(n11346), .I2(n10895), .O(n11074) );
  INV_GATE U11480 ( .I1(n10903), .O(n10897) );
  NAND_GATE U11481 ( .I1(n10898), .I2(n10897), .O(n10896) );
  NAND_GATE U11482 ( .I1(n482), .I2(n10896), .O(n10901) );
  NAND_GATE U11483 ( .I1(n10901), .I2(n10900), .O(n10905) );
  NAND_GATE U11484 ( .I1(n279), .I2(n10903), .O(n10904) );
  NAND_GATE U11485 ( .I1(n10905), .I2(n10904), .O(n11075) );
  NAND_GATE U11486 ( .I1(n11074), .I2(n11075), .O(n10907) );
  NAND_GATE U11487 ( .I1(n1415), .I2(A[21]), .O(n11078) );
  INV_GATE U11488 ( .I1(n11078), .O(n10906) );
  NAND_GATE U11489 ( .I1(n10906), .I2(n11075), .O(n11070) );
  NAND_GATE U11490 ( .I1(n10906), .I2(n11074), .O(n11071) );
  NAND3_GATE U11491 ( .I1(n10907), .I2(n11070), .I3(n11071), .O(n11362) );
  NAND_GATE U11492 ( .I1(n11355), .I2(n11357), .O(n10908) );
  NAND_GATE U11493 ( .I1(n10909), .I2(n11066), .O(n11063) );
  AND_GATE U11494 ( .I1(n11065), .I2(n11063), .O(n10914) );
  NAND_GATE U11495 ( .I1(n10910), .I2(n11057), .O(n10911) );
  NAND_GATE U11496 ( .I1(n10912), .I2(n10911), .O(n11064) );
  NAND_GATE U11497 ( .I1(n11066), .I2(n11064), .O(n10913) );
  NAND_GATE U11498 ( .I1(n11374), .I2(n11375), .O(n10915) );
  NAND_GATE U11499 ( .I1(n287), .I2(n10915), .O(n10916) );
  NAND_GATE U11500 ( .I1(n11372), .I2(n10916), .O(n11046) );
  NAND_GATE U11501 ( .I1(n10921), .I2(n11046), .O(n11037) );
  NAND_GATE U11502 ( .I1(n968), .I2(n10924), .O(n10917) );
  NAND_GATE U11503 ( .I1(n884), .I2(n10917), .O(n10918) );
  NAND_GATE U11504 ( .I1(n10921), .I2(n11048), .O(n10922) );
  INV_GATE U11505 ( .I1(n10922), .O(n11042) );
  NAND3_GATE U11506 ( .I1(n10925), .I2(n10924), .I3(n10923), .O(n10927) );
  NAND_GATE U11507 ( .I1(n884), .I2(n10927), .O(n10928) );
  NAND_GATE U11508 ( .I1(n10929), .I2(n10928), .O(n11043) );
  NAND_GATE U11509 ( .I1(n11044), .I2(n11043), .O(n11041) );
  NAND3_GATE U11510 ( .I1(n11046), .I2(n11048), .I3(n11041), .O(n10930) );
  NAND3_GATE U11511 ( .I1(n11037), .I2(n10931), .I3(n10930), .O(n11394) );
  NAND_GATE U11512 ( .I1(n11390), .I2(n11394), .O(n10933) );
  NAND3_GATE U11513 ( .I1(n11392), .I2(n11394), .I3(n11386), .O(n10932) );
  NAND3_GATE U11514 ( .I1(n10934), .I2(n10933), .I3(n10932), .O(n11026) );
  NAND_GATE U11515 ( .I1(n11033), .I2(n11026), .O(n11030) );
  NAND3_GATE U11516 ( .I1(n10935), .I2(n10938), .I3(n677), .O(n11020) );
  INV_GATE U11517 ( .I1(n10938), .O(n10936) );
  NAND_GATE U11518 ( .I1(n10935), .I2(n10940), .O(n11019) );
  NAND_GATE U11519 ( .I1(n10937), .I2(n10936), .O(n10940) );
  NAND_GATE U11520 ( .I1(n677), .I2(n10938), .O(n10939) );
  NAND_GATE U11521 ( .I1(n10940), .I2(n10939), .O(n11021) );
  NAND_GATE U11522 ( .I1(n11019), .I2(n11024), .O(n10941) );
  NAND_GATE U11523 ( .I1(n11020), .I2(n10941), .O(n11031) );
  NAND_GATE U11524 ( .I1(n11033), .I2(n11031), .O(n10943) );
  NAND_GATE U11525 ( .I1(n11026), .I2(n11031), .O(n10942) );
  NAND3_GATE U11526 ( .I1(n11030), .I2(n10943), .I3(n10942), .O(n11004) );
  NAND3_GATE U11527 ( .I1(n10945), .I2(n10944), .I3(n11004), .O(n10946) );
  NAND_GATE U11528 ( .I1(n11013), .I2(n11004), .O(n11014) );
  NAND3_GATE U11529 ( .I1(n10947), .I2(n10946), .I3(n11014), .O(n10995) );
  NAND_GATE U11530 ( .I1(n10999), .I2(n10995), .O(n10954) );
  NAND_GATE U11531 ( .I1(n10949), .I2(n10948), .O(n10950) );
  NAND_GATE U11532 ( .I1(n10951), .I2(n10950), .O(n10952) );
  NAND_GATE U11533 ( .I1(n10952), .I2(n10992), .O(n10994) );
  NAND3_GATE U11534 ( .I1(n10955), .I2(n10954), .I3(n10953), .O(n10981) );
  INV_GATE U11535 ( .I1(n10962), .O(n10960) );
  NAND_GATE U11536 ( .I1(n10961), .I2(n10960), .O(n10958) );
  NAND3_GATE U11537 ( .I1(n10959), .I2(n10958), .I3(n10957), .O(n10966) );
  NAND_GATE U11538 ( .I1(n10966), .I2(n10967), .O(n10980) );
  NAND_GATE U11539 ( .I1(n1415), .I2(A[30]), .O(n10984) );
  INV_GATE U11540 ( .I1(n10984), .O(n10965) );
  NAND_GATE U11541 ( .I1(n10965), .I2(n10981), .O(n10978) );
  NAND3_GATE U11542 ( .I1(n10967), .I2(n10966), .I3(n10965), .O(n10977) );
  NAND3_GATE U11543 ( .I1(n10971), .I2(n10972), .I3(n951), .O(n10968) );
  NAND_GATE U11544 ( .I1(n10973), .I2(n10968), .O(n10976) );
  NAND_GATE U11545 ( .I1(n1320), .I2(n10976), .O(n10970) );
  INV_GATE U11546 ( .I1(n10976), .O(n14819) );
  NAND_GATE U11547 ( .I1(n10970), .I2(n10969), .O(\A1[38] ) );
  NAND3_GATE U11548 ( .I1(n10972), .I2(n951), .I3(n10971), .O(n10974) );
  OR_GATE U11549 ( .I1(n10974), .I2(n10973), .O(n10975) );
  NAND_GATE U11550 ( .I1(n10976), .I2(n10975), .O(n11411) );
  OR_GATE U11551 ( .I1(n10977), .I2(n10981), .O(n10987) );
  INV_GATE U11552 ( .I1(n10978), .O(n10979) );
  NAND_GATE U11553 ( .I1(n10981), .I2(n10980), .O(n10982) );
  NAND3_GATE U11554 ( .I1(n10984), .I2(n10983), .I3(n10982), .O(n10985) );
  NAND3_GATE U11555 ( .I1(n10987), .I2(n10986), .I3(n10985), .O(n11414) );
  NAND_GATE U11556 ( .I1(n1413), .I2(A[30]), .O(n11790) );
  NAND_GATE U11557 ( .I1(n10989), .I2(n10988), .O(n10992) );
  INV_GATE U11558 ( .I1(n10995), .O(n10997) );
  NAND3_GATE U11559 ( .I1(n10998), .I2(n10992), .I3(n10997), .O(n10990) );
  AND_GATE U11560 ( .I1(n10991), .I2(n10990), .O(n11788) );
  NAND_GATE U11561 ( .I1(n10998), .I2(n10992), .O(n10993) );
  NAND_GATE U11562 ( .I1(n10995), .I2(n10993), .O(n11787) );
  AND_GATE U11563 ( .I1(n11788), .I2(n11787), .O(n11002) );
  NAND4_GATE U11564 ( .I1(n10996), .I2(n10995), .I3(n10999), .I4(n10994), .O(
        n11001) );
  NAND4_GATE U11565 ( .I1(n10999), .I2(n10998), .I3(n10992), .I4(n10997), .O(
        n11000) );
  NAND_GATE U11566 ( .I1(n11001), .I2(n11000), .O(n11786) );
  OR_GATE U11567 ( .I1(n11002), .I2(n11786), .O(n11789) );
  NAND_GATE U11568 ( .I1(n10944), .I2(n10945), .O(n11003) );
  NAND_GATE U11569 ( .I1(n11004), .I2(n11003), .O(n11007) );
  NAND3_GATE U11570 ( .I1(n10944), .I2(n10945), .I3(n11012), .O(n11006) );
  NAND3_GATE U11571 ( .I1(n11007), .I2(n11006), .I3(n11005), .O(n11018) );
  NAND_GATE U11572 ( .I1(n11011), .I2(n11010), .O(n11015) );
  NAND3_GATE U11573 ( .I1(n11013), .I2(n11012), .I3(n11015), .O(n11017) );
  OR_GATE U11574 ( .I1(n11015), .I2(n11014), .O(n11016) );
  NAND3_GATE U11575 ( .I1(n11018), .I2(n11017), .I3(n11016), .O(n11416) );
  NAND_GATE U11576 ( .I1(n1413), .I2(A[29]), .O(n11809) );
  INV_GATE U11577 ( .I1(n11809), .O(n11807) );
  NAND_GATE U11578 ( .I1(n781), .I2(n11807), .O(n11409) );
  NAND_GATE U11579 ( .I1(n1413), .I2(A[28]), .O(n11827) );
  INV_GATE U11580 ( .I1(n11827), .O(n11774) );
  INV_GATE U11581 ( .I1(n11026), .O(n11032) );
  NAND_GATE U11582 ( .I1(n11022), .I2(n11021), .O(n11024) );
  NAND3_GATE U11583 ( .I1(n11023), .I2(n11032), .I3(n11024), .O(n11028) );
  NAND_GATE U11584 ( .I1(n11024), .I2(n11023), .O(n11025) );
  NAND_GATE U11585 ( .I1(n11026), .I2(n11025), .O(n11027) );
  NAND3_GATE U11586 ( .I1(n11029), .I2(n11028), .I3(n11027), .O(n11036) );
  OR_GATE U11587 ( .I1(n11031), .I2(n11030), .O(n11035) );
  NAND3_GATE U11588 ( .I1(n11033), .I2(n11032), .I3(n11031), .O(n11034) );
  NAND3_GATE U11589 ( .I1(n11036), .I2(n11035), .I3(n11034), .O(n11776) );
  NAND_GATE U11590 ( .I1(n11774), .I2(n11778), .O(n11406) );
  NAND_GATE U11591 ( .I1(n1413), .I2(A[27]), .O(n11842) );
  INV_GATE U11592 ( .I1(n11842), .O(n11768) );
  NAND_GATE U11593 ( .I1(n1413), .I2(A[26]), .O(n11850) );
  INV_GATE U11594 ( .I1(n11037), .O(n11038) );
  NAND3_GATE U11595 ( .I1(n11040), .I2(n11039), .I3(n11038), .O(n11054) );
  INV_GATE U11596 ( .I1(n11046), .O(n11047) );
  NAND3_GATE U11597 ( .I1(n11042), .I2(n11041), .I3(n11047), .O(n11053) );
  NAND_GATE U11598 ( .I1(n11048), .I2(n11041), .O(n11045) );
  NAND_GATE U11599 ( .I1(n11046), .I2(n11045), .O(n11051) );
  NAND3_GATE U11600 ( .I1(n11048), .I2(n11041), .I3(n11047), .O(n11050) );
  NAND3_GATE U11601 ( .I1(n11051), .I2(n11050), .I3(n11049), .O(n11052) );
  NAND3_GATE U11602 ( .I1(n11054), .I2(n11053), .I3(n11052), .O(n11851) );
  NAND_GATE U11603 ( .I1(n1413), .I2(A[25]), .O(n11427) );
  INV_GATE U11604 ( .I1(n11427), .O(n11422) );
  NAND_GATE U11605 ( .I1(n11056), .I2(n11055), .O(n11057) );
  NAND3_GATE U11606 ( .I1(n11057), .I2(n636), .I3(n11058), .O(n11062) );
  NAND_GATE U11607 ( .I1(n11058), .I2(n11057), .O(n11059) );
  NAND_GATE U11608 ( .I1(n11066), .I2(n11059), .O(n11061) );
  NAND3_GATE U11609 ( .I1(n11062), .I2(n11061), .I3(n11060), .O(n11069) );
  OR_GATE U11610 ( .I1(n11064), .I2(n11063), .O(n11068) );
  OR_GATE U11611 ( .I1(n11066), .I2(n11065), .O(n11067) );
  NAND3_GATE U11612 ( .I1(n11069), .I2(n11068), .I3(n11067), .O(n11751) );
  INV_GATE U11613 ( .I1(n11751), .O(n11748) );
  NAND_GATE U11614 ( .I1(n1413), .I2(A[24]), .O(n11749) );
  INV_GATE U11615 ( .I1(n11749), .O(n11743) );
  NAND_GATE U11616 ( .I1(n11748), .I2(n11743), .O(n11744) );
  NAND_GATE U11617 ( .I1(n1413), .I2(A[23]), .O(n11434) );
  INV_GATE U11618 ( .I1(n11434), .O(n11365) );
  OR_GATE U11619 ( .I1(n11070), .I2(n11074), .O(n11073) );
  OR_GATE U11620 ( .I1(n11075), .I2(n11071), .O(n11072) );
  NAND_GATE U11621 ( .I1(n469), .I2(n11075), .O(n11076) );
  NAND3_GATE U11622 ( .I1(n11078), .I2(n11077), .I3(n11076), .O(n11079) );
  INV_GATE U11623 ( .I1(n11729), .O(n11731) );
  NAND_GATE U11624 ( .I1(n1413), .I2(A[22]), .O(n11890) );
  INV_GATE U11625 ( .I1(n11890), .O(n11725) );
  NAND_GATE U11626 ( .I1(n11731), .I2(n11725), .O(n11726) );
  NAND_GATE U11627 ( .I1(n1413), .I2(A[21]), .O(n11445) );
  INV_GATE U11628 ( .I1(n11445), .O(n11446) );
  NAND_GATE U11629 ( .I1(n1413), .I2(A[19]), .O(n11461) );
  INV_GATE U11630 ( .I1(n11461), .O(n11320) );
  OR_GATE U11631 ( .I1(n11080), .I2(n11085), .O(n11083) );
  OR_GATE U11632 ( .I1(n11084), .I2(n11081), .O(n11082) );
  NAND_GATE U11633 ( .I1(n129), .I2(n11084), .O(n11088) );
  NAND3_GATE U11634 ( .I1(n11088), .I2(n11087), .I3(n11086), .O(n11089) );
  INV_GATE U11635 ( .I1(n11704), .O(n11706) );
  NAND_GATE U11636 ( .I1(n1413), .I2(A[18]), .O(n11707) );
  INV_GATE U11637 ( .I1(n11707), .O(n11702) );
  NAND_GATE U11638 ( .I1(n11706), .I2(n11702), .O(n11699) );
  NAND_GATE U11639 ( .I1(n1413), .I2(A[17]), .O(n11471) );
  INV_GATE U11640 ( .I1(n11471), .O(n11306) );
  NAND_GATE U11641 ( .I1(n1413), .I2(A[16]), .O(n11691) );
  INV_GATE U11642 ( .I1(n11691), .O(n11685) );
  NAND_GATE U11643 ( .I1(n1413), .I2(A[15]), .O(n11676) );
  INV_GATE U11644 ( .I1(n11676), .O(n11281) );
  OR_GATE U11645 ( .I1(n11091), .I2(n11090), .O(n11101) );
  NAND_GATE U11646 ( .I1(n11092), .I2(n11091), .O(n11097) );
  NAND_GATE U11647 ( .I1(n11093), .I2(n11097), .O(n11100) );
  NAND_GATE U11648 ( .I1(n11097), .I2(n11096), .O(n11098) );
  NAND_GATE U11649 ( .I1(n11281), .I2(n11674), .O(n11671) );
  NAND_GATE U11650 ( .I1(n1413), .I2(A[14]), .O(n11483) );
  INV_GATE U11651 ( .I1(n11483), .O(n11477) );
  OR_GATE U11652 ( .I1(n11103), .I2(n11102), .O(n11115) );
  NAND_GATE U11653 ( .I1(n11104), .I2(n11103), .O(n11109) );
  NAND_GATE U11654 ( .I1(n11105), .I2(n11109), .O(n11113) );
  NAND_GATE U11655 ( .I1(n11107), .I2(n11106), .O(n11108) );
  NAND_GATE U11656 ( .I1(n11109), .I2(n11108), .O(n11110) );
  NAND_GATE U11657 ( .I1(n11111), .I2(n11110), .O(n11112) );
  NAND_GATE U11658 ( .I1(n11113), .I2(n11112), .O(n11114) );
  NAND_GATE U11659 ( .I1(n11115), .I2(n11114), .O(n11492) );
  OR_GATE U11660 ( .I1(n11116), .I2(n11120), .O(n11119) );
  OR_GATE U11661 ( .I1(n11117), .I2(n11121), .O(n11118) );
  NAND_GATE U11662 ( .I1(n11120), .I2(n1052), .O(n11124) );
  NAND3_GATE U11663 ( .I1(n11124), .I2(n11123), .I3(n11122), .O(n11125) );
  INV_GATE U11664 ( .I1(n11500), .O(n11503) );
  OR_GATE U11665 ( .I1(n11126), .I2(n11128), .O(n11139) );
  NAND_GATE U11666 ( .I1(n11128), .I2(n11127), .O(n11133) );
  NAND_GATE U11667 ( .I1(n11129), .I2(n11133), .O(n11137) );
  NAND_GATE U11668 ( .I1(n11131), .I2(n11130), .O(n11132) );
  NAND_GATE U11669 ( .I1(n11133), .I2(n11132), .O(n11134) );
  NAND_GATE U11670 ( .I1(n11135), .I2(n11134), .O(n11136) );
  NAND_GATE U11671 ( .I1(n11137), .I2(n11136), .O(n11138) );
  NAND_GATE U11672 ( .I1(n11139), .I2(n11138), .O(n11516) );
  OR_GATE U11673 ( .I1(n11140), .I2(n11144), .O(n11143) );
  OR_GATE U11674 ( .I1(n11141), .I2(n11145), .O(n11142) );
  NAND_GATE U11675 ( .I1(n11144), .I2(n1065), .O(n11148) );
  NAND3_GATE U11676 ( .I1(n11148), .I2(n11147), .I3(n11146), .O(n11149) );
  INV_GATE U11677 ( .I1(n11524), .O(n11527) );
  OR_GATE U11678 ( .I1(n11150), .I2(n11152), .O(n11163) );
  NAND_GATE U11679 ( .I1(n11152), .I2(n11151), .O(n11157) );
  NAND_GATE U11680 ( .I1(n11153), .I2(n11157), .O(n11161) );
  NAND_GATE U11681 ( .I1(n11155), .I2(n11154), .O(n11156) );
  NAND_GATE U11682 ( .I1(n11157), .I2(n11156), .O(n11158) );
  NAND_GATE U11683 ( .I1(n11159), .I2(n11158), .O(n11160) );
  NAND_GATE U11684 ( .I1(n11161), .I2(n11160), .O(n11162) );
  NAND_GATE U11685 ( .I1(n11163), .I2(n11162), .O(n11540) );
  OR_GATE U11686 ( .I1(n11164), .I2(n11168), .O(n11167) );
  OR_GATE U11687 ( .I1(n11165), .I2(n11169), .O(n11166) );
  AND_GATE U11688 ( .I1(n11167), .I2(n11166), .O(n11174) );
  NAND_GATE U11689 ( .I1(n11168), .I2(n1074), .O(n11172) );
  NAND3_GATE U11690 ( .I1(n11172), .I2(n11171), .I3(n11170), .O(n11173) );
  NAND_GATE U11691 ( .I1(n11174), .I2(n11173), .O(n11549) );
  INV_GATE U11692 ( .I1(n11549), .O(n11552) );
  OR_GATE U11693 ( .I1(n11175), .I2(n11177), .O(n11188) );
  NAND_GATE U11694 ( .I1(n11177), .I2(n11176), .O(n11182) );
  NAND_GATE U11695 ( .I1(n11178), .I2(n11182), .O(n11186) );
  NAND_GATE U11696 ( .I1(n11180), .I2(n11179), .O(n11181) );
  NAND_GATE U11697 ( .I1(n11182), .I2(n11181), .O(n11183) );
  NAND_GATE U11698 ( .I1(n11184), .I2(n11183), .O(n11185) );
  NAND_GATE U11699 ( .I1(n11186), .I2(n11185), .O(n11187) );
  NAND_GATE U11700 ( .I1(n11188), .I2(n11187), .O(n11565) );
  OR_GATE U11701 ( .I1(n11189), .I2(n11193), .O(n11192) );
  OR_GATE U11702 ( .I1(n11190), .I2(n11194), .O(n11191) );
  AND_GATE U11703 ( .I1(n11192), .I2(n11191), .O(n11199) );
  NAND_GATE U11704 ( .I1(n11193), .I2(n1184), .O(n11197) );
  NAND3_GATE U11705 ( .I1(n11197), .I2(n11196), .I3(n11195), .O(n11198) );
  NAND_GATE U11706 ( .I1(n11199), .I2(n11198), .O(n11574) );
  INV_GATE U11707 ( .I1(n11574), .O(n11577) );
  OR_GATE U11708 ( .I1(n11200), .I2(n11202), .O(n11213) );
  NAND_GATE U11709 ( .I1(n11202), .I2(n11201), .O(n11207) );
  NAND_GATE U11710 ( .I1(n11203), .I2(n11207), .O(n11211) );
  NAND_GATE U11711 ( .I1(n11205), .I2(n11204), .O(n11206) );
  NAND_GATE U11712 ( .I1(n11207), .I2(n11206), .O(n11208) );
  NAND_GATE U11713 ( .I1(n11209), .I2(n11208), .O(n11210) );
  NAND_GATE U11714 ( .I1(n11211), .I2(n11210), .O(n11212) );
  NAND_GATE U11715 ( .I1(n11213), .I2(n11212), .O(n11590) );
  OR_GATE U11716 ( .I1(n11214), .I2(n11218), .O(n11217) );
  OR_GATE U11717 ( .I1(n11215), .I2(n11219), .O(n11216) );
  AND_GATE U11718 ( .I1(n11217), .I2(n11216), .O(n11224) );
  NAND_GATE U11719 ( .I1(n11218), .I2(n1244), .O(n11222) );
  NAND3_GATE U11720 ( .I1(n11222), .I2(n11221), .I3(n11220), .O(n11223) );
  NAND_GATE U11721 ( .I1(n11224), .I2(n11223), .O(n11599) );
  INV_GATE U11722 ( .I1(n11599), .O(n11602) );
  INV_GATE U11723 ( .I1(n11225), .O(n11226) );
  NAND_GATE U11724 ( .I1(n11230), .I2(n11226), .O(n11238) );
  NAND_GATE U11725 ( .I1(n11228), .I2(n11232), .O(n11236) );
  NAND_GATE U11726 ( .I1(n11230), .I2(n11229), .O(n11231) );
  NAND_GATE U11727 ( .I1(n11232), .I2(n11231), .O(n11233) );
  NAND_GATE U11728 ( .I1(n11234), .I2(n11233), .O(n11235) );
  NAND_GATE U11729 ( .I1(n11236), .I2(n11235), .O(n11237) );
  NAND_GATE U11730 ( .I1(n11238), .I2(n11237), .O(n11615) );
  NAND_GATE U11731 ( .I1(n1417), .I2(A[0]), .O(n11239) );
  NAND_GATE U11732 ( .I1(n14241), .I2(n11239), .O(n11240) );
  NAND_GATE U11733 ( .I1(n1418), .I2(n11240), .O(n11244) );
  NAND_GATE U11734 ( .I1(n1419), .I2(A[1]), .O(n11241) );
  NAND_GATE U11735 ( .I1(n724), .I2(n11241), .O(n11242) );
  NAND_GATE U11736 ( .I1(n1415), .I2(n11242), .O(n11243) );
  NAND_GATE U11737 ( .I1(n11244), .I2(n11243), .O(n11627) );
  NAND_GATE U11738 ( .I1(n1413), .I2(A[2]), .O(n11631) );
  NAND3_GATE U11739 ( .I1(n1413), .I2(n1415), .I3(n1254), .O(n11624) );
  NAND_GATE U11740 ( .I1(n11631), .I2(n11624), .O(n11245) );
  NAND_GATE U11741 ( .I1(n11627), .I2(n11245), .O(n11246) );
  INV_GATE U11742 ( .I1(n11631), .O(n11625) );
  INV_GATE U11743 ( .I1(n11624), .O(n11626) );
  NAND_GATE U11744 ( .I1(n11625), .I2(n11626), .O(n11622) );
  NAND_GATE U11745 ( .I1(n11246), .I2(n11622), .O(n11616) );
  NAND_GATE U11746 ( .I1(n11615), .I2(n11616), .O(n11248) );
  NAND_GATE U11747 ( .I1(n1413), .I2(A[3]), .O(n11617) );
  INV_GATE U11748 ( .I1(n11617), .O(n11247) );
  NAND_GATE U11749 ( .I1(n11615), .I2(n11247), .O(n11612) );
  NAND_GATE U11750 ( .I1(n11616), .I2(n11247), .O(n11611) );
  NAND3_GATE U11751 ( .I1(n11248), .I2(n11612), .I3(n11611), .O(n11601) );
  INV_GATE U11752 ( .I1(n11601), .O(n11598) );
  NAND_GATE U11753 ( .I1(n1413), .I2(A[4]), .O(n11606) );
  NAND_GATE U11754 ( .I1(n11598), .I2(n11606), .O(n11249) );
  NAND_GATE U11755 ( .I1(n11602), .I2(n11249), .O(n11250) );
  INV_GATE U11756 ( .I1(n11606), .O(n11600) );
  NAND_GATE U11757 ( .I1(n11601), .I2(n11600), .O(n11597) );
  NAND_GATE U11758 ( .I1(n11250), .I2(n11597), .O(n11591) );
  NAND_GATE U11759 ( .I1(n11590), .I2(n11591), .O(n11252) );
  NAND_GATE U11760 ( .I1(n1413), .I2(A[5]), .O(n11592) );
  INV_GATE U11761 ( .I1(n11592), .O(n11251) );
  NAND_GATE U11762 ( .I1(n11590), .I2(n11251), .O(n11587) );
  NAND_GATE U11763 ( .I1(n11591), .I2(n11251), .O(n11586) );
  NAND3_GATE U11764 ( .I1(n11252), .I2(n11587), .I3(n11586), .O(n11576) );
  INV_GATE U11765 ( .I1(n11576), .O(n11573) );
  NAND_GATE U11766 ( .I1(n1413), .I2(A[6]), .O(n11581) );
  NAND_GATE U11767 ( .I1(n11573), .I2(n11581), .O(n11253) );
  NAND_GATE U11768 ( .I1(n11577), .I2(n11253), .O(n11254) );
  INV_GATE U11769 ( .I1(n11581), .O(n11575) );
  NAND_GATE U11770 ( .I1(n11576), .I2(n11575), .O(n11572) );
  NAND_GATE U11771 ( .I1(n11254), .I2(n11572), .O(n11566) );
  NAND_GATE U11772 ( .I1(n11565), .I2(n11566), .O(n11256) );
  NAND_GATE U11773 ( .I1(n1413), .I2(A[7]), .O(n11567) );
  INV_GATE U11774 ( .I1(n11567), .O(n11255) );
  NAND_GATE U11775 ( .I1(n11565), .I2(n11255), .O(n11562) );
  NAND_GATE U11776 ( .I1(n11566), .I2(n11255), .O(n11561) );
  NAND3_GATE U11777 ( .I1(n11256), .I2(n11562), .I3(n11561), .O(n11551) );
  INV_GATE U11778 ( .I1(n11551), .O(n11548) );
  NAND_GATE U11779 ( .I1(n1413), .I2(A[8]), .O(n11556) );
  NAND_GATE U11780 ( .I1(n11548), .I2(n11556), .O(n11257) );
  NAND_GATE U11781 ( .I1(n11552), .I2(n11257), .O(n11258) );
  INV_GATE U11782 ( .I1(n11556), .O(n11550) );
  NAND_GATE U11783 ( .I1(n11551), .I2(n11550), .O(n11547) );
  NAND_GATE U11784 ( .I1(n11258), .I2(n11547), .O(n11541) );
  NAND_GATE U11785 ( .I1(n11540), .I2(n11541), .O(n11260) );
  NAND_GATE U11786 ( .I1(n1413), .I2(A[9]), .O(n11542) );
  INV_GATE U11787 ( .I1(n11542), .O(n11259) );
  NAND_GATE U11788 ( .I1(n11540), .I2(n11259), .O(n11537) );
  NAND_GATE U11789 ( .I1(n11541), .I2(n11259), .O(n11536) );
  NAND3_GATE U11790 ( .I1(n11260), .I2(n11537), .I3(n11536), .O(n11526) );
  INV_GATE U11791 ( .I1(n11526), .O(n11523) );
  NAND_GATE U11792 ( .I1(n1413), .I2(A[10]), .O(n11531) );
  NAND_GATE U11793 ( .I1(n11523), .I2(n11531), .O(n11261) );
  NAND_GATE U11794 ( .I1(n11527), .I2(n11261), .O(n11262) );
  INV_GATE U11795 ( .I1(n11531), .O(n11525) );
  NAND_GATE U11796 ( .I1(n11526), .I2(n11525), .O(n11522) );
  NAND_GATE U11797 ( .I1(n11262), .I2(n11522), .O(n11517) );
  NAND_GATE U11798 ( .I1(n11516), .I2(n11517), .O(n11264) );
  NAND_GATE U11799 ( .I1(n1413), .I2(A[11]), .O(n11518) );
  INV_GATE U11800 ( .I1(n11518), .O(n11263) );
  NAND_GATE U11801 ( .I1(n11516), .I2(n11263), .O(n11513) );
  NAND_GATE U11802 ( .I1(n11517), .I2(n11263), .O(n11512) );
  NAND3_GATE U11803 ( .I1(n11264), .I2(n11513), .I3(n11512), .O(n11502) );
  INV_GATE U11804 ( .I1(n11502), .O(n11499) );
  NAND_GATE U11805 ( .I1(n1413), .I2(A[12]), .O(n11507) );
  NAND_GATE U11806 ( .I1(n11499), .I2(n11507), .O(n11265) );
  NAND_GATE U11807 ( .I1(n11503), .I2(n11265), .O(n11266) );
  INV_GATE U11808 ( .I1(n11507), .O(n11501) );
  NAND_GATE U11809 ( .I1(n11502), .I2(n11501), .O(n11498) );
  NAND_GATE U11810 ( .I1(n11266), .I2(n11498), .O(n11493) );
  NAND_GATE U11811 ( .I1(n11492), .I2(n11493), .O(n11268) );
  NAND_GATE U11812 ( .I1(n1413), .I2(A[13]), .O(n11494) );
  INV_GATE U11813 ( .I1(n11494), .O(n11267) );
  NAND_GATE U11814 ( .I1(n11492), .I2(n11267), .O(n11489) );
  NAND_GATE U11815 ( .I1(n11493), .I2(n11267), .O(n11488) );
  NAND_GATE U11816 ( .I1(n11477), .I2(n11479), .O(n11475) );
  OR_GATE U11817 ( .I1(n11269), .I2(n11273), .O(n11272) );
  OR_GATE U11818 ( .I1(n11274), .I2(n11270), .O(n11271) );
  NAND_GATE U11819 ( .I1(n11273), .I2(n1034), .O(n11277) );
  NAND3_GATE U11820 ( .I1(n11277), .I2(n11276), .I3(n11275), .O(n11278) );
  INV_GATE U11821 ( .I1(n11476), .O(n11478) );
  NAND_GATE U11822 ( .I1(n11483), .I2(n751), .O(n11279) );
  NAND_GATE U11823 ( .I1(n11478), .I2(n11279), .O(n11280) );
  NAND_GATE U11824 ( .I1(n11475), .I2(n11280), .O(n11675) );
  NAND_GATE U11825 ( .I1(n11674), .I2(n11675), .O(n11282) );
  NAND_GATE U11826 ( .I1(n11281), .I2(n11675), .O(n11670) );
  NAND3_GATE U11827 ( .I1(n11671), .I2(n11282), .I3(n11670), .O(n11687) );
  NAND_GATE U11828 ( .I1(n11685), .I2(n11687), .O(n11682) );
  OR_GATE U11829 ( .I1(n11283), .I2(n11287), .O(n11286) );
  OR_GATE U11830 ( .I1(n11288), .I2(n11284), .O(n11285) );
  NAND_GATE U11831 ( .I1(n11287), .I2(n1001), .O(n11291) );
  NAND3_GATE U11832 ( .I1(n11291), .I2(n11290), .I3(n11289), .O(n11292) );
  INV_GATE U11833 ( .I1(n11683), .O(n11686) );
  INV_GATE U11834 ( .I1(n11687), .O(n11684) );
  NAND_GATE U11835 ( .I1(n11686), .I2(n11293), .O(n11294) );
  NAND_GATE U11836 ( .I1(n11682), .I2(n11294), .O(n11470) );
  OR_GATE U11837 ( .I1(n11299), .I2(n11295), .O(n11305) );
  NAND_GATE U11838 ( .I1(n11296), .I2(n11300), .O(n11304) );
  NAND_GATE U11839 ( .I1(n11298), .I2(n11297), .O(n11301) );
  NAND_GATE U11840 ( .I1(n35), .I2(n11299), .O(n11300) );
  NAND_GATE U11841 ( .I1(n11301), .I2(n11300), .O(n11302) );
  NAND_GATE U11842 ( .I1(n11470), .I2(n11469), .O(n11307) );
  NAND_GATE U11843 ( .I1(n11306), .I2(n11469), .O(n11465) );
  NAND3_GATE U11844 ( .I1(n11466), .I2(n11307), .I3(n11465), .O(n11705) );
  NAND_GATE U11845 ( .I1(n11704), .I2(n11707), .O(n11308) );
  NAND_GATE U11846 ( .I1(n11705), .I2(n11308), .O(n11309) );
  NAND_GATE U11847 ( .I1(n11699), .I2(n11309), .O(n11456) );
  NAND_GATE U11848 ( .I1(n11320), .I2(n11456), .O(n11453) );
  NAND_GATE U11849 ( .I1(n11314), .I2(n11313), .O(n11311) );
  NAND3_GATE U11850 ( .I1(n11312), .I2(n11311), .I3(n11315), .O(n11319) );
  NAND_GATE U11851 ( .I1(n11315), .I2(n11311), .O(n11316) );
  NAND_GATE U11852 ( .I1(n11317), .I2(n11316), .O(n11318) );
  NAND_GATE U11853 ( .I1(n11319), .I2(n11318), .O(n11455) );
  NAND_GATE U11854 ( .I1(n11456), .I2(n11457), .O(n11321) );
  NAND_GATE U11855 ( .I1(n11320), .I2(n11457), .O(n11452) );
  NAND_GATE U11856 ( .I1(n1413), .I2(A[20]), .O(n11920) );
  OR_GATE U11857 ( .I1(n11322), .I2(n11327), .O(n11335) );
  NAND_GATE U11858 ( .I1(n1021), .I2(n11332), .O(n11329) );
  NAND3_GATE U11859 ( .I1(n11330), .I2(n11329), .I3(n11328), .O(n11334) );
  OR_GATE U11860 ( .I1(n11332), .I2(n11331), .O(n11333) );
  NAND3_GATE U11861 ( .I1(n11335), .I2(n11334), .I3(n11333), .O(n11720) );
  NAND_GATE U11862 ( .I1(n11920), .I2(n11720), .O(n11336) );
  NAND_GATE U11863 ( .I1(n11719), .I2(n11336), .O(n11338) );
  INV_GATE U11864 ( .I1(n11920), .O(n11717) );
  INV_GATE U11865 ( .I1(n11720), .O(n11718) );
  NAND_GATE U11866 ( .I1(n11717), .I2(n11718), .O(n11337) );
  NAND_GATE U11867 ( .I1(n11338), .I2(n11337), .O(n11442) );
  INV_GATE U11868 ( .I1(n11347), .O(n11341) );
  NAND_GATE U11869 ( .I1(n11342), .I2(n11341), .O(n11339) );
  NAND_GATE U11870 ( .I1(n11340), .I2(n11339), .O(n11345) );
  NAND_GATE U11871 ( .I1(n11345), .I2(n11344), .O(n11350) );
  INV_GATE U11872 ( .I1(n11346), .O(n11348) );
  NAND_GATE U11873 ( .I1(n11348), .I2(n11347), .O(n11349) );
  NAND_GATE U11874 ( .I1(n11350), .I2(n11349), .O(n11448) );
  NAND_GATE U11875 ( .I1(n11442), .I2(n11448), .O(n11352) );
  NAND_GATE U11876 ( .I1(n11446), .I2(n11448), .O(n11351) );
  NAND3_GATE U11877 ( .I1(n11447), .I2(n11352), .I3(n11351), .O(n11730) );
  NAND_GATE U11878 ( .I1(n11729), .I2(n11890), .O(n11353) );
  NAND_GATE U11879 ( .I1(n11730), .I2(n11353), .O(n11354) );
  NAND_GATE U11880 ( .I1(n11726), .I2(n11354), .O(n11431) );
  NAND_GATE U11881 ( .I1(n11365), .I2(n11431), .O(n11435) );
  INV_GATE U11882 ( .I1(n11362), .O(n11356) );
  NAND3_GATE U11883 ( .I1(n11357), .I2(n11356), .I3(n11355), .O(n11360) );
  NAND_GATE U11884 ( .I1(n11358), .I2(n11362), .O(n11359) );
  NAND3_GATE U11885 ( .I1(n11361), .I2(n11360), .I3(n11359), .O(n11364) );
  NAND_GATE U11886 ( .I1(n1275), .I2(n11362), .O(n11363) );
  NAND_GATE U11887 ( .I1(n11364), .I2(n11363), .O(n11436) );
  NAND_GATE U11888 ( .I1(n11431), .I2(n11436), .O(n11366) );
  NAND_GATE U11889 ( .I1(n11365), .I2(n11436), .O(n11439) );
  NAND3_GATE U11890 ( .I1(n11435), .I2(n11366), .I3(n11439), .O(n11747) );
  NAND_GATE U11891 ( .I1(n11751), .I2(n11749), .O(n11367) );
  NAND_GATE U11892 ( .I1(n11747), .I2(n11367), .O(n11368) );
  NAND_GATE U11893 ( .I1(n11422), .I2(n11423), .O(n11419) );
  NAND_GATE U11894 ( .I1(n11375), .I2(n1389), .O(n11369) );
  NAND_GATE U11895 ( .I1(n11377), .I2(n11369), .O(n11370) );
  NAND_GATE U11896 ( .I1(n11374), .I2(n11370), .O(n11420) );
  NAND_GATE U11897 ( .I1(n11371), .I2(n11369), .O(n11378) );
  INV_GATE U11898 ( .I1(n11378), .O(n11373) );
  NAND_GATE U11899 ( .I1(n11373), .I2(n11380), .O(n11421) );
  NAND3_GATE U11900 ( .I1(n11420), .I2(n11422), .I3(n11421), .O(n11382) );
  NAND_GATE U11901 ( .I1(n392), .I2(n287), .O(n11377) );
  NAND3_GATE U11902 ( .I1(n11375), .I2(n1389), .I3(n11374), .O(n11376) );
  NAND3_GATE U11903 ( .I1(n11378), .I2(n11377), .I3(n11376), .O(n11379) );
  NAND_GATE U11904 ( .I1(n11380), .I2(n11379), .O(n11424) );
  NAND_GATE U11905 ( .I1(n11423), .I2(n11424), .O(n11381) );
  NAND_GATE U11906 ( .I1(n11850), .I2(n11851), .O(n11383) );
  NAND_GATE U11907 ( .I1(n11768), .I2(n11836), .O(n11403) );
  AND_GATE U11908 ( .I1(n11390), .I2(n11384), .O(n11389) );
  NAND_GATE U11909 ( .I1(n11387), .I2(n11386), .O(n11388) );
  NAND3_GATE U11910 ( .I1(n11389), .I2(n11388), .I3(n11394), .O(n11400) );
  INV_GATE U11911 ( .I1(n11394), .O(n11391) );
  NAND4_GATE U11912 ( .I1(n11392), .I2(n11386), .I3(n11390), .I4(n11391), .O(
        n11399) );
  NAND3_GATE U11913 ( .I1(n11392), .I2(n11386), .I3(n11391), .O(n11396) );
  NAND_GATE U11914 ( .I1(n11392), .I2(n11386), .O(n11393) );
  NAND_GATE U11915 ( .I1(n11394), .I2(n11393), .O(n11395) );
  NAND3_GATE U11916 ( .I1(n11397), .I2(n11396), .I3(n11395), .O(n11398) );
  NAND4_GATE U11917 ( .I1(n11400), .I2(n11399), .I3(n11398), .I4(n11836), .O(
        n11402) );
  NAND3_GATE U11918 ( .I1(n11400), .I2(n11399), .I3(n11398), .O(n11835) );
  NAND_GATE U11919 ( .I1(n11768), .I2(n715), .O(n11401) );
  NAND3_GATE U11920 ( .I1(n11403), .I2(n11402), .I3(n11401), .O(n11777) );
  NAND_GATE U11921 ( .I1(n11827), .I2(n11776), .O(n11404) );
  NAND_GATE U11922 ( .I1(n11777), .I2(n11404), .O(n11405) );
  NAND_GATE U11923 ( .I1(n11406), .I2(n11405), .O(n11417) );
  NAND_GATE U11924 ( .I1(n11416), .I2(n11809), .O(n11407) );
  NAND_GATE U11925 ( .I1(n11417), .I2(n11407), .O(n11408) );
  NAND_GATE U11926 ( .I1(n11790), .I2(n11789), .O(n11410) );
  NAND_GATE U11927 ( .I1(n11411), .I2(n1390), .O(n11412) );
  NAND_GATE U11928 ( .I1(n11413), .I2(n11412), .O(\A1[37] ) );
  INV_GATE U11929 ( .I1(n11417), .O(n11415) );
  NAND_GATE U11930 ( .I1(n11416), .I2(n11415), .O(n11806) );
  NAND3_GATE U11931 ( .I1(n11807), .I2(n11417), .I3(n781), .O(n11811) );
  NAND3_GATE U11932 ( .I1(n11806), .I2(n11811), .I3(n11807), .O(n11800) );
  NAND_GATE U11933 ( .I1(n781), .I2(n11417), .O(n11418) );
  NAND_GATE U11934 ( .I1(n11806), .I2(n11418), .O(n11808) );
  NAND_GATE U11935 ( .I1(B[6]), .I2(A[29]), .O(n11825) );
  INV_GATE U11936 ( .I1(n11825), .O(n11831) );
  NAND_GATE U11937 ( .I1(B[6]), .I2(A[28]), .O(n12650) );
  INV_GATE U11938 ( .I1(n12650), .O(n11769) );
  NAND_GATE U11939 ( .I1(B[6]), .I2(A[26]), .O(n12273) );
  INV_GATE U11940 ( .I1(n12273), .O(n11867) );
  OR_GATE U11941 ( .I1(n11424), .I2(n11419), .O(n11430) );
  NAND4_GATE U11942 ( .I1(n11422), .I2(n647), .I3(n11421), .I4(n11420), .O(
        n11429) );
  NAND_GATE U11943 ( .I1(n647), .I2(n11424), .O(n11425) );
  NAND3_GATE U11944 ( .I1(n11427), .I2(n11426), .I3(n11425), .O(n11428) );
  NAND3_GATE U11945 ( .I1(n11430), .I2(n11429), .I3(n11428), .O(n11870) );
  NAND_GATE U11946 ( .I1(n11867), .I2(n390), .O(n11868) );
  NAND_GATE U11947 ( .I1(B[6]), .I2(A[25]), .O(n11882) );
  INV_GATE U11948 ( .I1(n11882), .O(n11877) );
  NAND_GATE U11949 ( .I1(B[6]), .I2(A[24]), .O(n12607) );
  INV_GATE U11950 ( .I1(n11431), .O(n11440) );
  NAND_GATE U11951 ( .I1(n11440), .I2(n11436), .O(n11432) );
  NAND3_GATE U11952 ( .I1(n11434), .I2(n11433), .I3(n11432), .O(n11438) );
  OR_GATE U11953 ( .I1(n11436), .I2(n11435), .O(n11437) );
  NAND_GATE U11954 ( .I1(n11438), .I2(n11437), .O(n11738) );
  NAND_GATE U11955 ( .I1(n12607), .I2(n11738), .O(n11737) );
  INV_GATE U11956 ( .I1(n11739), .O(n11441) );
  NAND_GATE U11957 ( .I1(n11441), .I2(n12607), .O(n11736) );
  NAND_GATE U11958 ( .I1(B[6]), .I2(A[23]), .O(n11904) );
  INV_GATE U11959 ( .I1(n11904), .O(n11896) );
  NAND_GATE U11960 ( .I1(B[6]), .I2(A[22]), .O(n11905) );
  NAND_GATE U11961 ( .I1(n77), .I2(n11448), .O(n11443) );
  NAND3_GATE U11962 ( .I1(n11445), .I2(n11444), .I3(n11443), .O(n11451) );
  NAND3_GATE U11963 ( .I1(n77), .I2(n11446), .I3(n11448), .O(n11450) );
  OR_GATE U11964 ( .I1(n11448), .I2(n11447), .O(n11449) );
  NAND3_GATE U11965 ( .I1(n11451), .I2(n11450), .I3(n11449), .O(n11907) );
  NAND_GATE U11966 ( .I1(B[6]), .I2(A[21]), .O(n11925) );
  INV_GATE U11967 ( .I1(n11925), .O(n11721) );
  OR_GATE U11968 ( .I1(n11452), .I2(n11456), .O(n11464) );
  INV_GATE U11969 ( .I1(n11453), .O(n11454) );
  NAND_GATE U11970 ( .I1(n11454), .I2(n11455), .O(n11463) );
  NAND_GATE U11971 ( .I1(n11456), .I2(n11455), .O(n11460) );
  INV_GATE U11972 ( .I1(n11456), .O(n11458) );
  NAND_GATE U11973 ( .I1(n11458), .I2(n11457), .O(n11459) );
  NAND3_GATE U11974 ( .I1(n11461), .I2(n11460), .I3(n11459), .O(n11462) );
  NAND3_GATE U11975 ( .I1(n11464), .I2(n11463), .I3(n11462), .O(n12198) );
  NAND_GATE U11976 ( .I1(B[6]), .I2(A[20]), .O(n12201) );
  NAND_GATE U11977 ( .I1(n84), .I2(n434), .O(n12196) );
  NAND_GATE U11978 ( .I1(B[6]), .I2(A[19]), .O(n11937) );
  INV_GATE U11979 ( .I1(n11937), .O(n11712) );
  OR_GATE U11980 ( .I1(n11465), .I2(n11470), .O(n11468) );
  OR_GATE U11981 ( .I1(n11469), .I2(n11466), .O(n11467) );
  NAND_GATE U11982 ( .I1(n110), .I2(n11469), .O(n11473) );
  NAND3_GATE U11983 ( .I1(n11473), .I2(n11472), .I3(n11471), .O(n11474) );
  INV_GATE U11984 ( .I1(n12182), .O(n12184) );
  NAND_GATE U11985 ( .I1(B[6]), .I2(A[18]), .O(n12187) );
  INV_GATE U11986 ( .I1(n12187), .O(n12180) );
  NAND_GATE U11987 ( .I1(n12184), .I2(n12180), .O(n12177) );
  NAND_GATE U11988 ( .I1(B[6]), .I2(A[17]), .O(n11947) );
  INV_GATE U11989 ( .I1(n11947), .O(n11695) );
  NAND_GATE U11990 ( .I1(B[6]), .I2(A[16]), .O(n11960) );
  INV_GATE U11991 ( .I1(n11960), .O(n11954) );
  OR_GATE U11992 ( .I1(n11476), .I2(n11475), .O(n11487) );
  NAND_GATE U11993 ( .I1(n751), .I2(n11476), .O(n11481) );
  NAND_GATE U11994 ( .I1(n11477), .I2(n11481), .O(n11485) );
  NAND_GATE U11995 ( .I1(n11479), .I2(n11478), .O(n11480) );
  NAND_GATE U11996 ( .I1(n11481), .I2(n11480), .O(n11482) );
  NAND_GATE U11997 ( .I1(n11483), .I2(n11482), .O(n11484) );
  NAND_GATE U11998 ( .I1(n11485), .I2(n11484), .O(n11486) );
  NAND_GATE U11999 ( .I1(n11487), .I2(n11486), .O(n11967) );
  OR_GATE U12000 ( .I1(n11488), .I2(n11492), .O(n11491) );
  OR_GATE U12001 ( .I1(n11489), .I2(n11493), .O(n11490) );
  NAND_GATE U12002 ( .I1(n11492), .I2(n1039), .O(n11496) );
  NAND3_GATE U12003 ( .I1(n11496), .I2(n11495), .I3(n11494), .O(n11497) );
  INV_GATE U12004 ( .I1(n11976), .O(n11979) );
  OR_GATE U12005 ( .I1(n11498), .I2(n11500), .O(n11511) );
  NAND_GATE U12006 ( .I1(n11500), .I2(n11499), .O(n11505) );
  NAND_GATE U12007 ( .I1(n11501), .I2(n11505), .O(n11509) );
  NAND_GATE U12008 ( .I1(n11503), .I2(n11502), .O(n11504) );
  NAND_GATE U12009 ( .I1(n11505), .I2(n11504), .O(n11506) );
  NAND_GATE U12010 ( .I1(n11507), .I2(n11506), .O(n11508) );
  NAND_GATE U12011 ( .I1(n11509), .I2(n11508), .O(n11510) );
  NAND_GATE U12012 ( .I1(n11511), .I2(n11510), .O(n11992) );
  OR_GATE U12013 ( .I1(n11512), .I2(n11516), .O(n11515) );
  OR_GATE U12014 ( .I1(n11513), .I2(n11517), .O(n11514) );
  NAND_GATE U12015 ( .I1(n11516), .I2(n1060), .O(n11520) );
  NAND3_GATE U12016 ( .I1(n11520), .I2(n11519), .I3(n11518), .O(n11521) );
  INV_GATE U12017 ( .I1(n12000), .O(n12003) );
  OR_GATE U12018 ( .I1(n11522), .I2(n11524), .O(n11535) );
  NAND_GATE U12019 ( .I1(n11524), .I2(n11523), .O(n11529) );
  NAND_GATE U12020 ( .I1(n11525), .I2(n11529), .O(n11533) );
  NAND_GATE U12021 ( .I1(n11527), .I2(n11526), .O(n11528) );
  NAND_GATE U12022 ( .I1(n11529), .I2(n11528), .O(n11530) );
  NAND_GATE U12023 ( .I1(n11531), .I2(n11530), .O(n11532) );
  NAND_GATE U12024 ( .I1(n11533), .I2(n11532), .O(n11534) );
  NAND_GATE U12025 ( .I1(n11535), .I2(n11534), .O(n12016) );
  OR_GATE U12026 ( .I1(n11536), .I2(n11540), .O(n11539) );
  OR_GATE U12027 ( .I1(n11537), .I2(n11541), .O(n11538) );
  AND_GATE U12028 ( .I1(n11539), .I2(n11538), .O(n11546) );
  NAND_GATE U12029 ( .I1(n11540), .I2(n1070), .O(n11544) );
  NAND3_GATE U12030 ( .I1(n11544), .I2(n11543), .I3(n11542), .O(n11545) );
  NAND_GATE U12031 ( .I1(n11546), .I2(n11545), .O(n12025) );
  INV_GATE U12032 ( .I1(n12025), .O(n12028) );
  OR_GATE U12033 ( .I1(n11547), .I2(n11549), .O(n11560) );
  NAND_GATE U12034 ( .I1(n11549), .I2(n11548), .O(n11554) );
  NAND_GATE U12035 ( .I1(n11550), .I2(n11554), .O(n11558) );
  NAND_GATE U12036 ( .I1(n11552), .I2(n11551), .O(n11553) );
  NAND_GATE U12037 ( .I1(n11554), .I2(n11553), .O(n11555) );
  NAND_GATE U12038 ( .I1(n11556), .I2(n11555), .O(n11557) );
  NAND_GATE U12039 ( .I1(n11558), .I2(n11557), .O(n11559) );
  NAND_GATE U12040 ( .I1(n11560), .I2(n11559), .O(n12041) );
  OR_GATE U12041 ( .I1(n11561), .I2(n11565), .O(n11564) );
  OR_GATE U12042 ( .I1(n11562), .I2(n11566), .O(n11563) );
  AND_GATE U12043 ( .I1(n11564), .I2(n11563), .O(n11571) );
  NAND_GATE U12044 ( .I1(n11565), .I2(n1080), .O(n11569) );
  NAND3_GATE U12045 ( .I1(n11569), .I2(n11568), .I3(n11567), .O(n11570) );
  NAND_GATE U12046 ( .I1(n11571), .I2(n11570), .O(n12050) );
  INV_GATE U12047 ( .I1(n12050), .O(n12053) );
  OR_GATE U12048 ( .I1(n11572), .I2(n11574), .O(n11585) );
  NAND_GATE U12049 ( .I1(n11574), .I2(n11573), .O(n11579) );
  NAND_GATE U12050 ( .I1(n11575), .I2(n11579), .O(n11583) );
  NAND_GATE U12051 ( .I1(n11577), .I2(n11576), .O(n11578) );
  NAND_GATE U12052 ( .I1(n11579), .I2(n11578), .O(n11580) );
  NAND_GATE U12053 ( .I1(n11581), .I2(n11580), .O(n11582) );
  NAND_GATE U12054 ( .I1(n11583), .I2(n11582), .O(n11584) );
  NAND_GATE U12055 ( .I1(n11585), .I2(n11584), .O(n12066) );
  OR_GATE U12056 ( .I1(n11586), .I2(n11590), .O(n11589) );
  OR_GATE U12057 ( .I1(n11587), .I2(n11591), .O(n11588) );
  AND_GATE U12058 ( .I1(n11589), .I2(n11588), .O(n11596) );
  NAND_GATE U12059 ( .I1(n11590), .I2(n1186), .O(n11594) );
  NAND3_GATE U12060 ( .I1(n11594), .I2(n11593), .I3(n11592), .O(n11595) );
  NAND_GATE U12061 ( .I1(n11596), .I2(n11595), .O(n12075) );
  INV_GATE U12062 ( .I1(n12075), .O(n12078) );
  OR_GATE U12063 ( .I1(n11597), .I2(n11599), .O(n11610) );
  NAND_GATE U12064 ( .I1(n11599), .I2(n11598), .O(n11604) );
  NAND_GATE U12065 ( .I1(n11600), .I2(n11604), .O(n11608) );
  NAND_GATE U12066 ( .I1(n11602), .I2(n11601), .O(n11603) );
  NAND_GATE U12067 ( .I1(n11604), .I2(n11603), .O(n11605) );
  NAND_GATE U12068 ( .I1(n11606), .I2(n11605), .O(n11607) );
  NAND_GATE U12069 ( .I1(n11608), .I2(n11607), .O(n11609) );
  NAND_GATE U12070 ( .I1(n11610), .I2(n11609), .O(n12091) );
  OR_GATE U12071 ( .I1(n11611), .I2(n11615), .O(n11614) );
  OR_GATE U12072 ( .I1(n11612), .I2(n11616), .O(n11613) );
  AND_GATE U12073 ( .I1(n11614), .I2(n11613), .O(n11621) );
  NAND_GATE U12074 ( .I1(n11615), .I2(n1245), .O(n11619) );
  NAND3_GATE U12075 ( .I1(n11619), .I2(n11618), .I3(n11617), .O(n11620) );
  NAND_GATE U12076 ( .I1(n11621), .I2(n11620), .O(n12100) );
  INV_GATE U12077 ( .I1(n12100), .O(n12103) );
  INV_GATE U12078 ( .I1(n11622), .O(n11623) );
  NAND_GATE U12079 ( .I1(n11627), .I2(n11623), .O(n11635) );
  NAND_GATE U12080 ( .I1(n11625), .I2(n11629), .O(n11633) );
  NAND_GATE U12081 ( .I1(n11627), .I2(n11626), .O(n11628) );
  NAND_GATE U12082 ( .I1(n11629), .I2(n11628), .O(n11630) );
  NAND_GATE U12083 ( .I1(n11631), .I2(n11630), .O(n11632) );
  NAND_GATE U12084 ( .I1(n11633), .I2(n11632), .O(n11634) );
  NAND_GATE U12085 ( .I1(n11635), .I2(n11634), .O(n12116) );
  NAND_GATE U12086 ( .I1(n1414), .I2(A[0]), .O(n11636) );
  NAND_GATE U12087 ( .I1(n14241), .I2(n11636), .O(n11637) );
  NAND_GATE U12088 ( .I1(n1415), .I2(n11637), .O(n11641) );
  NAND_GATE U12089 ( .I1(n1417), .I2(A[1]), .O(n11638) );
  NAND_GATE U12090 ( .I1(n724), .I2(n11638), .O(n11639) );
  NAND_GATE U12091 ( .I1(n1413), .I2(n11639), .O(n11640) );
  NAND_GATE U12092 ( .I1(n11641), .I2(n11640), .O(n12128) );
  NAND_GATE U12093 ( .I1(B[6]), .I2(A[2]), .O(n12132) );
  NAND3_GATE U12094 ( .I1(B[6]), .I2(n1413), .I3(n1254), .O(n12125) );
  NAND_GATE U12095 ( .I1(n12132), .I2(n12125), .O(n11642) );
  NAND_GATE U12096 ( .I1(n12128), .I2(n11642), .O(n11643) );
  INV_GATE U12097 ( .I1(n12132), .O(n12126) );
  INV_GATE U12098 ( .I1(n12125), .O(n12127) );
  NAND_GATE U12099 ( .I1(n12126), .I2(n12127), .O(n12123) );
  NAND_GATE U12100 ( .I1(n11643), .I2(n12123), .O(n12117) );
  NAND_GATE U12101 ( .I1(n12116), .I2(n12117), .O(n11645) );
  NAND_GATE U12102 ( .I1(B[6]), .I2(A[3]), .O(n12118) );
  INV_GATE U12103 ( .I1(n12118), .O(n11644) );
  NAND_GATE U12104 ( .I1(n12116), .I2(n11644), .O(n12113) );
  NAND_GATE U12105 ( .I1(n12117), .I2(n11644), .O(n12112) );
  NAND3_GATE U12106 ( .I1(n11645), .I2(n12113), .I3(n12112), .O(n12102) );
  INV_GATE U12107 ( .I1(n12102), .O(n12099) );
  NAND_GATE U12108 ( .I1(B[6]), .I2(A[4]), .O(n12107) );
  NAND_GATE U12109 ( .I1(n12099), .I2(n12107), .O(n11646) );
  NAND_GATE U12110 ( .I1(n12103), .I2(n11646), .O(n11647) );
  INV_GATE U12111 ( .I1(n12107), .O(n12101) );
  NAND_GATE U12112 ( .I1(n12102), .I2(n12101), .O(n12098) );
  NAND_GATE U12113 ( .I1(n11647), .I2(n12098), .O(n12092) );
  NAND_GATE U12114 ( .I1(n12091), .I2(n12092), .O(n11649) );
  NAND_GATE U12115 ( .I1(B[6]), .I2(A[5]), .O(n12093) );
  INV_GATE U12116 ( .I1(n12093), .O(n11648) );
  NAND_GATE U12117 ( .I1(n12091), .I2(n11648), .O(n12088) );
  NAND_GATE U12118 ( .I1(n12092), .I2(n11648), .O(n12087) );
  NAND3_GATE U12119 ( .I1(n11649), .I2(n12088), .I3(n12087), .O(n12077) );
  INV_GATE U12120 ( .I1(n12077), .O(n12074) );
  NAND_GATE U12121 ( .I1(B[6]), .I2(A[6]), .O(n12082) );
  NAND_GATE U12122 ( .I1(n12074), .I2(n12082), .O(n11650) );
  NAND_GATE U12123 ( .I1(n12078), .I2(n11650), .O(n11651) );
  INV_GATE U12124 ( .I1(n12082), .O(n12076) );
  NAND_GATE U12125 ( .I1(n12077), .I2(n12076), .O(n12073) );
  NAND_GATE U12126 ( .I1(n11651), .I2(n12073), .O(n12067) );
  NAND_GATE U12127 ( .I1(n12066), .I2(n12067), .O(n11653) );
  NAND_GATE U12128 ( .I1(B[6]), .I2(A[7]), .O(n12068) );
  INV_GATE U12129 ( .I1(n12068), .O(n11652) );
  NAND_GATE U12130 ( .I1(n12066), .I2(n11652), .O(n12063) );
  NAND_GATE U12131 ( .I1(n12067), .I2(n11652), .O(n12062) );
  NAND3_GATE U12132 ( .I1(n11653), .I2(n12063), .I3(n12062), .O(n12052) );
  INV_GATE U12133 ( .I1(n12052), .O(n12049) );
  NAND_GATE U12134 ( .I1(B[6]), .I2(A[8]), .O(n12057) );
  NAND_GATE U12135 ( .I1(n12049), .I2(n12057), .O(n11654) );
  NAND_GATE U12136 ( .I1(n12053), .I2(n11654), .O(n11655) );
  INV_GATE U12137 ( .I1(n12057), .O(n12051) );
  NAND_GATE U12138 ( .I1(n12052), .I2(n12051), .O(n12048) );
  NAND_GATE U12139 ( .I1(n11655), .I2(n12048), .O(n12042) );
  NAND_GATE U12140 ( .I1(n12041), .I2(n12042), .O(n11657) );
  NAND_GATE U12141 ( .I1(B[6]), .I2(A[9]), .O(n12043) );
  INV_GATE U12142 ( .I1(n12043), .O(n11656) );
  NAND_GATE U12143 ( .I1(n12041), .I2(n11656), .O(n12038) );
  NAND_GATE U12144 ( .I1(n12042), .I2(n11656), .O(n12037) );
  NAND3_GATE U12145 ( .I1(n11657), .I2(n12038), .I3(n12037), .O(n12027) );
  INV_GATE U12146 ( .I1(n12027), .O(n12024) );
  NAND_GATE U12147 ( .I1(B[6]), .I2(A[10]), .O(n12032) );
  NAND_GATE U12148 ( .I1(n12024), .I2(n12032), .O(n11658) );
  NAND_GATE U12149 ( .I1(n12028), .I2(n11658), .O(n11659) );
  INV_GATE U12150 ( .I1(n12032), .O(n12026) );
  NAND_GATE U12151 ( .I1(n12027), .I2(n12026), .O(n12023) );
  NAND_GATE U12152 ( .I1(n11659), .I2(n12023), .O(n12017) );
  NAND_GATE U12153 ( .I1(n12016), .I2(n12017), .O(n11661) );
  NAND_GATE U12154 ( .I1(B[6]), .I2(A[11]), .O(n12018) );
  INV_GATE U12155 ( .I1(n12018), .O(n11660) );
  NAND_GATE U12156 ( .I1(n12016), .I2(n11660), .O(n12013) );
  NAND_GATE U12157 ( .I1(n12017), .I2(n11660), .O(n12012) );
  NAND3_GATE U12158 ( .I1(n11661), .I2(n12013), .I3(n12012), .O(n12002) );
  INV_GATE U12159 ( .I1(n12002), .O(n11999) );
  NAND_GATE U12160 ( .I1(B[6]), .I2(A[12]), .O(n12007) );
  NAND_GATE U12161 ( .I1(n11999), .I2(n12007), .O(n11662) );
  NAND_GATE U12162 ( .I1(n12003), .I2(n11662), .O(n11663) );
  INV_GATE U12163 ( .I1(n12007), .O(n12001) );
  NAND_GATE U12164 ( .I1(n12002), .I2(n12001), .O(n11998) );
  NAND_GATE U12165 ( .I1(n11663), .I2(n11998), .O(n11993) );
  NAND_GATE U12166 ( .I1(n11992), .I2(n11993), .O(n11665) );
  NAND_GATE U12167 ( .I1(B[6]), .I2(A[13]), .O(n11994) );
  INV_GATE U12168 ( .I1(n11994), .O(n11664) );
  NAND_GATE U12169 ( .I1(n11992), .I2(n11664), .O(n11989) );
  NAND_GATE U12170 ( .I1(n11993), .I2(n11664), .O(n11988) );
  NAND3_GATE U12171 ( .I1(n11665), .I2(n11989), .I3(n11988), .O(n11978) );
  INV_GATE U12172 ( .I1(n11978), .O(n11975) );
  NAND_GATE U12173 ( .I1(B[6]), .I2(A[14]), .O(n11983) );
  NAND_GATE U12174 ( .I1(n11975), .I2(n11983), .O(n11666) );
  NAND_GATE U12175 ( .I1(n11979), .I2(n11666), .O(n11667) );
  INV_GATE U12176 ( .I1(n11983), .O(n11977) );
  NAND_GATE U12177 ( .I1(n11978), .I2(n11977), .O(n11974) );
  NAND_GATE U12178 ( .I1(n11667), .I2(n11974), .O(n11968) );
  NAND_GATE U12179 ( .I1(n11967), .I2(n11968), .O(n11669) );
  NAND_GATE U12180 ( .I1(B[6]), .I2(A[15]), .O(n11969) );
  INV_GATE U12181 ( .I1(n11969), .O(n11668) );
  NAND_GATE U12182 ( .I1(n11968), .I2(n11668), .O(n11963) );
  NAND3_GATE U12183 ( .I1(n11669), .I2(n11964), .I3(n11963), .O(n11956) );
  NAND_GATE U12184 ( .I1(n11954), .I2(n11956), .O(n11952) );
  OR_GATE U12185 ( .I1(n11670), .I2(n11674), .O(n11673) );
  OR_GATE U12186 ( .I1(n11675), .I2(n11671), .O(n11672) );
  NAND_GATE U12187 ( .I1(n11674), .I2(n1006), .O(n11678) );
  NAND3_GATE U12188 ( .I1(n11678), .I2(n11677), .I3(n11676), .O(n11679) );
  INV_GATE U12189 ( .I1(n11953), .O(n11955) );
  NAND_GATE U12190 ( .I1(n11960), .I2(n771), .O(n11680) );
  NAND_GATE U12191 ( .I1(n11955), .I2(n11680), .O(n11681) );
  NAND_GATE U12192 ( .I1(n11952), .I2(n11681), .O(n11946) );
  NAND_GATE U12193 ( .I1(n11695), .I2(n11946), .O(n11942) );
  OR_GATE U12194 ( .I1(n11683), .I2(n11682), .O(n11694) );
  NAND_GATE U12195 ( .I1(n11684), .I2(n11683), .O(n11689) );
  NAND_GATE U12196 ( .I1(n11685), .I2(n11689), .O(n11693) );
  NAND_GATE U12197 ( .I1(n11687), .I2(n11686), .O(n11688) );
  NAND_GATE U12198 ( .I1(n11689), .I2(n11688), .O(n11690) );
  NAND_GATE U12199 ( .I1(n11691), .I2(n11690), .O(n11692) );
  NAND_GATE U12200 ( .I1(n11946), .I2(n11945), .O(n11696) );
  NAND3_GATE U12201 ( .I1(n11942), .I2(n11696), .I3(n11941), .O(n12183) );
  NAND_GATE U12202 ( .I1(n12182), .I2(n12187), .O(n11697) );
  NAND_GATE U12203 ( .I1(n12183), .I2(n11697), .O(n11698) );
  NAND_GATE U12204 ( .I1(n12177), .I2(n11698), .O(n11936) );
  NAND_GATE U12205 ( .I1(n11712), .I2(n11936), .O(n11932) );
  INV_GATE U12206 ( .I1(n11699), .O(n11700) );
  NAND_GATE U12207 ( .I1(n11700), .I2(n11705), .O(n11711) );
  INV_GATE U12208 ( .I1(n11705), .O(n11703) );
  NAND_GATE U12209 ( .I1(n11704), .I2(n11703), .O(n11701) );
  NAND_GATE U12210 ( .I1(n11702), .I2(n11701), .O(n11709) );
  NAND_GATE U12211 ( .I1(n11709), .I2(n11708), .O(n11710) );
  NAND_GATE U12212 ( .I1(n11711), .I2(n11710), .O(n11935) );
  NAND_GATE U12213 ( .I1(n11936), .I2(n11935), .O(n11713) );
  NAND_GATE U12214 ( .I1(n11712), .I2(n11935), .O(n11931) );
  NAND3_GATE U12215 ( .I1(n11932), .I2(n11713), .I3(n11931), .O(n12199) );
  NAND_GATE U12216 ( .I1(n12198), .I2(n12201), .O(n11714) );
  NAND_GATE U12217 ( .I1(n12199), .I2(n11714), .O(n11715) );
  NAND_GATE U12218 ( .I1(n12196), .I2(n11715), .O(n11926) );
  NAND_GATE U12219 ( .I1(n11721), .I2(n11926), .O(n11916) );
  NAND_GATE U12220 ( .I1(n300), .I2(n11720), .O(n11716) );
  NAND3_GATE U12221 ( .I1(n11718), .I2(n11717), .I3(n11719), .O(n11919) );
  NAND_GATE U12222 ( .I1(n83), .I2(n11919), .O(n11921) );
  NAND3_GATE U12223 ( .I1(n11926), .I2(n11921), .I3(n11914), .O(n11722) );
  NAND3_GATE U12224 ( .I1(n11721), .I2(n11921), .I3(n11914), .O(n11927) );
  NAND3_GATE U12225 ( .I1(n11916), .I2(n11722), .I3(n11927), .O(n11911) );
  NAND_GATE U12226 ( .I1(n11905), .I2(n11907), .O(n11723) );
  NAND_GATE U12227 ( .I1(n11729), .I2(n11728), .O(n11724) );
  NAND_GATE U12228 ( .I1(n11725), .I2(n11724), .O(n11891) );
  INV_GATE U12229 ( .I1(n11891), .O(n11727) );
  NAND_GATE U12230 ( .I1(n11727), .I2(n11894), .O(n11733) );
  NAND3_GATE U12231 ( .I1(n11892), .I2(n11733), .I3(n11732), .O(n11735) );
  NAND3_GATE U12232 ( .I1(n11896), .I2(n11733), .I3(n11732), .O(n11734) );
  NAND3_GATE U12233 ( .I1(n11895), .I2(n11735), .I3(n11734), .O(n11887) );
  NAND3_GATE U12234 ( .I1(n11737), .I2(n11736), .I3(n11887), .O(n11741) );
  INV_GATE U12235 ( .I1(n12607), .O(n11886) );
  NAND_GATE U12236 ( .I1(n11886), .I2(n1395), .O(n11740) );
  NAND_GATE U12237 ( .I1(n11741), .I2(n11740), .O(n11874) );
  NAND_GATE U12238 ( .I1(n11877), .I2(n11874), .O(n11758) );
  NAND_GATE U12239 ( .I1(n11751), .I2(n11750), .O(n11742) );
  NAND_GATE U12240 ( .I1(n11743), .I2(n11742), .O(n11753) );
  NAND_GATE U12241 ( .I1(n756), .I2(n11755), .O(n11876) );
  NAND_GATE U12242 ( .I1(n11748), .I2(n11747), .O(n11745) );
  NAND_GATE U12243 ( .I1(n11745), .I2(n11742), .O(n11746) );
  NAND_GATE U12244 ( .I1(n11749), .I2(n11746), .O(n11875) );
  NAND3_GATE U12245 ( .I1(n11877), .I2(n11876), .I3(n11875), .O(n11757) );
  NAND3_GATE U12246 ( .I1(n11751), .I2(n11750), .I3(n11749), .O(n11752) );
  NAND3_GATE U12247 ( .I1(n11753), .I2(n11745), .I3(n11752), .O(n11754) );
  NAND_GATE U12248 ( .I1(n11755), .I2(n11754), .O(n11873) );
  NAND_GATE U12249 ( .I1(n11874), .I2(n11873), .O(n11756) );
  NAND_GATE U12250 ( .I1(n12273), .I2(n11870), .O(n11759) );
  NAND_GATE U12251 ( .I1(n11869), .I2(n11759), .O(n11760) );
  NAND_GATE U12252 ( .I1(n11868), .I2(n11760), .O(n11858) );
  NAND_GATE U12253 ( .I1(n11851), .I2(n372), .O(n11761) );
  NAND_GATE U12254 ( .I1(n11853), .I2(n11761), .O(n11762) );
  NAND_GATE U12255 ( .I1(n11850), .I2(n11762), .O(n11764) );
  INV_GATE U12256 ( .I1(n11854), .O(n11763) );
  NAND_GATE U12257 ( .I1(n1356), .I2(n11849), .O(n11856) );
  NAND_GATE U12258 ( .I1(n11763), .I2(n11856), .O(n11765) );
  NAND3_GATE U12259 ( .I1(n11858), .I2(n11764), .I3(n11765), .O(n11767) );
  NAND_GATE U12260 ( .I1(B[6]), .I2(A[27]), .O(n11863) );
  INV_GATE U12261 ( .I1(n11863), .O(n11766) );
  NAND3_GATE U12262 ( .I1(n11766), .I2(n11765), .I3(n11764), .O(n11857) );
  NAND_GATE U12263 ( .I1(n11766), .I2(n11858), .O(n11848) );
  NAND3_GATE U12264 ( .I1(n11767), .I2(n11857), .I3(n11848), .O(n11844) );
  NAND_GATE U12265 ( .I1(n11769), .I2(n11844), .O(n11840) );
  NAND_GATE U12266 ( .I1(n11768), .I2(n11770), .O(n11837) );
  NAND_GATE U12267 ( .I1(n655), .I2(n11835), .O(n11770) );
  NAND_GATE U12268 ( .I1(n11838), .I2(n11770), .O(n11841) );
  NAND_GATE U12269 ( .I1(n992), .I2(n11846), .O(n11772) );
  NAND3_GATE U12270 ( .I1(n11844), .I2(n11847), .I3(n11846), .O(n11771) );
  NAND3_GATE U12271 ( .I1(n11840), .I2(n11772), .I3(n11771), .O(n11822) );
  NAND_GATE U12272 ( .I1(n11831), .I2(n11822), .O(n11828) );
  INV_GATE U12273 ( .I1(n11777), .O(n11775) );
  NAND_GATE U12274 ( .I1(n11776), .I2(n11775), .O(n11773) );
  NAND_GATE U12275 ( .I1(n11774), .I2(n11773), .O(n11819) );
  NAND_GATE U12276 ( .I1(n11819), .I2(n11779), .O(n11780) );
  NAND_GATE U12277 ( .I1(n11826), .I2(n11780), .O(n11781) );
  NAND_GATE U12278 ( .I1(n11831), .I2(n11781), .O(n11783) );
  NAND_GATE U12279 ( .I1(n11822), .I2(n11781), .O(n11782) );
  NAND3_GATE U12280 ( .I1(n11828), .I2(n11783), .I3(n11782), .O(n11802) );
  NAND3_GATE U12281 ( .I1(n11800), .I2(n11799), .I3(n11802), .O(n11785) );
  NAND_GATE U12282 ( .I1(B[6]), .I2(A[30]), .O(n11803) );
  INV_GATE U12283 ( .I1(n11803), .O(n11813) );
  NAND3_GATE U12284 ( .I1(n11800), .I2(n11799), .I3(n11813), .O(n11784) );
  NAND_GATE U12285 ( .I1(n11813), .I2(n11802), .O(n11814) );
  AND3_GATE U12286 ( .I1(n11785), .I2(n11784), .I3(n11814), .O(n12234) );
  NAND_GATE U12287 ( .I1(n1412), .I2(A[31]), .O(n12233) );
  NAND3_GATE U12288 ( .I1(n11790), .I2(n911), .I3(n11789), .O(n11791) );
  NAND3_GATE U12289 ( .I1(n11793), .I2(n11792), .I3(n11791), .O(n11795) );
  NAND_GATE U12290 ( .I1(n928), .I2(n357), .O(n11794) );
  NAND_GATE U12291 ( .I1(n11795), .I2(n11794), .O(n12235) );
  NAND_GATE U12292 ( .I1(n12236), .I2(n12235), .O(n12238) );
  NAND_GATE U12293 ( .I1(n11796), .I2(n350), .O(n11797) );
  NAND_GATE U12294 ( .I1(n11798), .I2(n11797), .O(\A1[36] ) );
  INV_GATE U12295 ( .I1(n11802), .O(n11812) );
  NAND_GATE U12296 ( .I1(n11800), .I2(n11799), .O(n11801) );
  NAND_GATE U12297 ( .I1(n11802), .I2(n11801), .O(n11804) );
  NAND3_GATE U12298 ( .I1(n11805), .I2(n11804), .I3(n11803), .O(n11818) );
  NAND_GATE U12299 ( .I1(n11807), .I2(n11806), .O(n11810) );
  NAND3_GATE U12300 ( .I1(n11813), .I2(n11812), .I3(n11815), .O(n11817) );
  OR_GATE U12301 ( .I1(n11815), .I2(n11814), .O(n11816) );
  NAND3_GATE U12302 ( .I1(n11818), .I2(n11817), .I3(n11816), .O(n12643) );
  NAND3_GATE U12303 ( .I1(n11779), .I2(n11820), .I3(n286), .O(n11824) );
  NAND_GATE U12304 ( .I1(n11820), .I2(n11779), .O(n11821) );
  NAND_GATE U12305 ( .I1(n11822), .I2(n11821), .O(n11823) );
  NAND3_GATE U12306 ( .I1(n11825), .I2(n11824), .I3(n11823), .O(n11834) );
  AND_GATE U12307 ( .I1(n11830), .I2(n11779), .O(n11829) );
  OR_GATE U12308 ( .I1(n11829), .I2(n11828), .O(n11833) );
  NAND4_GATE U12309 ( .I1(n11831), .I2(n11830), .I3(n11779), .I4(n286), .O(
        n11832) );
  NAND3_GATE U12310 ( .I1(n11834), .I2(n11833), .I3(n11832), .O(n13082) );
  NAND_GATE U12311 ( .I1(n1410), .I2(A[30]), .O(n13086) );
  INV_GATE U12312 ( .I1(n13086), .O(n12244) );
  NAND_GATE U12313 ( .I1(n716), .I2(n12244), .O(n12232) );
  INV_GATE U12314 ( .I1(n11844), .O(n11845) );
  NAND3_GATE U12315 ( .I1(n11846), .I2(n992), .I3(n11845), .O(n12247) );
  NAND_GATE U12316 ( .I1(n1410), .I2(A[29]), .O(n12250) );
  INV_GATE U12317 ( .I1(n12250), .O(n12655) );
  NAND3_GATE U12318 ( .I1(n11835), .I2(n655), .I3(n11842), .O(n11839) );
  NAND_GATE U12319 ( .I1(n11836), .I2(n715), .O(n11838) );
  NAND_GATE U12320 ( .I1(n11842), .I2(n11841), .O(n11846) );
  NAND_GATE U12321 ( .I1(n11847), .I2(n11846), .O(n11843) );
  NAND_GATE U12322 ( .I1(n11844), .I2(n11843), .O(n12649) );
  NAND3_GATE U12323 ( .I1(n11847), .I2(n11846), .I3(n11845), .O(n12651) );
  NAND3_GATE U12324 ( .I1(n12649), .I2(n12651), .I3(n12650), .O(n12248) );
  NAND4_GATE U12325 ( .I1(n12247), .I2(n12655), .I3(n12246), .I4(n12248), .O(
        n12249) );
  NAND_GATE U12326 ( .I1(n1410), .I2(A[28]), .O(n12258) );
  NAND_GATE U12327 ( .I1(n885), .I2(n11849), .O(n11853) );
  NAND3_GATE U12328 ( .I1(n11851), .I2(n372), .I3(n11850), .O(n11852) );
  NAND3_GATE U12329 ( .I1(n11854), .I2(n11853), .I3(n11852), .O(n11855) );
  NAND_GATE U12330 ( .I1(n11856), .I2(n11855), .O(n11859) );
  INV_GATE U12331 ( .I1(n11858), .O(n11860) );
  NAND_GATE U12332 ( .I1(n11860), .I2(n11859), .O(n11861) );
  NAND3_GATE U12333 ( .I1(n11862), .I2(n11861), .I3(n11863), .O(n12255) );
  NAND4_GATE U12334 ( .I1(n11863), .I2(n11862), .I3(n12258), .I4(n11861), .O(
        n12225) );
  NAND_GATE U12335 ( .I1(n11865), .I2(n11864), .O(n11866) );
  NAND_GATE U12336 ( .I1(n1410), .I2(A[27]), .O(n12279) );
  INV_GATE U12337 ( .I1(n12279), .O(n12221) );
  NAND_GATE U12338 ( .I1(n523), .I2(n12274), .O(n12222) );
  NAND_GATE U12339 ( .I1(n390), .I2(n11869), .O(n11872) );
  NAND_GATE U12340 ( .I1(n11870), .I2(n1278), .O(n11871) );
  NAND_GATE U12341 ( .I1(n11872), .I2(n11871), .O(n12272) );
  NAND3_GATE U12342 ( .I1(n12221), .I2(n12222), .I3(n12266), .O(n12271) );
  NAND_GATE U12343 ( .I1(n1410), .I2(A[26]), .O(n12689) );
  INV_GATE U12344 ( .I1(n12689), .O(n12622) );
  NAND_GATE U12345 ( .I1(n11874), .I2(n495), .O(n11883) );
  AND3_GATE U12346 ( .I1(n11884), .I2(n11882), .I3(n11883), .O(n11880) );
  NAND3_GATE U12347 ( .I1(n11874), .I2(n495), .I3(n11877), .O(n11879) );
  NAND_GATE U12348 ( .I1(n11879), .I2(n11878), .O(n11881) );
  OR_GATE U12349 ( .I1(n11880), .I2(n11881), .O(n12620) );
  NAND_GATE U12350 ( .I1(n12622), .I2(n12623), .O(n12220) );
  NAND_GATE U12351 ( .I1(n12689), .I2(n11881), .O(n12218) );
  NAND4_GATE U12352 ( .I1(n11884), .I2(n11883), .I3(n12689), .I4(n11882), .O(
        n12217) );
  NAND_GATE U12353 ( .I1(n1410), .I2(A[25]), .O(n12606) );
  INV_GATE U12354 ( .I1(n12606), .O(n12612) );
  NAND_GATE U12355 ( .I1(n158), .I2(n11888), .O(n11885) );
  NAND_GATE U12356 ( .I1(n11886), .I2(n11885), .O(n12608) );
  NAND3_GATE U12357 ( .I1(n11887), .I2(n11886), .I3(n1395), .O(n12610) );
  NAND_GATE U12358 ( .I1(n11887), .I2(n1395), .O(n11889) );
  NAND3_GATE U12359 ( .I1(n12612), .I2(n12613), .I3(n12611), .O(n12216) );
  NAND_GATE U12360 ( .I1(n1410), .I2(A[24]), .O(n12716) );
  INV_GATE U12361 ( .I1(n12716), .O(n12283) );
  NAND_GATE U12362 ( .I1(n11891), .I2(n11732), .O(n11893) );
  NAND3_GATE U12363 ( .I1(n11893), .I2(n11894), .I3(n11892), .O(n11903) );
  NAND_GATE U12364 ( .I1(n11894), .I2(n11893), .O(n11897) );
  NAND_GATE U12365 ( .I1(n470), .I2(n11897), .O(n11902) );
  AND3_GATE U12366 ( .I1(n11903), .I2(n11902), .I3(n11904), .O(n11900) );
  OR_GATE U12367 ( .I1(n11897), .I2(n11895), .O(n11899) );
  NAND3_GATE U12368 ( .I1(n470), .I2(n11897), .I3(n11896), .O(n11898) );
  NAND_GATE U12369 ( .I1(n11899), .I2(n11898), .O(n11901) );
  NAND_GATE U12370 ( .I1(n12716), .I2(n11901), .O(n12213) );
  NAND4_GATE U12371 ( .I1(n11904), .I2(n11903), .I3(n12716), .I4(n11902), .O(
        n12212) );
  NAND_GATE U12372 ( .I1(n1410), .I2(A[23]), .O(n12296) );
  INV_GATE U12373 ( .I1(n12296), .O(n12210) );
  INV_GATE U12374 ( .I1(n11911), .O(n11906) );
  NAND3_GATE U12375 ( .I1(n11907), .I2(n11906), .I3(n11905), .O(n11908) );
  NAND3_GATE U12376 ( .I1(n11910), .I2(n11909), .I3(n11908), .O(n11913) );
  NAND_GATE U12377 ( .I1(n1383), .I2(n11911), .O(n11912) );
  NAND_GATE U12378 ( .I1(n11913), .I2(n11912), .O(n12293) );
  NAND_GATE U12379 ( .I1(n12210), .I2(n12293), .O(n12288) );
  NAND_GATE U12380 ( .I1(n11915), .I2(n11914), .O(n11918) );
  INV_GATE U12381 ( .I1(n11916), .O(n11917) );
  NAND3_GATE U12382 ( .I1(n11919), .I2(n11918), .I3(n11917), .O(n11930) );
  NAND_GATE U12383 ( .I1(n11921), .I2(n11914), .O(n11922) );
  NAND_GATE U12384 ( .I1(n11926), .I2(n11922), .O(n11924) );
  OR_GATE U12385 ( .I1(n11922), .I2(n11926), .O(n11923) );
  NAND3_GATE U12386 ( .I1(n11925), .I2(n11924), .I3(n11923), .O(n11929) );
  OR_GATE U12387 ( .I1(n11927), .I2(n11926), .O(n11928) );
  NAND3_GATE U12388 ( .I1(n11930), .I2(n11929), .I3(n11928), .O(n12303) );
  NAND_GATE U12389 ( .I1(n1410), .I2(A[22]), .O(n12301) );
  INV_GATE U12390 ( .I1(n12301), .O(n12299) );
  NAND_GATE U12391 ( .I1(n438), .I2(n12299), .O(n12297) );
  NAND_GATE U12392 ( .I1(n1409), .I2(A[21]), .O(n12307) );
  INV_GATE U12393 ( .I1(n12307), .O(n12206) );
  OR_GATE U12394 ( .I1(n11931), .I2(n11936), .O(n11934) );
  OR_GATE U12395 ( .I1(n11935), .I2(n11932), .O(n11933) );
  NAND_GATE U12396 ( .I1(n996), .I2(n11935), .O(n11939) );
  NAND3_GATE U12397 ( .I1(n11939), .I2(n11938), .I3(n11937), .O(n11940) );
  NAND_GATE U12398 ( .I1(n1409), .I2(A[20]), .O(n12586) );
  INV_GATE U12399 ( .I1(n12586), .O(n12581) );
  NAND_GATE U12400 ( .I1(n12585), .I2(n12581), .O(n12578) );
  NAND_GATE U12401 ( .I1(n1409), .I2(A[19]), .O(n12323) );
  INV_GATE U12402 ( .I1(n12323), .O(n12192) );
  OR_GATE U12403 ( .I1(n11941), .I2(n11946), .O(n11944) );
  OR_GATE U12404 ( .I1(n11945), .I2(n11942), .O(n11943) );
  AND_GATE U12405 ( .I1(n11944), .I2(n11943), .O(n11951) );
  NAND_GATE U12406 ( .I1(n999), .I2(n11945), .O(n11949) );
  NAND3_GATE U12407 ( .I1(n11949), .I2(n11948), .I3(n11947), .O(n11950) );
  NAND_GATE U12408 ( .I1(n11951), .I2(n11950), .O(n12330) );
  NAND_GATE U12409 ( .I1(n1409), .I2(A[18]), .O(n12333) );
  NAND_GATE U12410 ( .I1(n85), .I2(n461), .O(n12327) );
  OR_GATE U12411 ( .I1(n771), .I2(n111), .O(n11962) );
  NAND_GATE U12412 ( .I1(n771), .I2(n11953), .O(n11958) );
  NAND_GATE U12413 ( .I1(n11954), .I2(n11958), .O(n11961) );
  NAND_GATE U12414 ( .I1(n11956), .I2(n11955), .O(n11957) );
  NAND_GATE U12415 ( .I1(n11958), .I2(n11957), .O(n11959) );
  OR_GATE U12416 ( .I1(n11963), .I2(n11967), .O(n11966) );
  OR_GATE U12417 ( .I1(n11964), .I2(n11968), .O(n11965) );
  AND_GATE U12418 ( .I1(n11966), .I2(n11965), .O(n11973) );
  NAND_GATE U12419 ( .I1(n11967), .I2(n1036), .O(n11971) );
  NAND3_GATE U12420 ( .I1(n11971), .I2(n11970), .I3(n11969), .O(n11972) );
  NAND_GATE U12421 ( .I1(n11973), .I2(n11972), .O(n12340) );
  INV_GATE U12422 ( .I1(n12340), .O(n12343) );
  OR_GATE U12423 ( .I1(n11974), .I2(n11976), .O(n11987) );
  NAND_GATE U12424 ( .I1(n11976), .I2(n11975), .O(n11981) );
  NAND_GATE U12425 ( .I1(n11977), .I2(n11981), .O(n11985) );
  NAND_GATE U12426 ( .I1(n11979), .I2(n11978), .O(n11980) );
  NAND_GATE U12427 ( .I1(n11981), .I2(n11980), .O(n11982) );
  NAND_GATE U12428 ( .I1(n11983), .I2(n11982), .O(n11984) );
  NAND_GATE U12429 ( .I1(n11985), .I2(n11984), .O(n11986) );
  NAND_GATE U12430 ( .I1(n11987), .I2(n11986), .O(n12354) );
  OR_GATE U12431 ( .I1(n11988), .I2(n11992), .O(n11991) );
  OR_GATE U12432 ( .I1(n11989), .I2(n11993), .O(n11990) );
  NAND_GATE U12433 ( .I1(n11992), .I2(n1054), .O(n11996) );
  NAND3_GATE U12434 ( .I1(n11996), .I2(n11995), .I3(n11994), .O(n11997) );
  INV_GATE U12435 ( .I1(n12362), .O(n12365) );
  OR_GATE U12436 ( .I1(n11998), .I2(n12000), .O(n12011) );
  NAND_GATE U12437 ( .I1(n12000), .I2(n11999), .O(n12005) );
  NAND_GATE U12438 ( .I1(n12001), .I2(n12005), .O(n12009) );
  NAND_GATE U12439 ( .I1(n12003), .I2(n12002), .O(n12004) );
  NAND_GATE U12440 ( .I1(n12005), .I2(n12004), .O(n12006) );
  NAND_GATE U12441 ( .I1(n12007), .I2(n12006), .O(n12008) );
  NAND_GATE U12442 ( .I1(n12009), .I2(n12008), .O(n12010) );
  NAND_GATE U12443 ( .I1(n12011), .I2(n12010), .O(n12378) );
  OR_GATE U12444 ( .I1(n12012), .I2(n12016), .O(n12015) );
  OR_GATE U12445 ( .I1(n12013), .I2(n12017), .O(n12014) );
  AND_GATE U12446 ( .I1(n12015), .I2(n12014), .O(n12022) );
  NAND_GATE U12447 ( .I1(n12016), .I2(n1066), .O(n12020) );
  NAND3_GATE U12448 ( .I1(n12020), .I2(n12019), .I3(n12018), .O(n12021) );
  NAND_GATE U12449 ( .I1(n12022), .I2(n12021), .O(n12387) );
  INV_GATE U12450 ( .I1(n12387), .O(n12390) );
  OR_GATE U12451 ( .I1(n12023), .I2(n12025), .O(n12036) );
  NAND_GATE U12452 ( .I1(n12025), .I2(n12024), .O(n12030) );
  NAND_GATE U12453 ( .I1(n12026), .I2(n12030), .O(n12034) );
  NAND_GATE U12454 ( .I1(n12028), .I2(n12027), .O(n12029) );
  NAND_GATE U12455 ( .I1(n12030), .I2(n12029), .O(n12031) );
  NAND_GATE U12456 ( .I1(n12032), .I2(n12031), .O(n12033) );
  NAND_GATE U12457 ( .I1(n12034), .I2(n12033), .O(n12035) );
  NAND_GATE U12458 ( .I1(n12036), .I2(n12035), .O(n12403) );
  OR_GATE U12459 ( .I1(n12037), .I2(n12041), .O(n12040) );
  OR_GATE U12460 ( .I1(n12038), .I2(n12042), .O(n12039) );
  AND_GATE U12461 ( .I1(n12040), .I2(n12039), .O(n12047) );
  NAND_GATE U12462 ( .I1(n12041), .I2(n1075), .O(n12045) );
  NAND3_GATE U12463 ( .I1(n12045), .I2(n12044), .I3(n12043), .O(n12046) );
  NAND_GATE U12464 ( .I1(n12047), .I2(n12046), .O(n12412) );
  INV_GATE U12465 ( .I1(n12412), .O(n12415) );
  OR_GATE U12466 ( .I1(n12048), .I2(n12050), .O(n12061) );
  NAND_GATE U12467 ( .I1(n12050), .I2(n12049), .O(n12055) );
  NAND_GATE U12468 ( .I1(n12051), .I2(n12055), .O(n12059) );
  NAND_GATE U12469 ( .I1(n12053), .I2(n12052), .O(n12054) );
  NAND_GATE U12470 ( .I1(n12055), .I2(n12054), .O(n12056) );
  NAND_GATE U12471 ( .I1(n12057), .I2(n12056), .O(n12058) );
  NAND_GATE U12472 ( .I1(n12059), .I2(n12058), .O(n12060) );
  NAND_GATE U12473 ( .I1(n12061), .I2(n12060), .O(n12428) );
  OR_GATE U12474 ( .I1(n12062), .I2(n12066), .O(n12065) );
  OR_GATE U12475 ( .I1(n12063), .I2(n12067), .O(n12064) );
  AND_GATE U12476 ( .I1(n12065), .I2(n12064), .O(n12072) );
  NAND_GATE U12477 ( .I1(n12066), .I2(n1083), .O(n12070) );
  NAND3_GATE U12478 ( .I1(n12070), .I2(n12069), .I3(n12068), .O(n12071) );
  NAND_GATE U12479 ( .I1(n12072), .I2(n12071), .O(n12437) );
  INV_GATE U12480 ( .I1(n12437), .O(n12440) );
  OR_GATE U12481 ( .I1(n12073), .I2(n12075), .O(n12086) );
  NAND_GATE U12482 ( .I1(n12075), .I2(n12074), .O(n12080) );
  NAND_GATE U12483 ( .I1(n12076), .I2(n12080), .O(n12084) );
  NAND_GATE U12484 ( .I1(n12078), .I2(n12077), .O(n12079) );
  NAND_GATE U12485 ( .I1(n12080), .I2(n12079), .O(n12081) );
  NAND_GATE U12486 ( .I1(n12082), .I2(n12081), .O(n12083) );
  NAND_GATE U12487 ( .I1(n12084), .I2(n12083), .O(n12085) );
  NAND_GATE U12488 ( .I1(n12086), .I2(n12085), .O(n12453) );
  OR_GATE U12489 ( .I1(n12087), .I2(n12091), .O(n12090) );
  OR_GATE U12490 ( .I1(n12088), .I2(n12092), .O(n12089) );
  AND_GATE U12491 ( .I1(n12090), .I2(n12089), .O(n12097) );
  NAND_GATE U12492 ( .I1(n12091), .I2(n1187), .O(n12095) );
  NAND3_GATE U12493 ( .I1(n12095), .I2(n12094), .I3(n12093), .O(n12096) );
  NAND_GATE U12494 ( .I1(n12097), .I2(n12096), .O(n12462) );
  INV_GATE U12495 ( .I1(n12462), .O(n12465) );
  OR_GATE U12496 ( .I1(n12098), .I2(n12100), .O(n12111) );
  NAND_GATE U12497 ( .I1(n12100), .I2(n12099), .O(n12105) );
  NAND_GATE U12498 ( .I1(n12101), .I2(n12105), .O(n12109) );
  NAND_GATE U12499 ( .I1(n12103), .I2(n12102), .O(n12104) );
  NAND_GATE U12500 ( .I1(n12105), .I2(n12104), .O(n12106) );
  NAND_GATE U12501 ( .I1(n12107), .I2(n12106), .O(n12108) );
  NAND_GATE U12502 ( .I1(n12109), .I2(n12108), .O(n12110) );
  NAND_GATE U12503 ( .I1(n12111), .I2(n12110), .O(n12478) );
  OR_GATE U12504 ( .I1(n12112), .I2(n12116), .O(n12115) );
  OR_GATE U12505 ( .I1(n12113), .I2(n12117), .O(n12114) );
  AND_GATE U12506 ( .I1(n12115), .I2(n12114), .O(n12122) );
  NAND_GATE U12507 ( .I1(n12116), .I2(n1246), .O(n12120) );
  NAND3_GATE U12508 ( .I1(n12120), .I2(n12119), .I3(n12118), .O(n12121) );
  NAND_GATE U12509 ( .I1(n12122), .I2(n12121), .O(n12487) );
  INV_GATE U12510 ( .I1(n12487), .O(n12490) );
  INV_GATE U12511 ( .I1(n12123), .O(n12124) );
  NAND_GATE U12512 ( .I1(n12128), .I2(n12124), .O(n12136) );
  NAND_GATE U12513 ( .I1(n12126), .I2(n12130), .O(n12134) );
  NAND_GATE U12514 ( .I1(n12128), .I2(n12127), .O(n12129) );
  NAND_GATE U12515 ( .I1(n12130), .I2(n12129), .O(n12131) );
  NAND_GATE U12516 ( .I1(n12132), .I2(n12131), .O(n12133) );
  NAND_GATE U12517 ( .I1(n12134), .I2(n12133), .O(n12135) );
  NAND_GATE U12518 ( .I1(n12136), .I2(n12135), .O(n12503) );
  NAND_GATE U12519 ( .I1(n1412), .I2(A[0]), .O(n12137) );
  NAND_GATE U12520 ( .I1(n14241), .I2(n12137), .O(n12138) );
  NAND_GATE U12521 ( .I1(n1413), .I2(n12138), .O(n12142) );
  NAND_GATE U12522 ( .I1(n1414), .I2(A[1]), .O(n12139) );
  NAND_GATE U12523 ( .I1(n724), .I2(n12139), .O(n12140) );
  NAND_GATE U12524 ( .I1(B[6]), .I2(n12140), .O(n12141) );
  NAND_GATE U12525 ( .I1(n12142), .I2(n12141), .O(n12515) );
  NAND_GATE U12526 ( .I1(n1409), .I2(A[2]), .O(n12519) );
  NAND3_GATE U12527 ( .I1(n1409), .I2(B[6]), .I3(n1254), .O(n12512) );
  NAND_GATE U12528 ( .I1(n12519), .I2(n12512), .O(n12143) );
  NAND_GATE U12529 ( .I1(n12515), .I2(n12143), .O(n12144) );
  INV_GATE U12530 ( .I1(n12519), .O(n12513) );
  INV_GATE U12531 ( .I1(n12512), .O(n12514) );
  NAND_GATE U12532 ( .I1(n12513), .I2(n12514), .O(n12510) );
  NAND_GATE U12533 ( .I1(n12144), .I2(n12510), .O(n12504) );
  NAND_GATE U12534 ( .I1(n12503), .I2(n12504), .O(n12146) );
  NAND_GATE U12535 ( .I1(n1409), .I2(A[3]), .O(n12505) );
  INV_GATE U12536 ( .I1(n12505), .O(n12145) );
  NAND_GATE U12537 ( .I1(n12503), .I2(n12145), .O(n12500) );
  NAND_GATE U12538 ( .I1(n12504), .I2(n12145), .O(n12499) );
  NAND3_GATE U12539 ( .I1(n12146), .I2(n12500), .I3(n12499), .O(n12489) );
  INV_GATE U12540 ( .I1(n12489), .O(n12486) );
  NAND_GATE U12541 ( .I1(n1409), .I2(A[4]), .O(n12494) );
  NAND_GATE U12542 ( .I1(n12486), .I2(n12494), .O(n12147) );
  NAND_GATE U12543 ( .I1(n12490), .I2(n12147), .O(n12148) );
  INV_GATE U12544 ( .I1(n12494), .O(n12488) );
  NAND_GATE U12545 ( .I1(n12489), .I2(n12488), .O(n12485) );
  NAND_GATE U12546 ( .I1(n12148), .I2(n12485), .O(n12479) );
  NAND_GATE U12547 ( .I1(n12478), .I2(n12479), .O(n12150) );
  NAND_GATE U12548 ( .I1(n1409), .I2(A[5]), .O(n12480) );
  INV_GATE U12549 ( .I1(n12480), .O(n12149) );
  NAND_GATE U12550 ( .I1(n12478), .I2(n12149), .O(n12475) );
  NAND_GATE U12551 ( .I1(n12479), .I2(n12149), .O(n12474) );
  NAND3_GATE U12552 ( .I1(n12150), .I2(n12475), .I3(n12474), .O(n12464) );
  INV_GATE U12553 ( .I1(n12464), .O(n12461) );
  NAND_GATE U12554 ( .I1(n1410), .I2(A[6]), .O(n12469) );
  NAND_GATE U12555 ( .I1(n12461), .I2(n12469), .O(n12151) );
  NAND_GATE U12556 ( .I1(n12465), .I2(n12151), .O(n12152) );
  INV_GATE U12557 ( .I1(n12469), .O(n12463) );
  NAND_GATE U12558 ( .I1(n12464), .I2(n12463), .O(n12460) );
  NAND_GATE U12559 ( .I1(n12152), .I2(n12460), .O(n12454) );
  NAND_GATE U12560 ( .I1(n12453), .I2(n12454), .O(n12154) );
  NAND_GATE U12561 ( .I1(n1410), .I2(A[7]), .O(n12455) );
  INV_GATE U12562 ( .I1(n12455), .O(n12153) );
  NAND_GATE U12563 ( .I1(n12453), .I2(n12153), .O(n12450) );
  NAND_GATE U12564 ( .I1(n12454), .I2(n12153), .O(n12449) );
  NAND3_GATE U12565 ( .I1(n12154), .I2(n12450), .I3(n12449), .O(n12439) );
  INV_GATE U12566 ( .I1(n12439), .O(n12436) );
  NAND_GATE U12567 ( .I1(n1410), .I2(A[8]), .O(n12444) );
  NAND_GATE U12568 ( .I1(n12436), .I2(n12444), .O(n12155) );
  NAND_GATE U12569 ( .I1(n12440), .I2(n12155), .O(n12156) );
  INV_GATE U12570 ( .I1(n12444), .O(n12438) );
  NAND_GATE U12571 ( .I1(n12439), .I2(n12438), .O(n12435) );
  NAND_GATE U12572 ( .I1(n12156), .I2(n12435), .O(n12429) );
  NAND_GATE U12573 ( .I1(n12428), .I2(n12429), .O(n12158) );
  NAND_GATE U12574 ( .I1(n1410), .I2(A[9]), .O(n12430) );
  INV_GATE U12575 ( .I1(n12430), .O(n12157) );
  NAND_GATE U12576 ( .I1(n12428), .I2(n12157), .O(n12425) );
  NAND_GATE U12577 ( .I1(n12429), .I2(n12157), .O(n12424) );
  NAND3_GATE U12578 ( .I1(n12158), .I2(n12425), .I3(n12424), .O(n12414) );
  INV_GATE U12579 ( .I1(n12414), .O(n12411) );
  NAND_GATE U12580 ( .I1(n1410), .I2(A[10]), .O(n12419) );
  NAND_GATE U12581 ( .I1(n12411), .I2(n12419), .O(n12159) );
  NAND_GATE U12582 ( .I1(n12415), .I2(n12159), .O(n12160) );
  INV_GATE U12583 ( .I1(n12419), .O(n12413) );
  NAND_GATE U12584 ( .I1(n12414), .I2(n12413), .O(n12410) );
  NAND_GATE U12585 ( .I1(n12160), .I2(n12410), .O(n12404) );
  NAND_GATE U12586 ( .I1(n12403), .I2(n12404), .O(n12162) );
  NAND_GATE U12587 ( .I1(n1410), .I2(A[11]), .O(n12405) );
  INV_GATE U12588 ( .I1(n12405), .O(n12161) );
  NAND_GATE U12589 ( .I1(n12403), .I2(n12161), .O(n12400) );
  NAND_GATE U12590 ( .I1(n12404), .I2(n12161), .O(n12399) );
  NAND3_GATE U12591 ( .I1(n12162), .I2(n12400), .I3(n12399), .O(n12389) );
  INV_GATE U12592 ( .I1(n12389), .O(n12386) );
  NAND_GATE U12593 ( .I1(n1410), .I2(A[12]), .O(n12394) );
  NAND_GATE U12594 ( .I1(n12386), .I2(n12394), .O(n12163) );
  NAND_GATE U12595 ( .I1(n12390), .I2(n12163), .O(n12164) );
  INV_GATE U12596 ( .I1(n12394), .O(n12388) );
  NAND_GATE U12597 ( .I1(n12389), .I2(n12388), .O(n12385) );
  NAND_GATE U12598 ( .I1(n12164), .I2(n12385), .O(n12379) );
  NAND_GATE U12599 ( .I1(n12378), .I2(n12379), .O(n12166) );
  NAND_GATE U12600 ( .I1(n1410), .I2(A[13]), .O(n12380) );
  INV_GATE U12601 ( .I1(n12380), .O(n12165) );
  NAND_GATE U12602 ( .I1(n12378), .I2(n12165), .O(n12375) );
  NAND_GATE U12603 ( .I1(n12379), .I2(n12165), .O(n12374) );
  NAND3_GATE U12604 ( .I1(n12166), .I2(n12375), .I3(n12374), .O(n12364) );
  INV_GATE U12605 ( .I1(n12364), .O(n12361) );
  NAND_GATE U12606 ( .I1(n1410), .I2(A[14]), .O(n12369) );
  NAND_GATE U12607 ( .I1(n12361), .I2(n12369), .O(n12167) );
  NAND_GATE U12608 ( .I1(n12365), .I2(n12167), .O(n12168) );
  INV_GATE U12609 ( .I1(n12369), .O(n12363) );
  NAND_GATE U12610 ( .I1(n12364), .I2(n12363), .O(n12360) );
  NAND_GATE U12611 ( .I1(n12168), .I2(n12360), .O(n12355) );
  NAND_GATE U12612 ( .I1(n12354), .I2(n12355), .O(n12170) );
  NAND_GATE U12613 ( .I1(n1410), .I2(A[15]), .O(n12356) );
  INV_GATE U12614 ( .I1(n12356), .O(n12169) );
  NAND_GATE U12615 ( .I1(n12354), .I2(n12169), .O(n12351) );
  NAND_GATE U12616 ( .I1(n12355), .I2(n12169), .O(n12350) );
  NAND3_GATE U12617 ( .I1(n12170), .I2(n12351), .I3(n12350), .O(n12342) );
  INV_GATE U12618 ( .I1(n12342), .O(n12339) );
  NAND_GATE U12619 ( .I1(n1410), .I2(A[16]), .O(n12347) );
  NAND_GATE U12620 ( .I1(n12339), .I2(n12347), .O(n12171) );
  NAND_GATE U12621 ( .I1(n12343), .I2(n12171), .O(n12172) );
  INV_GATE U12622 ( .I1(n12347), .O(n12341) );
  NAND_GATE U12623 ( .I1(n12342), .I2(n12341), .O(n12338) );
  NAND_GATE U12624 ( .I1(n12172), .I2(n12338), .O(n12567) );
  NAND_GATE U12625 ( .I1(n12566), .I2(n12567), .O(n12174) );
  NAND_GATE U12626 ( .I1(n1410), .I2(A[17]), .O(n12568) );
  INV_GATE U12627 ( .I1(n12568), .O(n12173) );
  NAND_GATE U12628 ( .I1(n12567), .I2(n12173), .O(n12563) );
  NAND_GATE U12629 ( .I1(n12566), .I2(n12173), .O(n12562) );
  NAND3_GATE U12630 ( .I1(n12174), .I2(n12563), .I3(n12562), .O(n12331) );
  NAND_GATE U12631 ( .I1(n12330), .I2(n12333), .O(n12175) );
  NAND_GATE U12632 ( .I1(n12331), .I2(n12175), .O(n12176) );
  NAND_GATE U12633 ( .I1(n12327), .I2(n12176), .O(n12322) );
  NAND_GATE U12634 ( .I1(n12192), .I2(n12322), .O(n12318) );
  INV_GATE U12635 ( .I1(n12177), .O(n12178) );
  NAND_GATE U12636 ( .I1(n12178), .I2(n12183), .O(n12191) );
  INV_GATE U12637 ( .I1(n12183), .O(n12181) );
  NAND_GATE U12638 ( .I1(n12182), .I2(n12181), .O(n12179) );
  NAND_GATE U12639 ( .I1(n12180), .I2(n12179), .O(n12189) );
  NAND_GATE U12640 ( .I1(n12179), .I2(n12185), .O(n12186) );
  NAND_GATE U12641 ( .I1(n12187), .I2(n12186), .O(n12188) );
  NAND_GATE U12642 ( .I1(n12189), .I2(n12188), .O(n12190) );
  NAND_GATE U12643 ( .I1(n12191), .I2(n12190), .O(n12321) );
  NAND_GATE U12644 ( .I1(n12322), .I2(n12321), .O(n12193) );
  NAND_GATE U12645 ( .I1(n12192), .I2(n12321), .O(n12317) );
  NAND3_GATE U12646 ( .I1(n12318), .I2(n12193), .I3(n12317), .O(n12584) );
  NAND_GATE U12647 ( .I1(n12583), .I2(n12586), .O(n12194) );
  NAND_GATE U12648 ( .I1(n12584), .I2(n12194), .O(n12195) );
  NAND_GATE U12649 ( .I1(n12578), .I2(n12195), .O(n12310) );
  NAND_GATE U12650 ( .I1(n12206), .I2(n12310), .O(n12312) );
  INV_GATE U12651 ( .I1(n12196), .O(n12197) );
  NAND_GATE U12652 ( .I1(n12197), .I2(n12199), .O(n12205) );
  NAND_GATE U12653 ( .I1(n434), .I2(n12200), .O(n12203) );
  NAND_GATE U12654 ( .I1(n12203), .I2(n12202), .O(n12204) );
  NAND_GATE U12655 ( .I1(n12205), .I2(n12204), .O(n12313) );
  NAND_GATE U12656 ( .I1(n12310), .I2(n12313), .O(n12207) );
  NAND_GATE U12657 ( .I1(n12206), .I2(n12313), .O(n12311) );
  NAND3_GATE U12658 ( .I1(n12312), .I2(n12207), .I3(n12311), .O(n12300) );
  NAND_GATE U12659 ( .I1(n12303), .I2(n12301), .O(n12208) );
  NAND_GATE U12660 ( .I1(n12300), .I2(n12208), .O(n12209) );
  NAND_GATE U12661 ( .I1(n12297), .I2(n12209), .O(n12292) );
  NAND_GATE U12662 ( .I1(n12293), .I2(n12292), .O(n12211) );
  NAND_GATE U12663 ( .I1(n12210), .I2(n12292), .O(n12289) );
  NAND3_GATE U12664 ( .I1(n12288), .I2(n12211), .I3(n12289), .O(n12285) );
  NAND3_GATE U12665 ( .I1(n12213), .I2(n12212), .I3(n12285), .O(n12214) );
  NAND_GATE U12666 ( .I1(n12284), .I2(n12214), .O(n12604) );
  NAND3_GATE U12667 ( .I1(n12604), .I2(n12613), .I3(n12611), .O(n12215) );
  NAND_GATE U12668 ( .I1(n12612), .I2(n12604), .O(n12609) );
  NAND3_GATE U12669 ( .I1(n12218), .I2(n12217), .I3(n494), .O(n12219) );
  NAND_GATE U12670 ( .I1(n12220), .I2(n12219), .O(n12276) );
  NAND_GATE U12671 ( .I1(n12221), .I2(n12276), .O(n12268) );
  NAND3_GATE U12672 ( .I1(n12276), .I2(n12266), .I3(n12222), .O(n12223) );
  NAND3_GATE U12673 ( .I1(n12271), .I2(n12268), .I3(n12223), .O(n12263) );
  NAND3_GATE U12674 ( .I1(n12225), .I2(n12224), .I3(n12263), .O(n12226) );
  NAND_GATE U12675 ( .I1(n12262), .I2(n12226), .O(n12634) );
  NAND4_GATE U12676 ( .I1(n12247), .I2(n12246), .I3(n12248), .I4(n12634), .O(
        n12228) );
  NAND_GATE U12677 ( .I1(n12655), .I2(n12634), .O(n12227) );
  NAND3_GATE U12678 ( .I1(n12249), .I2(n12228), .I3(n12227), .O(n13080) );
  NAND_GATE U12679 ( .I1(n13082), .I2(n13086), .O(n12229) );
  NAND_GATE U12680 ( .I1(n13080), .I2(n12229), .O(n12231) );
  NAND_GATE U12681 ( .I1(n1411), .I2(A[31]), .O(n12230) );
  NAND3_GATE U12682 ( .I1(n12232), .I2(n12231), .I3(n12230), .O(n12641) );
  NAND_GATE U12683 ( .I1(n12640), .I2(n12641), .O(n12240) );
  INV_GATE U12684 ( .I1(n12240), .O(n14821) );
  NAND_GATE U12685 ( .I1(n12234), .I2(n12233), .O(n12236) );
  OR_GATE U12686 ( .I1(n12236), .I2(n12235), .O(n12237) );
  NAND_GATE U12687 ( .I1(n12238), .I2(n12237), .O(n12239) );
  NAND_GATE U12688 ( .I1(n14821), .I2(n12239), .O(n12242) );
  NAND_GATE U12689 ( .I1(n12240), .I2(n14820), .O(n12241) );
  NAND_GATE U12690 ( .I1(n12242), .I2(n12241), .O(\A1[35] ) );
  INV_GATE U12691 ( .I1(n13080), .O(n13081) );
  NAND3_GATE U12692 ( .I1(n13086), .I2(n13081), .I3(n13082), .O(n12243) );
  NAND_GATE U12693 ( .I1(n12244), .I2(n13083), .O(n13078) );
  NAND3_GATE U12694 ( .I1(n13084), .I2(n12243), .I3(n13078), .O(n12245) );
  NAND3_GATE U12695 ( .I1(n12244), .I2(n13080), .I3(n716), .O(n13079) );
  NAND_GATE U12696 ( .I1(n12245), .I2(n13079), .O(n12639) );
  NAND_GATE U12697 ( .I1(n12247), .I2(n12246), .O(n12648) );
  NAND3_GATE U12698 ( .I1(n12250), .I2(n12634), .I3(n873), .O(n12656) );
  NAND3_GATE U12699 ( .I1(n12250), .I2(n12652), .I3(n12633), .O(n12658) );
  NAND_GATE U12700 ( .I1(B[4]), .I2(A[30]), .O(n12667) );
  INV_GATE U12701 ( .I1(n12667), .O(n12632) );
  INV_GATE U12702 ( .I1(n12249), .O(n12635) );
  NAND3_GATE U12703 ( .I1(n12634), .I2(n12632), .I3(n12635), .O(n12253) );
  NAND3_GATE U12704 ( .I1(n12632), .I2(n12652), .I3(n12633), .O(n12252) );
  NAND_GATE U12705 ( .I1(n12250), .I2(n12632), .O(n12251) );
  NAND3_GATE U12706 ( .I1(n12253), .I2(n12252), .I3(n12251), .O(n12254) );
  NAND_GATE U12707 ( .I1(n993), .I2(n12254), .O(n13077) );
  NAND_GATE U12708 ( .I1(B[4]), .I2(A[29]), .O(n12677) );
  INV_GATE U12709 ( .I1(n12677), .O(n12670) );
  INV_GATE U12710 ( .I1(n12263), .O(n12257) );
  NAND3_GATE U12711 ( .I1(n12258), .I2(n12257), .I3(n12256), .O(n12259) );
  NAND3_GATE U12712 ( .I1(n12261), .I2(n12260), .I3(n12259), .O(n12265) );
  NAND_GATE U12713 ( .I1(n912), .I2(n12263), .O(n12264) );
  NAND_GATE U12714 ( .I1(n12265), .I2(n12264), .O(n12673) );
  NAND_GATE U12715 ( .I1(n12670), .I2(n12673), .O(n12631) );
  NAND_GATE U12716 ( .I1(B[4]), .I2(A[28]), .O(n13103) );
  NAND_GATE U12717 ( .I1(n12273), .I2(n12272), .O(n12266) );
  NAND_GATE U12718 ( .I1(n12267), .I2(n12266), .O(n12270) );
  INV_GATE U12719 ( .I1(n12268), .O(n12269) );
  NAND3_GATE U12720 ( .I1(n12270), .I2(n12269), .I3(n12274), .O(n12282) );
  OR_GATE U12721 ( .I1(n12276), .I2(n12271), .O(n12281) );
  NAND3_GATE U12722 ( .I1(n12266), .I2(n658), .I3(n12222), .O(n12278) );
  NAND_GATE U12723 ( .I1(n12222), .I2(n12266), .O(n12275) );
  NAND_GATE U12724 ( .I1(n12276), .I2(n12275), .O(n12277) );
  NAND3_GATE U12725 ( .I1(n12279), .I2(n12278), .I3(n12277), .O(n12280) );
  NAND3_GATE U12726 ( .I1(n12282), .I2(n12281), .I3(n12280), .O(n13102) );
  NAND_GATE U12727 ( .I1(B[4]), .I2(A[27]), .O(n12687) );
  INV_GATE U12728 ( .I1(n12687), .O(n12695) );
  NAND_GATE U12729 ( .I1(n12283), .I2(n12287), .O(n12717) );
  NAND_GATE U12730 ( .I1(n1374), .I2(n12285), .O(n12286) );
  NAND_GATE U12731 ( .I1(n12287), .I2(n12286), .O(n12715) );
  NAND_GATE U12732 ( .I1(n12716), .I2(n12715), .O(n12707) );
  NAND_GATE U12733 ( .I1(B[4]), .I2(A[24]), .O(n13046) );
  OR_GATE U12734 ( .I1(n12292), .I2(n12288), .O(n12291) );
  OR_GATE U12735 ( .I1(n12289), .I2(n12293), .O(n12290) );
  NAND_GATE U12736 ( .I1(n12293), .I2(n269), .O(n12294) );
  NAND3_GATE U12737 ( .I1(n12296), .I2(n12295), .I3(n12294), .O(n12597) );
  NAND_GATE U12738 ( .I1(B[4]), .I2(A[23]), .O(n12727) );
  INV_GATE U12739 ( .I1(n12727), .O(n12595) );
  INV_GATE U12740 ( .I1(n12300), .O(n12302) );
  NAND_GATE U12741 ( .I1(n12299), .I2(n12298), .O(n12306) );
  NAND_GATE U12742 ( .I1(n438), .I2(n12300), .O(n12305) );
  NAND3_GATE U12743 ( .I1(n12303), .I2(n12302), .I3(n12301), .O(n12304) );
  NAND3_GATE U12744 ( .I1(n12306), .I2(n12305), .I3(n12304), .O(n12726) );
  NAND_GATE U12745 ( .I1(n12725), .I2(n12726), .O(n12732) );
  NAND_GATE U12746 ( .I1(n12595), .I2(n12732), .O(n12730) );
  NAND_GATE U12747 ( .I1(n134), .I2(n12313), .O(n12309) );
  NAND3_GATE U12748 ( .I1(n12309), .I2(n12308), .I3(n12307), .O(n12316) );
  OR_GATE U12749 ( .I1(n12311), .I2(n12310), .O(n12315) );
  OR_GATE U12750 ( .I1(n12313), .I2(n12312), .O(n12314) );
  NAND3_GATE U12751 ( .I1(n12316), .I2(n12315), .I3(n12314), .O(n13032) );
  INV_GATE U12752 ( .I1(n13032), .O(n13034) );
  NAND_GATE U12753 ( .I1(B[4]), .I2(A[22]), .O(n13035) );
  INV_GATE U12754 ( .I1(n13035), .O(n13031) );
  NAND_GATE U12755 ( .I1(n13034), .I2(n13031), .O(n13028) );
  NAND_GATE U12756 ( .I1(B[4]), .I2(A[21]), .O(n12743) );
  INV_GATE U12757 ( .I1(n12743), .O(n12591) );
  OR_GATE U12758 ( .I1(n12317), .I2(n12322), .O(n12320) );
  OR_GATE U12759 ( .I1(n12321), .I2(n12318), .O(n12319) );
  NAND_GATE U12760 ( .I1(n1028), .I2(n12321), .O(n12325) );
  NAND3_GATE U12761 ( .I1(n12325), .I2(n12324), .I3(n12323), .O(n12326) );
  NAND_GATE U12762 ( .I1(B[4]), .I2(A[20]), .O(n12752) );
  INV_GATE U12763 ( .I1(n12327), .O(n12328) );
  NAND_GATE U12764 ( .I1(n12328), .I2(n12331), .O(n12337) );
  INV_GATE U12765 ( .I1(n12331), .O(n12329) );
  NAND_GATE U12766 ( .I1(n12330), .I2(n12329), .O(n12332) );
  NAND_GATE U12767 ( .I1(n461), .I2(n12332), .O(n12335) );
  NAND_GATE U12768 ( .I1(n12335), .I2(n12334), .O(n12336) );
  NAND_GATE U12769 ( .I1(n12337), .I2(n12336), .O(n13016) );
  OR_GATE U12770 ( .I1(n12338), .I2(n12340), .O(n12349) );
  NAND_GATE U12771 ( .I1(n12340), .I2(n12339), .O(n12345) );
  NAND_GATE U12772 ( .I1(n12341), .I2(n12345), .O(n12348) );
  NAND_GATE U12773 ( .I1(n12343), .I2(n12342), .O(n12344) );
  NAND_GATE U12774 ( .I1(n12345), .I2(n12344), .O(n12346) );
  OR_GATE U12775 ( .I1(n12350), .I2(n12354), .O(n12353) );
  OR_GATE U12776 ( .I1(n12351), .I2(n12355), .O(n12352) );
  NAND_GATE U12777 ( .I1(n12354), .I2(n1042), .O(n12358) );
  NAND3_GATE U12778 ( .I1(n12358), .I2(n12357), .I3(n12356), .O(n12359) );
  INV_GATE U12779 ( .I1(n12773), .O(n12776) );
  OR_GATE U12780 ( .I1(n12360), .I2(n12362), .O(n12373) );
  NAND_GATE U12781 ( .I1(n12362), .I2(n12361), .O(n12367) );
  NAND_GATE U12782 ( .I1(n12363), .I2(n12367), .O(n12371) );
  NAND_GATE U12783 ( .I1(n12365), .I2(n12364), .O(n12366) );
  NAND_GATE U12784 ( .I1(n12367), .I2(n12366), .O(n12368) );
  NAND_GATE U12785 ( .I1(n12369), .I2(n12368), .O(n12370) );
  NAND_GATE U12786 ( .I1(n12371), .I2(n12370), .O(n12372) );
  NAND_GATE U12787 ( .I1(n12373), .I2(n12372), .O(n12789) );
  OR_GATE U12788 ( .I1(n12374), .I2(n12378), .O(n12377) );
  OR_GATE U12789 ( .I1(n12375), .I2(n12379), .O(n12376) );
  AND_GATE U12790 ( .I1(n12377), .I2(n12376), .O(n12384) );
  NAND_GATE U12791 ( .I1(n12378), .I2(n1061), .O(n12382) );
  NAND3_GATE U12792 ( .I1(n12382), .I2(n12381), .I3(n12380), .O(n12383) );
  NAND_GATE U12793 ( .I1(n12384), .I2(n12383), .O(n12798) );
  INV_GATE U12794 ( .I1(n12798), .O(n12801) );
  OR_GATE U12795 ( .I1(n12385), .I2(n12387), .O(n12398) );
  NAND_GATE U12796 ( .I1(n12387), .I2(n12386), .O(n12392) );
  NAND_GATE U12797 ( .I1(n12388), .I2(n12392), .O(n12396) );
  NAND_GATE U12798 ( .I1(n12390), .I2(n12389), .O(n12391) );
  NAND_GATE U12799 ( .I1(n12392), .I2(n12391), .O(n12393) );
  NAND_GATE U12800 ( .I1(n12394), .I2(n12393), .O(n12395) );
  NAND_GATE U12801 ( .I1(n12396), .I2(n12395), .O(n12397) );
  NAND_GATE U12802 ( .I1(n12398), .I2(n12397), .O(n12814) );
  OR_GATE U12803 ( .I1(n12399), .I2(n12403), .O(n12402) );
  OR_GATE U12804 ( .I1(n12400), .I2(n12404), .O(n12401) );
  AND_GATE U12805 ( .I1(n12402), .I2(n12401), .O(n12409) );
  NAND_GATE U12806 ( .I1(n12403), .I2(n1071), .O(n12407) );
  NAND3_GATE U12807 ( .I1(n12407), .I2(n12406), .I3(n12405), .O(n12408) );
  NAND_GATE U12808 ( .I1(n12409), .I2(n12408), .O(n12823) );
  INV_GATE U12809 ( .I1(n12823), .O(n12826) );
  OR_GATE U12810 ( .I1(n12410), .I2(n12412), .O(n12423) );
  NAND_GATE U12811 ( .I1(n12412), .I2(n12411), .O(n12417) );
  NAND_GATE U12812 ( .I1(n12413), .I2(n12417), .O(n12421) );
  NAND_GATE U12813 ( .I1(n12415), .I2(n12414), .O(n12416) );
  NAND_GATE U12814 ( .I1(n12417), .I2(n12416), .O(n12418) );
  NAND_GATE U12815 ( .I1(n12419), .I2(n12418), .O(n12420) );
  NAND_GATE U12816 ( .I1(n12421), .I2(n12420), .O(n12422) );
  NAND_GATE U12817 ( .I1(n12423), .I2(n12422), .O(n12839) );
  OR_GATE U12818 ( .I1(n12424), .I2(n12428), .O(n12427) );
  OR_GATE U12819 ( .I1(n12425), .I2(n12429), .O(n12426) );
  AND_GATE U12820 ( .I1(n12427), .I2(n12426), .O(n12434) );
  NAND_GATE U12821 ( .I1(n12428), .I2(n1079), .O(n12432) );
  NAND3_GATE U12822 ( .I1(n12432), .I2(n12431), .I3(n12430), .O(n12433) );
  NAND_GATE U12823 ( .I1(n12434), .I2(n12433), .O(n12848) );
  INV_GATE U12824 ( .I1(n12848), .O(n12851) );
  OR_GATE U12825 ( .I1(n12435), .I2(n12437), .O(n12448) );
  NAND_GATE U12826 ( .I1(n12437), .I2(n12436), .O(n12442) );
  NAND_GATE U12827 ( .I1(n12438), .I2(n12442), .O(n12446) );
  NAND_GATE U12828 ( .I1(n12440), .I2(n12439), .O(n12441) );
  NAND_GATE U12829 ( .I1(n12442), .I2(n12441), .O(n12443) );
  NAND_GATE U12830 ( .I1(n12444), .I2(n12443), .O(n12445) );
  NAND_GATE U12831 ( .I1(n12446), .I2(n12445), .O(n12447) );
  NAND_GATE U12832 ( .I1(n12448), .I2(n12447), .O(n12864) );
  OR_GATE U12833 ( .I1(n12449), .I2(n12453), .O(n12452) );
  OR_GATE U12834 ( .I1(n12450), .I2(n12454), .O(n12451) );
  AND_GATE U12835 ( .I1(n12452), .I2(n12451), .O(n12459) );
  NAND_GATE U12836 ( .I1(n12453), .I2(n1086), .O(n12457) );
  NAND3_GATE U12837 ( .I1(n12457), .I2(n12456), .I3(n12455), .O(n12458) );
  NAND_GATE U12838 ( .I1(n12459), .I2(n12458), .O(n12873) );
  INV_GATE U12839 ( .I1(n12873), .O(n12876) );
  OR_GATE U12840 ( .I1(n12460), .I2(n12462), .O(n12473) );
  NAND_GATE U12841 ( .I1(n12462), .I2(n12461), .O(n12467) );
  NAND_GATE U12842 ( .I1(n12463), .I2(n12467), .O(n12471) );
  NAND_GATE U12843 ( .I1(n12465), .I2(n12464), .O(n12466) );
  NAND_GATE U12844 ( .I1(n12467), .I2(n12466), .O(n12468) );
  NAND_GATE U12845 ( .I1(n12469), .I2(n12468), .O(n12470) );
  NAND_GATE U12846 ( .I1(n12471), .I2(n12470), .O(n12472) );
  NAND_GATE U12847 ( .I1(n12473), .I2(n12472), .O(n12889) );
  OR_GATE U12848 ( .I1(n12474), .I2(n12478), .O(n12477) );
  OR_GATE U12849 ( .I1(n12475), .I2(n12479), .O(n12476) );
  AND_GATE U12850 ( .I1(n12477), .I2(n12476), .O(n12484) );
  NAND_GATE U12851 ( .I1(n12478), .I2(n1189), .O(n12482) );
  NAND3_GATE U12852 ( .I1(n12482), .I2(n12481), .I3(n12480), .O(n12483) );
  NAND_GATE U12853 ( .I1(n12484), .I2(n12483), .O(n12898) );
  INV_GATE U12854 ( .I1(n12898), .O(n12901) );
  OR_GATE U12855 ( .I1(n12485), .I2(n12487), .O(n12498) );
  NAND_GATE U12856 ( .I1(n12487), .I2(n12486), .O(n12492) );
  NAND_GATE U12857 ( .I1(n12488), .I2(n12492), .O(n12496) );
  NAND_GATE U12858 ( .I1(n12490), .I2(n12489), .O(n12491) );
  NAND_GATE U12859 ( .I1(n12492), .I2(n12491), .O(n12493) );
  NAND_GATE U12860 ( .I1(n12494), .I2(n12493), .O(n12495) );
  NAND_GATE U12861 ( .I1(n12496), .I2(n12495), .O(n12497) );
  NAND_GATE U12862 ( .I1(n12498), .I2(n12497), .O(n12914) );
  OR_GATE U12863 ( .I1(n12499), .I2(n12503), .O(n12502) );
  OR_GATE U12864 ( .I1(n12500), .I2(n12504), .O(n12501) );
  AND_GATE U12865 ( .I1(n12502), .I2(n12501), .O(n12509) );
  NAND_GATE U12866 ( .I1(n12503), .I2(n1247), .O(n12507) );
  NAND3_GATE U12867 ( .I1(n12507), .I2(n12506), .I3(n12505), .O(n12508) );
  NAND_GATE U12868 ( .I1(n12509), .I2(n12508), .O(n12923) );
  INV_GATE U12869 ( .I1(n12923), .O(n12926) );
  INV_GATE U12870 ( .I1(n12510), .O(n12511) );
  NAND_GATE U12871 ( .I1(n12515), .I2(n12511), .O(n12523) );
  NAND_GATE U12872 ( .I1(n12513), .I2(n12517), .O(n12521) );
  NAND_GATE U12873 ( .I1(n12515), .I2(n12514), .O(n12516) );
  NAND_GATE U12874 ( .I1(n12517), .I2(n12516), .O(n12518) );
  NAND_GATE U12875 ( .I1(n12519), .I2(n12518), .O(n12520) );
  NAND_GATE U12876 ( .I1(n12521), .I2(n12520), .O(n12522) );
  NAND_GATE U12877 ( .I1(n12523), .I2(n12522), .O(n12939) );
  NAND_GATE U12878 ( .I1(n1411), .I2(A[0]), .O(n12524) );
  NAND_GATE U12879 ( .I1(n14241), .I2(n12524), .O(n12525) );
  NAND_GATE U12880 ( .I1(B[6]), .I2(n12525), .O(n12529) );
  NAND_GATE U12881 ( .I1(n1412), .I2(A[1]), .O(n12526) );
  NAND_GATE U12882 ( .I1(n724), .I2(n12526), .O(n12527) );
  NAND_GATE U12883 ( .I1(n1410), .I2(n12527), .O(n12528) );
  NAND_GATE U12884 ( .I1(n12529), .I2(n12528), .O(n12951) );
  NAND_GATE U12885 ( .I1(B[4]), .I2(A[2]), .O(n12955) );
  NAND3_GATE U12886 ( .I1(B[4]), .I2(n1410), .I3(n1254), .O(n12948) );
  NAND_GATE U12887 ( .I1(n12955), .I2(n12948), .O(n12530) );
  NAND_GATE U12888 ( .I1(n12951), .I2(n12530), .O(n12531) );
  INV_GATE U12889 ( .I1(n12955), .O(n12949) );
  INV_GATE U12890 ( .I1(n12948), .O(n12950) );
  NAND_GATE U12891 ( .I1(n12949), .I2(n12950), .O(n12946) );
  NAND_GATE U12892 ( .I1(n12531), .I2(n12946), .O(n12940) );
  NAND_GATE U12893 ( .I1(n12939), .I2(n12940), .O(n12533) );
  NAND_GATE U12894 ( .I1(B[4]), .I2(A[3]), .O(n12941) );
  INV_GATE U12895 ( .I1(n12941), .O(n12532) );
  NAND_GATE U12896 ( .I1(n12939), .I2(n12532), .O(n12936) );
  NAND_GATE U12897 ( .I1(n12940), .I2(n12532), .O(n12935) );
  NAND3_GATE U12898 ( .I1(n12533), .I2(n12936), .I3(n12935), .O(n12925) );
  INV_GATE U12899 ( .I1(n12925), .O(n12922) );
  NAND_GATE U12900 ( .I1(B[4]), .I2(A[4]), .O(n12930) );
  NAND_GATE U12901 ( .I1(n12922), .I2(n12930), .O(n12534) );
  NAND_GATE U12902 ( .I1(n12926), .I2(n12534), .O(n12535) );
  INV_GATE U12903 ( .I1(n12930), .O(n12924) );
  NAND_GATE U12904 ( .I1(n12925), .I2(n12924), .O(n12921) );
  NAND_GATE U12905 ( .I1(n12535), .I2(n12921), .O(n12915) );
  NAND_GATE U12906 ( .I1(n12914), .I2(n12915), .O(n12537) );
  NAND_GATE U12907 ( .I1(B[4]), .I2(A[5]), .O(n12916) );
  INV_GATE U12908 ( .I1(n12916), .O(n12536) );
  NAND_GATE U12909 ( .I1(n12914), .I2(n12536), .O(n12911) );
  NAND_GATE U12910 ( .I1(n12915), .I2(n12536), .O(n12910) );
  NAND3_GATE U12911 ( .I1(n12537), .I2(n12911), .I3(n12910), .O(n12900) );
  INV_GATE U12912 ( .I1(n12900), .O(n12897) );
  NAND_GATE U12913 ( .I1(B[4]), .I2(A[6]), .O(n12905) );
  NAND_GATE U12914 ( .I1(n12897), .I2(n12905), .O(n12538) );
  NAND_GATE U12915 ( .I1(n12901), .I2(n12538), .O(n12539) );
  INV_GATE U12916 ( .I1(n12905), .O(n12899) );
  NAND_GATE U12917 ( .I1(n12900), .I2(n12899), .O(n12896) );
  NAND_GATE U12918 ( .I1(n12539), .I2(n12896), .O(n12890) );
  NAND_GATE U12919 ( .I1(n12889), .I2(n12890), .O(n12541) );
  NAND_GATE U12920 ( .I1(B[4]), .I2(A[7]), .O(n12891) );
  INV_GATE U12921 ( .I1(n12891), .O(n12540) );
  NAND_GATE U12922 ( .I1(n12889), .I2(n12540), .O(n12886) );
  NAND_GATE U12923 ( .I1(n12890), .I2(n12540), .O(n12885) );
  NAND3_GATE U12924 ( .I1(n12541), .I2(n12886), .I3(n12885), .O(n12875) );
  INV_GATE U12925 ( .I1(n12875), .O(n12872) );
  NAND_GATE U12926 ( .I1(B[4]), .I2(A[8]), .O(n12880) );
  NAND_GATE U12927 ( .I1(n12872), .I2(n12880), .O(n12542) );
  NAND_GATE U12928 ( .I1(n12876), .I2(n12542), .O(n12543) );
  INV_GATE U12929 ( .I1(n12880), .O(n12874) );
  NAND_GATE U12930 ( .I1(n12875), .I2(n12874), .O(n12871) );
  NAND_GATE U12931 ( .I1(n12543), .I2(n12871), .O(n12865) );
  NAND_GATE U12932 ( .I1(n12864), .I2(n12865), .O(n12545) );
  NAND_GATE U12933 ( .I1(B[4]), .I2(A[9]), .O(n12866) );
  INV_GATE U12934 ( .I1(n12866), .O(n12544) );
  NAND_GATE U12935 ( .I1(n12864), .I2(n12544), .O(n12861) );
  NAND_GATE U12936 ( .I1(n12865), .I2(n12544), .O(n12860) );
  NAND3_GATE U12937 ( .I1(n12545), .I2(n12861), .I3(n12860), .O(n12850) );
  INV_GATE U12938 ( .I1(n12850), .O(n12847) );
  NAND_GATE U12939 ( .I1(B[4]), .I2(A[10]), .O(n12855) );
  NAND_GATE U12940 ( .I1(n12847), .I2(n12855), .O(n12546) );
  NAND_GATE U12941 ( .I1(n12851), .I2(n12546), .O(n12547) );
  INV_GATE U12942 ( .I1(n12855), .O(n12849) );
  NAND_GATE U12943 ( .I1(n12850), .I2(n12849), .O(n12846) );
  NAND_GATE U12944 ( .I1(n12547), .I2(n12846), .O(n12840) );
  NAND_GATE U12945 ( .I1(n12839), .I2(n12840), .O(n12549) );
  NAND_GATE U12946 ( .I1(B[4]), .I2(A[11]), .O(n12841) );
  INV_GATE U12947 ( .I1(n12841), .O(n12548) );
  NAND_GATE U12948 ( .I1(n12839), .I2(n12548), .O(n12836) );
  NAND_GATE U12949 ( .I1(n12840), .I2(n12548), .O(n12835) );
  NAND3_GATE U12950 ( .I1(n12549), .I2(n12836), .I3(n12835), .O(n12825) );
  INV_GATE U12951 ( .I1(n12825), .O(n12822) );
  NAND_GATE U12952 ( .I1(B[4]), .I2(A[12]), .O(n12830) );
  NAND_GATE U12953 ( .I1(n12822), .I2(n12830), .O(n12550) );
  NAND_GATE U12954 ( .I1(n12826), .I2(n12550), .O(n12551) );
  INV_GATE U12955 ( .I1(n12830), .O(n12824) );
  NAND_GATE U12956 ( .I1(n12825), .I2(n12824), .O(n12821) );
  NAND_GATE U12957 ( .I1(n12551), .I2(n12821), .O(n12815) );
  NAND_GATE U12958 ( .I1(n12814), .I2(n12815), .O(n12553) );
  NAND_GATE U12959 ( .I1(B[4]), .I2(A[13]), .O(n12816) );
  INV_GATE U12960 ( .I1(n12816), .O(n12552) );
  NAND_GATE U12961 ( .I1(n12814), .I2(n12552), .O(n12811) );
  NAND_GATE U12962 ( .I1(n12815), .I2(n12552), .O(n12810) );
  NAND3_GATE U12963 ( .I1(n12553), .I2(n12811), .I3(n12810), .O(n12800) );
  INV_GATE U12964 ( .I1(n12800), .O(n12797) );
  NAND_GATE U12965 ( .I1(B[4]), .I2(A[14]), .O(n12805) );
  NAND_GATE U12966 ( .I1(n12797), .I2(n12805), .O(n12554) );
  NAND_GATE U12967 ( .I1(n12801), .I2(n12554), .O(n12555) );
  INV_GATE U12968 ( .I1(n12805), .O(n12799) );
  NAND_GATE U12969 ( .I1(n12800), .I2(n12799), .O(n12796) );
  NAND_GATE U12970 ( .I1(n12555), .I2(n12796), .O(n12790) );
  NAND_GATE U12971 ( .I1(n12789), .I2(n12790), .O(n12557) );
  NAND_GATE U12972 ( .I1(B[4]), .I2(A[15]), .O(n12791) );
  INV_GATE U12973 ( .I1(n12791), .O(n12556) );
  NAND_GATE U12974 ( .I1(n12789), .I2(n12556), .O(n12786) );
  NAND_GATE U12975 ( .I1(n12790), .I2(n12556), .O(n12785) );
  NAND3_GATE U12976 ( .I1(n12557), .I2(n12786), .I3(n12785), .O(n12775) );
  INV_GATE U12977 ( .I1(n12775), .O(n12772) );
  NAND_GATE U12978 ( .I1(B[4]), .I2(A[16]), .O(n12780) );
  NAND_GATE U12979 ( .I1(n12772), .I2(n12780), .O(n12558) );
  NAND_GATE U12980 ( .I1(n12776), .I2(n12558), .O(n12559) );
  INV_GATE U12981 ( .I1(n12780), .O(n12774) );
  NAND_GATE U12982 ( .I1(n12775), .I2(n12774), .O(n12771) );
  NAND_GATE U12983 ( .I1(n12559), .I2(n12771), .O(n13003) );
  NAND_GATE U12984 ( .I1(n13002), .I2(n13003), .O(n12561) );
  NAND_GATE U12985 ( .I1(B[4]), .I2(A[17]), .O(n13004) );
  INV_GATE U12986 ( .I1(n13004), .O(n12560) );
  NAND_GATE U12987 ( .I1(n13003), .I2(n12560), .O(n12999) );
  NAND_GATE U12988 ( .I1(n13002), .I2(n12560), .O(n12998) );
  NAND3_GATE U12989 ( .I1(n12561), .I2(n12999), .I3(n12998), .O(n12762) );
  NAND_GATE U12990 ( .I1(B[4]), .I2(A[18]), .O(n12766) );
  OR_GATE U12991 ( .I1(n12562), .I2(n12567), .O(n12565) );
  OR_GATE U12992 ( .I1(n12563), .I2(n12566), .O(n12564) );
  NAND_GATE U12993 ( .I1(n12566), .I2(n1007), .O(n12570) );
  NAND3_GATE U12994 ( .I1(n12570), .I2(n12569), .I3(n12568), .O(n12571) );
  NAND_GATE U12995 ( .I1(n12766), .I2(n12759), .O(n12572) );
  NAND_GATE U12996 ( .I1(n12762), .I2(n12572), .O(n12573) );
  INV_GATE U12997 ( .I1(n12766), .O(n12760) );
  INV_GATE U12998 ( .I1(n12759), .O(n12761) );
  NAND_GATE U12999 ( .I1(n12760), .I2(n12761), .O(n12757) );
  NAND_GATE U13000 ( .I1(n12573), .I2(n12757), .O(n13017) );
  NAND_GATE U13001 ( .I1(n13016), .I2(n13017), .O(n12575) );
  NAND_GATE U13002 ( .I1(B[4]), .I2(A[19]), .O(n13018) );
  INV_GATE U13003 ( .I1(n13018), .O(n12574) );
  NAND_GATE U13004 ( .I1(n13017), .I2(n12574), .O(n13013) );
  NAND_GATE U13005 ( .I1(n13016), .I2(n12574), .O(n13012) );
  NAND3_GATE U13006 ( .I1(n12575), .I2(n13013), .I3(n13012), .O(n12750) );
  NAND_GATE U13007 ( .I1(n12749), .I2(n12752), .O(n12576) );
  NAND_GATE U13008 ( .I1(n12750), .I2(n12576), .O(n12577) );
  NAND_GATE U13009 ( .I1(n12747), .I2(n12577), .O(n12742) );
  INV_GATE U13010 ( .I1(n12578), .O(n12579) );
  NAND_GATE U13011 ( .I1(n12579), .I2(n12584), .O(n12590) );
  NAND_GATE U13012 ( .I1(n12583), .I2(n12582), .O(n12580) );
  NAND_GATE U13013 ( .I1(n12581), .I2(n12580), .O(n12588) );
  NAND_GATE U13014 ( .I1(n12588), .I2(n12587), .O(n12589) );
  NAND_GATE U13015 ( .I1(n12590), .I2(n12589), .O(n12741) );
  NAND_GATE U13016 ( .I1(n12742), .I2(n12741), .O(n12592) );
  NAND_GATE U13017 ( .I1(n12591), .I2(n12741), .O(n12737) );
  NAND3_GATE U13018 ( .I1(n12738), .I2(n12592), .I3(n12737), .O(n13033) );
  NAND_GATE U13019 ( .I1(n13032), .I2(n13035), .O(n12593) );
  NAND_GATE U13020 ( .I1(n13033), .I2(n12593), .O(n12594) );
  NAND_GATE U13021 ( .I1(n13028), .I2(n12594), .O(n12731) );
  NAND_GATE U13022 ( .I1(n12732), .I2(n12731), .O(n12596) );
  NAND_GATE U13023 ( .I1(n12595), .I2(n12731), .O(n12733) );
  NAND3_GATE U13024 ( .I1(n12730), .I2(n12596), .I3(n12733), .O(n13047) );
  NAND_GATE U13025 ( .I1(n13047), .I2(n12598), .O(n12599) );
  NAND_GATE U13026 ( .I1(n13044), .I2(n12706), .O(n12714) );
  NAND3_GATE U13027 ( .I1(n12708), .I2(n12707), .I3(n12714), .O(n12603) );
  NAND_GATE U13028 ( .I1(B[4]), .I2(A[25]), .O(n12712) );
  INV_GATE U13029 ( .I1(n12712), .O(n12600) );
  NAND3_GATE U13030 ( .I1(n12600), .I2(n12708), .I3(n12707), .O(n12713) );
  NAND_GATE U13031 ( .I1(n13044), .I2(n12599), .O(n12602) );
  NAND3_GATE U13032 ( .I1(n12602), .I2(n12601), .I3(n12600), .O(n12718) );
  NAND3_GATE U13033 ( .I1(n12603), .I2(n12713), .I3(n12718), .O(n12705) );
  NAND3_GATE U13034 ( .I1(n483), .I2(n12613), .I3(n12611), .O(n12605) );
  NAND4_GATE U13035 ( .I1(n12613), .I2(n483), .I3(n12612), .I4(n12611), .O(
        n12614) );
  NAND3_GATE U13036 ( .I1(n12705), .I2(n12616), .I3(n1262), .O(n12618) );
  NAND_GATE U13037 ( .I1(B[4]), .I2(A[26]), .O(n12704) );
  INV_GATE U13038 ( .I1(n12704), .O(n13483) );
  NAND_GATE U13039 ( .I1(n13483), .I2(n12705), .O(n12617) );
  NAND_GATE U13040 ( .I1(n1262), .I2(n12616), .O(n12702) );
  NAND3_GATE U13041 ( .I1(n12618), .I2(n12617), .I3(n12701), .O(n12684) );
  NAND_GATE U13042 ( .I1(n12695), .I2(n12684), .O(n12696) );
  NAND_GATE U13043 ( .I1(n12623), .I2(n494), .O(n12619) );
  NAND_GATE U13044 ( .I1(n12621), .I2(n12619), .O(n12688) );
  NAND_GATE U13045 ( .I1(n12620), .I2(n748), .O(n12621) );
  NAND_GATE U13046 ( .I1(n12622), .I2(n12621), .O(n12691) );
  INV_GATE U13047 ( .I1(n12691), .O(n12681) );
  NAND3_GATE U13048 ( .I1(n494), .I2(n12623), .I3(n12622), .O(n12693) );
  NAND_GATE U13049 ( .I1(n12681), .I2(n12693), .O(n12624) );
  NAND3_GATE U13050 ( .I1(n12690), .I2(n12624), .I3(n12684), .O(n12626) );
  NAND3_GATE U13051 ( .I1(n12624), .I2(n12695), .I3(n12690), .O(n12625) );
  NAND3_GATE U13052 ( .I1(n12696), .I2(n12626), .I3(n12625), .O(n13100) );
  NAND_GATE U13053 ( .I1(n13103), .I2(n13102), .O(n12627) );
  NAND_GATE U13054 ( .I1(n13100), .I2(n12627), .O(n12628) );
  NAND_GATE U13055 ( .I1(n13063), .I2(n12628), .O(n12674) );
  NAND_GATE U13056 ( .I1(n12674), .I2(n12673), .O(n12630) );
  NAND_GATE U13057 ( .I1(n12670), .I2(n12674), .O(n12629) );
  NAND3_GATE U13058 ( .I1(n12631), .I2(n12630), .I3(n12629), .O(n12664) );
  NAND_GATE U13059 ( .I1(n12632), .I2(n12664), .O(n13076) );
  NAND_GATE U13060 ( .I1(n1408), .I2(A[31]), .O(n13075) );
  NAND_GATE U13061 ( .I1(n12652), .I2(n12633), .O(n12636) );
  NAND_GATE U13062 ( .I1(n12635), .I2(n12634), .O(n12660) );
  NAND3_GATE U13063 ( .I1(n12655), .I2(n12636), .I3(n12660), .O(n12637) );
  NAND3_GATE U13064 ( .I1(n12637), .I2(n993), .I3(n12664), .O(n13074) );
  NAND4_GATE U13065 ( .I1(n13077), .I2(n13076), .I3(n13075), .I4(n13074), .O(
        n12638) );
  NAND_GATE U13066 ( .I1(n12639), .I2(n12638), .O(n13092) );
  INV_GATE U13067 ( .I1(n12641), .O(n12642) );
  NAND_GATE U13068 ( .I1(n12643), .I2(n12642), .O(n12644) );
  NAND_GATE U13069 ( .I1(n12240), .I2(n12644), .O(n12645) );
  NAND_GATE U13070 ( .I1(n280), .I2(n12645), .O(n12647) );
  NAND_GATE U13071 ( .I1(n12647), .I2(n12646), .O(\A1[34] ) );
  OR_GATE U13072 ( .I1(n13077), .I2(n12664), .O(n12662) );
  NAND_GATE U13073 ( .I1(n12652), .I2(n12648), .O(n12654) );
  NAND4_GATE U13074 ( .I1(n12652), .I2(n12651), .I3(n12650), .I4(n12649), .O(
        n12653) );
  NAND3_GATE U13075 ( .I1(n12655), .I2(n12654), .I3(n12653), .O(n12657) );
  NAND3_GATE U13076 ( .I1(n12658), .I2(n12657), .I3(n12656), .O(n12659) );
  NAND_GATE U13077 ( .I1(n12660), .I2(n12659), .O(n12663) );
  OR_GATE U13078 ( .I1(n12663), .I2(n13076), .O(n12661) );
  AND_GATE U13079 ( .I1(n12662), .I2(n12661), .O(n12669) );
  NAND_GATE U13080 ( .I1(n995), .I2(n12663), .O(n12666) );
  NAND3_GATE U13081 ( .I1(n12667), .I2(n12666), .I3(n12665), .O(n12668) );
  NAND_GATE U13082 ( .I1(n12669), .I2(n12668), .O(n13097) );
  NAND3_GATE U13083 ( .I1(n12670), .I2(n887), .I3(n12673), .O(n12671) );
  AND_GATE U13084 ( .I1(n12672), .I2(n12671), .O(n12679) );
  NAND_GATE U13085 ( .I1(n887), .I2(n12673), .O(n12676) );
  NAND3_GATE U13086 ( .I1(n12677), .I2(n12676), .I3(n12675), .O(n12678) );
  NAND_GATE U13087 ( .I1(n12679), .I2(n12678), .O(n13518) );
  INV_GATE U13088 ( .I1(n13518), .O(n13517) );
  NAND_GATE U13089 ( .I1(B[3]), .I2(A[30]), .O(n13516) );
  NAND_GATE U13090 ( .I1(n1407), .I2(A[31]), .O(n12680) );
  AND_GATE U13091 ( .I1(n13522), .I2(n12680), .O(n13073) );
  NAND_GATE U13092 ( .I1(B[3]), .I2(A[29]), .O(n13114) );
  INV_GATE U13093 ( .I1(n13114), .O(n13108) );
  NAND_GATE U13094 ( .I1(B[3]), .I2(A[28]), .O(n13502) );
  INV_GATE U13095 ( .I1(n13502), .O(n13506) );
  INV_GATE U13096 ( .I1(n12684), .O(n12694) );
  NAND_GATE U13097 ( .I1(n12682), .I2(n12690), .O(n12683) );
  NAND_GATE U13098 ( .I1(n12684), .I2(n12683), .O(n12685) );
  NAND3_GATE U13099 ( .I1(n12687), .I2(n12686), .I3(n12685), .O(n12700) );
  NAND_GATE U13100 ( .I1(n12691), .I2(n12690), .O(n12692) );
  NAND_GATE U13101 ( .I1(n12693), .I2(n12692), .O(n12697) );
  NAND3_GATE U13102 ( .I1(n12695), .I2(n12694), .I3(n12697), .O(n12699) );
  OR_GATE U13103 ( .I1(n12697), .I2(n12696), .O(n12698) );
  NAND3_GATE U13104 ( .I1(n12700), .I2(n12699), .I3(n12698), .O(n13504) );
  INV_GATE U13105 ( .I1(n13504), .O(n13503) );
  NAND_GATE U13106 ( .I1(n12702), .I2(n12703), .O(n13482) );
  NAND3_GATE U13107 ( .I1(n13482), .I2(n13488), .I3(n13483), .O(n13058) );
  NAND3_GATE U13108 ( .I1(n12704), .I2(n12703), .I3(n12702), .O(n13484) );
  NAND3_GATE U13109 ( .I1(n12705), .I2(n12704), .I3(n160), .O(n13485) );
  NAND_GATE U13110 ( .I1(B[3]), .I2(A[27]), .O(n13492) );
  INV_GATE U13111 ( .I1(n13492), .O(n13494) );
  NAND3_GATE U13112 ( .I1(n13058), .I2(n412), .I3(n13494), .O(n13060) );
  NAND4_GATE U13113 ( .I1(n13044), .I2(n12708), .I3(n12707), .I4(n12706), .O(
        n12711) );
  NAND_GATE U13114 ( .I1(n12708), .I2(n12707), .O(n12709) );
  NAND_GATE U13115 ( .I1(n12714), .I2(n12709), .O(n12710) );
  NAND3_GATE U13116 ( .I1(n12712), .I2(n12711), .I3(n12710), .O(n12724) );
  OR_GATE U13117 ( .I1(n12714), .I2(n12713), .O(n12723) );
  NAND_GATE U13118 ( .I1(n12717), .I2(n12707), .O(n12721) );
  INV_GATE U13119 ( .I1(n12718), .O(n12720) );
  NAND3_GATE U13120 ( .I1(n12721), .I2(n12720), .I3(n12719), .O(n12722) );
  NAND3_GATE U13121 ( .I1(n12724), .I2(n12723), .I3(n12722), .O(n13471) );
  INV_GATE U13122 ( .I1(n13471), .O(n13470) );
  NAND_GATE U13123 ( .I1(B[3]), .I2(A[26]), .O(n13473) );
  INV_GATE U13124 ( .I1(n13473), .O(n13468) );
  NAND_GATE U13125 ( .I1(n13470), .I2(n13468), .O(n13466) );
  NAND_GATE U13126 ( .I1(n12732), .I2(n487), .O(n12729) );
  NAND3_GATE U13127 ( .I1(n12726), .I2(n12725), .I3(n12731), .O(n12728) );
  NAND3_GATE U13128 ( .I1(n12729), .I2(n12728), .I3(n12727), .O(n12736) );
  OR_GATE U13129 ( .I1(n12731), .I2(n12730), .O(n12735) );
  OR_GATE U13130 ( .I1(n12733), .I2(n12732), .O(n12734) );
  NAND3_GATE U13131 ( .I1(n12736), .I2(n12735), .I3(n12734), .O(n13453) );
  NAND_GATE U13132 ( .I1(B[3]), .I2(A[24]), .O(n13456) );
  INV_GATE U13133 ( .I1(n13456), .O(n13452) );
  NAND_GATE U13134 ( .I1(n13455), .I2(n13452), .O(n13449) );
  NAND_GATE U13135 ( .I1(B[3]), .I2(A[23]), .O(n13138) );
  INV_GATE U13136 ( .I1(n13138), .O(n13040) );
  OR_GATE U13137 ( .I1(n12737), .I2(n12742), .O(n12740) );
  OR_GATE U13138 ( .I1(n12741), .I2(n12738), .O(n12739) );
  NAND_GATE U13139 ( .I1(n479), .I2(n12741), .O(n12745) );
  NAND3_GATE U13140 ( .I1(n12745), .I2(n12744), .I3(n12743), .O(n12746) );
  NAND_GATE U13141 ( .I1(B[3]), .I2(A[22]), .O(n13148) );
  INV_GATE U13142 ( .I1(n13148), .O(n13145) );
  NAND_GATE U13143 ( .I1(n451), .I2(n12750), .O(n12756) );
  INV_GATE U13144 ( .I1(n12750), .O(n12748) );
  NAND_GATE U13145 ( .I1(n12749), .I2(n12748), .O(n12751) );
  NAND_GATE U13146 ( .I1(n557), .I2(n12751), .O(n12754) );
  NAND_GATE U13147 ( .I1(n12754), .I2(n12753), .O(n12755) );
  NAND_GATE U13148 ( .I1(n12756), .I2(n12755), .O(n13436) );
  INV_GATE U13149 ( .I1(n12757), .O(n12758) );
  NAND_GATE U13150 ( .I1(n12762), .I2(n12758), .O(n12770) );
  NAND_GATE U13151 ( .I1(n12760), .I2(n12764), .O(n12768) );
  NAND_GATE U13152 ( .I1(n12762), .I2(n12761), .O(n12763) );
  NAND_GATE U13153 ( .I1(n12764), .I2(n12763), .O(n12765) );
  NAND_GATE U13154 ( .I1(n12766), .I2(n12765), .O(n12767) );
  NAND_GATE U13155 ( .I1(n12768), .I2(n12767), .O(n12769) );
  NAND_GATE U13156 ( .I1(n12770), .I2(n12769), .O(n13422) );
  OR_GATE U13157 ( .I1(n12771), .I2(n12773), .O(n12784) );
  NAND_GATE U13158 ( .I1(n12773), .I2(n12772), .O(n12778) );
  NAND_GATE U13159 ( .I1(n12774), .I2(n12778), .O(n12782) );
  NAND_GATE U13160 ( .I1(n12776), .I2(n12775), .O(n12777) );
  NAND_GATE U13161 ( .I1(n12778), .I2(n12777), .O(n12779) );
  NAND_GATE U13162 ( .I1(n12780), .I2(n12779), .O(n12781) );
  NAND_GATE U13163 ( .I1(n12782), .I2(n12781), .O(n12783) );
  NAND_GATE U13164 ( .I1(n12784), .I2(n12783), .O(n13407) );
  OR_GATE U13165 ( .I1(n12785), .I2(n12789), .O(n12788) );
  OR_GATE U13166 ( .I1(n12786), .I2(n12790), .O(n12787) );
  AND_GATE U13167 ( .I1(n12788), .I2(n12787), .O(n12795) );
  NAND_GATE U13168 ( .I1(n12789), .I2(n1056), .O(n12793) );
  NAND3_GATE U13169 ( .I1(n12793), .I2(n12792), .I3(n12791), .O(n12794) );
  NAND_GATE U13170 ( .I1(n12795), .I2(n12794), .O(n13178) );
  INV_GATE U13171 ( .I1(n13178), .O(n13181) );
  OR_GATE U13172 ( .I1(n12796), .I2(n12798), .O(n12809) );
  NAND_GATE U13173 ( .I1(n12798), .I2(n12797), .O(n12803) );
  NAND_GATE U13174 ( .I1(n12799), .I2(n12803), .O(n12807) );
  NAND_GATE U13175 ( .I1(n12801), .I2(n12800), .O(n12802) );
  NAND_GATE U13176 ( .I1(n12803), .I2(n12802), .O(n12804) );
  NAND_GATE U13177 ( .I1(n12805), .I2(n12804), .O(n12806) );
  NAND_GATE U13178 ( .I1(n12807), .I2(n12806), .O(n12808) );
  NAND_GATE U13179 ( .I1(n12809), .I2(n12808), .O(n13194) );
  OR_GATE U13180 ( .I1(n12810), .I2(n12814), .O(n12813) );
  OR_GATE U13181 ( .I1(n12811), .I2(n12815), .O(n12812) );
  AND_GATE U13182 ( .I1(n12813), .I2(n12812), .O(n12820) );
  NAND_GATE U13183 ( .I1(n12814), .I2(n1067), .O(n12818) );
  NAND3_GATE U13184 ( .I1(n12818), .I2(n12817), .I3(n12816), .O(n12819) );
  NAND_GATE U13185 ( .I1(n12820), .I2(n12819), .O(n13203) );
  INV_GATE U13186 ( .I1(n13203), .O(n13206) );
  OR_GATE U13187 ( .I1(n12821), .I2(n12823), .O(n12834) );
  NAND_GATE U13188 ( .I1(n12823), .I2(n12822), .O(n12828) );
  NAND_GATE U13189 ( .I1(n12824), .I2(n12828), .O(n12832) );
  NAND_GATE U13190 ( .I1(n12826), .I2(n12825), .O(n12827) );
  NAND_GATE U13191 ( .I1(n12828), .I2(n12827), .O(n12829) );
  NAND_GATE U13192 ( .I1(n12830), .I2(n12829), .O(n12831) );
  NAND_GATE U13193 ( .I1(n12832), .I2(n12831), .O(n12833) );
  NAND_GATE U13194 ( .I1(n12834), .I2(n12833), .O(n13219) );
  OR_GATE U13195 ( .I1(n12835), .I2(n12839), .O(n12838) );
  OR_GATE U13196 ( .I1(n12836), .I2(n12840), .O(n12837) );
  AND_GATE U13197 ( .I1(n12838), .I2(n12837), .O(n12845) );
  NAND_GATE U13198 ( .I1(n12839), .I2(n1076), .O(n12843) );
  NAND3_GATE U13199 ( .I1(n12843), .I2(n12842), .I3(n12841), .O(n12844) );
  NAND_GATE U13200 ( .I1(n12845), .I2(n12844), .O(n13228) );
  INV_GATE U13201 ( .I1(n13228), .O(n13231) );
  OR_GATE U13202 ( .I1(n12846), .I2(n12848), .O(n12859) );
  NAND_GATE U13203 ( .I1(n12848), .I2(n12847), .O(n12853) );
  NAND_GATE U13204 ( .I1(n12849), .I2(n12853), .O(n12857) );
  NAND_GATE U13205 ( .I1(n12851), .I2(n12850), .O(n12852) );
  NAND_GATE U13206 ( .I1(n12853), .I2(n12852), .O(n12854) );
  NAND_GATE U13207 ( .I1(n12855), .I2(n12854), .O(n12856) );
  NAND_GATE U13208 ( .I1(n12857), .I2(n12856), .O(n12858) );
  NAND_GATE U13209 ( .I1(n12859), .I2(n12858), .O(n13244) );
  OR_GATE U13210 ( .I1(n12860), .I2(n12864), .O(n12863) );
  OR_GATE U13211 ( .I1(n12861), .I2(n12865), .O(n12862) );
  AND_GATE U13212 ( .I1(n12863), .I2(n12862), .O(n12870) );
  NAND_GATE U13213 ( .I1(n12864), .I2(n1082), .O(n12868) );
  NAND3_GATE U13214 ( .I1(n12868), .I2(n12867), .I3(n12866), .O(n12869) );
  NAND_GATE U13215 ( .I1(n12870), .I2(n12869), .O(n13253) );
  INV_GATE U13216 ( .I1(n13253), .O(n13256) );
  OR_GATE U13217 ( .I1(n12871), .I2(n12873), .O(n12884) );
  NAND_GATE U13218 ( .I1(n12873), .I2(n12872), .O(n12878) );
  NAND_GATE U13219 ( .I1(n12874), .I2(n12878), .O(n12882) );
  NAND_GATE U13220 ( .I1(n12876), .I2(n12875), .O(n12877) );
  NAND_GATE U13221 ( .I1(n12878), .I2(n12877), .O(n12879) );
  NAND_GATE U13222 ( .I1(n12880), .I2(n12879), .O(n12881) );
  NAND_GATE U13223 ( .I1(n12882), .I2(n12881), .O(n12883) );
  NAND_GATE U13224 ( .I1(n12884), .I2(n12883), .O(n13269) );
  OR_GATE U13225 ( .I1(n12885), .I2(n12889), .O(n12888) );
  OR_GATE U13226 ( .I1(n12886), .I2(n12890), .O(n12887) );
  AND_GATE U13227 ( .I1(n12888), .I2(n12887), .O(n12895) );
  NAND_GATE U13228 ( .I1(n12889), .I2(n1088), .O(n12893) );
  NAND3_GATE U13229 ( .I1(n12893), .I2(n12892), .I3(n12891), .O(n12894) );
  NAND_GATE U13230 ( .I1(n12895), .I2(n12894), .O(n13278) );
  INV_GATE U13231 ( .I1(n13278), .O(n13281) );
  OR_GATE U13232 ( .I1(n12896), .I2(n12898), .O(n12909) );
  NAND_GATE U13233 ( .I1(n12898), .I2(n12897), .O(n12903) );
  NAND_GATE U13234 ( .I1(n12899), .I2(n12903), .O(n12907) );
  NAND_GATE U13235 ( .I1(n12901), .I2(n12900), .O(n12902) );
  NAND_GATE U13236 ( .I1(n12903), .I2(n12902), .O(n12904) );
  NAND_GATE U13237 ( .I1(n12905), .I2(n12904), .O(n12906) );
  NAND_GATE U13238 ( .I1(n12907), .I2(n12906), .O(n12908) );
  NAND_GATE U13239 ( .I1(n12909), .I2(n12908), .O(n13294) );
  OR_GATE U13240 ( .I1(n12910), .I2(n12914), .O(n12913) );
  OR_GATE U13241 ( .I1(n12911), .I2(n12915), .O(n12912) );
  AND_GATE U13242 ( .I1(n12913), .I2(n12912), .O(n12920) );
  NAND_GATE U13243 ( .I1(n12914), .I2(n1191), .O(n12918) );
  NAND3_GATE U13244 ( .I1(n12918), .I2(n12917), .I3(n12916), .O(n12919) );
  NAND_GATE U13245 ( .I1(n12920), .I2(n12919), .O(n13303) );
  INV_GATE U13246 ( .I1(n13303), .O(n13306) );
  OR_GATE U13247 ( .I1(n12921), .I2(n12923), .O(n12934) );
  NAND_GATE U13248 ( .I1(n12923), .I2(n12922), .O(n12928) );
  NAND_GATE U13249 ( .I1(n12924), .I2(n12928), .O(n12932) );
  NAND_GATE U13250 ( .I1(n12926), .I2(n12925), .O(n12927) );
  NAND_GATE U13251 ( .I1(n12928), .I2(n12927), .O(n12929) );
  NAND_GATE U13252 ( .I1(n12930), .I2(n12929), .O(n12931) );
  NAND_GATE U13253 ( .I1(n12932), .I2(n12931), .O(n12933) );
  NAND_GATE U13254 ( .I1(n12934), .I2(n12933), .O(n13319) );
  OR_GATE U13255 ( .I1(n12935), .I2(n12939), .O(n12938) );
  OR_GATE U13256 ( .I1(n12936), .I2(n12940), .O(n12937) );
  AND_GATE U13257 ( .I1(n12938), .I2(n12937), .O(n12945) );
  NAND_GATE U13258 ( .I1(n12939), .I2(n1248), .O(n12943) );
  NAND3_GATE U13259 ( .I1(n12943), .I2(n12942), .I3(n12941), .O(n12944) );
  NAND_GATE U13260 ( .I1(n12945), .I2(n12944), .O(n13328) );
  INV_GATE U13261 ( .I1(n13328), .O(n13331) );
  INV_GATE U13262 ( .I1(n12946), .O(n12947) );
  NAND_GATE U13263 ( .I1(n12951), .I2(n12947), .O(n12959) );
  NAND_GATE U13264 ( .I1(n12949), .I2(n12953), .O(n12957) );
  NAND_GATE U13265 ( .I1(n12951), .I2(n12950), .O(n12952) );
  NAND_GATE U13266 ( .I1(n12953), .I2(n12952), .O(n12954) );
  NAND_GATE U13267 ( .I1(n12955), .I2(n12954), .O(n12956) );
  NAND_GATE U13268 ( .I1(n12957), .I2(n12956), .O(n12958) );
  NAND_GATE U13269 ( .I1(n12959), .I2(n12958), .O(n13344) );
  NAND_GATE U13270 ( .I1(n1408), .I2(A[0]), .O(n12960) );
  NAND_GATE U13271 ( .I1(n14241), .I2(n12960), .O(n12961) );
  NAND_GATE U13272 ( .I1(n1410), .I2(n12961), .O(n12965) );
  NAND_GATE U13273 ( .I1(n1411), .I2(A[1]), .O(n12962) );
  NAND_GATE U13274 ( .I1(n724), .I2(n12962), .O(n12963) );
  NAND_GATE U13275 ( .I1(B[4]), .I2(n12963), .O(n12964) );
  NAND_GATE U13276 ( .I1(n12965), .I2(n12964), .O(n13356) );
  NAND_GATE U13277 ( .I1(B[3]), .I2(A[2]), .O(n13360) );
  NAND3_GATE U13278 ( .I1(B[3]), .I2(B[4]), .I3(n1254), .O(n13353) );
  NAND_GATE U13279 ( .I1(n13360), .I2(n13353), .O(n12966) );
  NAND_GATE U13280 ( .I1(n13356), .I2(n12966), .O(n12967) );
  INV_GATE U13281 ( .I1(n13360), .O(n13354) );
  INV_GATE U13282 ( .I1(n13353), .O(n13355) );
  NAND_GATE U13283 ( .I1(n13354), .I2(n13355), .O(n13351) );
  NAND_GATE U13284 ( .I1(n12967), .I2(n13351), .O(n13345) );
  NAND_GATE U13285 ( .I1(n13344), .I2(n13345), .O(n12969) );
  NAND_GATE U13286 ( .I1(B[3]), .I2(A[3]), .O(n13346) );
  INV_GATE U13287 ( .I1(n13346), .O(n12968) );
  NAND_GATE U13288 ( .I1(n13344), .I2(n12968), .O(n13341) );
  NAND_GATE U13289 ( .I1(n13345), .I2(n12968), .O(n13340) );
  NAND3_GATE U13290 ( .I1(n12969), .I2(n13341), .I3(n13340), .O(n13330) );
  INV_GATE U13291 ( .I1(n13330), .O(n13327) );
  NAND_GATE U13292 ( .I1(B[3]), .I2(A[4]), .O(n13335) );
  NAND_GATE U13293 ( .I1(n13327), .I2(n13335), .O(n12970) );
  NAND_GATE U13294 ( .I1(n13331), .I2(n12970), .O(n12971) );
  INV_GATE U13295 ( .I1(n13335), .O(n13329) );
  NAND_GATE U13296 ( .I1(n13330), .I2(n13329), .O(n13326) );
  NAND_GATE U13297 ( .I1(n12971), .I2(n13326), .O(n13320) );
  NAND_GATE U13298 ( .I1(n13319), .I2(n13320), .O(n12973) );
  NAND_GATE U13299 ( .I1(B[3]), .I2(A[5]), .O(n13321) );
  INV_GATE U13300 ( .I1(n13321), .O(n12972) );
  NAND_GATE U13301 ( .I1(n13319), .I2(n12972), .O(n13316) );
  NAND_GATE U13302 ( .I1(n13320), .I2(n12972), .O(n13315) );
  NAND3_GATE U13303 ( .I1(n12973), .I2(n13316), .I3(n13315), .O(n13305) );
  INV_GATE U13304 ( .I1(n13305), .O(n13302) );
  NAND_GATE U13305 ( .I1(B[3]), .I2(A[6]), .O(n13310) );
  NAND_GATE U13306 ( .I1(n13302), .I2(n13310), .O(n12974) );
  NAND_GATE U13307 ( .I1(n13306), .I2(n12974), .O(n12975) );
  INV_GATE U13308 ( .I1(n13310), .O(n13304) );
  NAND_GATE U13309 ( .I1(n13305), .I2(n13304), .O(n13301) );
  NAND_GATE U13310 ( .I1(n12975), .I2(n13301), .O(n13295) );
  NAND_GATE U13311 ( .I1(n13294), .I2(n13295), .O(n12977) );
  NAND_GATE U13312 ( .I1(B[3]), .I2(A[7]), .O(n13296) );
  INV_GATE U13313 ( .I1(n13296), .O(n12976) );
  NAND_GATE U13314 ( .I1(n13294), .I2(n12976), .O(n13291) );
  NAND_GATE U13315 ( .I1(n13295), .I2(n12976), .O(n13290) );
  NAND3_GATE U13316 ( .I1(n12977), .I2(n13291), .I3(n13290), .O(n13280) );
  INV_GATE U13317 ( .I1(n13280), .O(n13277) );
  NAND_GATE U13318 ( .I1(B[3]), .I2(A[8]), .O(n13285) );
  NAND_GATE U13319 ( .I1(n13277), .I2(n13285), .O(n12978) );
  NAND_GATE U13320 ( .I1(n13281), .I2(n12978), .O(n12979) );
  INV_GATE U13321 ( .I1(n13285), .O(n13279) );
  NAND_GATE U13322 ( .I1(n13280), .I2(n13279), .O(n13276) );
  NAND_GATE U13323 ( .I1(n12979), .I2(n13276), .O(n13270) );
  NAND_GATE U13324 ( .I1(n13269), .I2(n13270), .O(n12981) );
  NAND_GATE U13325 ( .I1(B[3]), .I2(A[9]), .O(n13271) );
  INV_GATE U13326 ( .I1(n13271), .O(n12980) );
  NAND_GATE U13327 ( .I1(n13269), .I2(n12980), .O(n13266) );
  NAND_GATE U13328 ( .I1(n13270), .I2(n12980), .O(n13265) );
  NAND3_GATE U13329 ( .I1(n12981), .I2(n13266), .I3(n13265), .O(n13255) );
  INV_GATE U13330 ( .I1(n13255), .O(n13252) );
  NAND_GATE U13331 ( .I1(B[3]), .I2(A[10]), .O(n13260) );
  NAND_GATE U13332 ( .I1(n13252), .I2(n13260), .O(n12982) );
  NAND_GATE U13333 ( .I1(n13256), .I2(n12982), .O(n12983) );
  INV_GATE U13334 ( .I1(n13260), .O(n13254) );
  NAND_GATE U13335 ( .I1(n13255), .I2(n13254), .O(n13251) );
  NAND_GATE U13336 ( .I1(n12983), .I2(n13251), .O(n13245) );
  NAND_GATE U13337 ( .I1(n13244), .I2(n13245), .O(n12985) );
  NAND_GATE U13338 ( .I1(B[3]), .I2(A[11]), .O(n13246) );
  INV_GATE U13339 ( .I1(n13246), .O(n12984) );
  NAND_GATE U13340 ( .I1(n13244), .I2(n12984), .O(n13241) );
  NAND_GATE U13341 ( .I1(n13245), .I2(n12984), .O(n13240) );
  NAND3_GATE U13342 ( .I1(n12985), .I2(n13241), .I3(n13240), .O(n13230) );
  INV_GATE U13343 ( .I1(n13230), .O(n13227) );
  NAND_GATE U13344 ( .I1(B[3]), .I2(A[12]), .O(n13235) );
  NAND_GATE U13345 ( .I1(n13227), .I2(n13235), .O(n12986) );
  NAND_GATE U13346 ( .I1(n13231), .I2(n12986), .O(n12987) );
  INV_GATE U13347 ( .I1(n13235), .O(n13229) );
  NAND_GATE U13348 ( .I1(n13230), .I2(n13229), .O(n13226) );
  NAND_GATE U13349 ( .I1(n12987), .I2(n13226), .O(n13220) );
  NAND_GATE U13350 ( .I1(n13219), .I2(n13220), .O(n12989) );
  NAND_GATE U13351 ( .I1(B[3]), .I2(A[13]), .O(n13221) );
  INV_GATE U13352 ( .I1(n13221), .O(n12988) );
  NAND_GATE U13353 ( .I1(n13219), .I2(n12988), .O(n13216) );
  NAND_GATE U13354 ( .I1(n13220), .I2(n12988), .O(n13215) );
  NAND3_GATE U13355 ( .I1(n12989), .I2(n13216), .I3(n13215), .O(n13205) );
  INV_GATE U13356 ( .I1(n13205), .O(n13202) );
  NAND_GATE U13357 ( .I1(B[3]), .I2(A[14]), .O(n13210) );
  NAND_GATE U13358 ( .I1(n13202), .I2(n13210), .O(n12990) );
  NAND_GATE U13359 ( .I1(n13206), .I2(n12990), .O(n12991) );
  INV_GATE U13360 ( .I1(n13210), .O(n13204) );
  NAND_GATE U13361 ( .I1(n13205), .I2(n13204), .O(n13201) );
  NAND_GATE U13362 ( .I1(n12991), .I2(n13201), .O(n13195) );
  NAND_GATE U13363 ( .I1(n13194), .I2(n13195), .O(n12993) );
  NAND_GATE U13364 ( .I1(B[3]), .I2(A[15]), .O(n13196) );
  INV_GATE U13365 ( .I1(n13196), .O(n12992) );
  NAND_GATE U13366 ( .I1(n13194), .I2(n12992), .O(n13191) );
  NAND_GATE U13367 ( .I1(n13195), .I2(n12992), .O(n13190) );
  NAND3_GATE U13368 ( .I1(n12993), .I2(n13191), .I3(n13190), .O(n13180) );
  INV_GATE U13369 ( .I1(n13180), .O(n13177) );
  NAND_GATE U13370 ( .I1(B[3]), .I2(A[16]), .O(n13185) );
  NAND_GATE U13371 ( .I1(n13177), .I2(n13185), .O(n12994) );
  NAND_GATE U13372 ( .I1(n13181), .I2(n12994), .O(n12995) );
  INV_GATE U13373 ( .I1(n13185), .O(n13179) );
  NAND_GATE U13374 ( .I1(n13180), .I2(n13179), .O(n13176) );
  NAND_GATE U13375 ( .I1(n12995), .I2(n13176), .O(n13408) );
  NAND_GATE U13376 ( .I1(n13407), .I2(n13408), .O(n12997) );
  NAND_GATE U13377 ( .I1(B[3]), .I2(A[17]), .O(n13409) );
  INV_GATE U13378 ( .I1(n13409), .O(n12996) );
  NAND_GATE U13379 ( .I1(n13408), .I2(n12996), .O(n13404) );
  NAND_GATE U13380 ( .I1(n13407), .I2(n12996), .O(n13403) );
  NAND3_GATE U13381 ( .I1(n12997), .I2(n13404), .I3(n13403), .O(n13167) );
  NAND_GATE U13382 ( .I1(B[3]), .I2(A[18]), .O(n13171) );
  OR_GATE U13383 ( .I1(n12998), .I2(n13003), .O(n13001) );
  OR_GATE U13384 ( .I1(n12999), .I2(n13002), .O(n13000) );
  NAND_GATE U13385 ( .I1(n13002), .I2(n1037), .O(n13006) );
  NAND3_GATE U13386 ( .I1(n13006), .I2(n13005), .I3(n13004), .O(n13007) );
  NAND_GATE U13387 ( .I1(n13171), .I2(n13165), .O(n13008) );
  NAND_GATE U13388 ( .I1(n13167), .I2(n13008), .O(n13009) );
  INV_GATE U13389 ( .I1(n13171), .O(n13166) );
  NAND_GATE U13390 ( .I1(n13166), .I2(n136), .O(n13163) );
  NAND_GATE U13391 ( .I1(n13009), .I2(n13163), .O(n13423) );
  NAND_GATE U13392 ( .I1(n13422), .I2(n13423), .O(n13011) );
  NAND_GATE U13393 ( .I1(B[3]), .I2(A[19]), .O(n13424) );
  INV_GATE U13394 ( .I1(n13424), .O(n13010) );
  NAND_GATE U13395 ( .I1(n13423), .I2(n13010), .O(n13419) );
  NAND_GATE U13396 ( .I1(n13422), .I2(n13010), .O(n13418) );
  NAND3_GATE U13397 ( .I1(n13011), .I2(n13419), .I3(n13418), .O(n13156) );
  NAND_GATE U13398 ( .I1(B[3]), .I2(A[20]), .O(n13160) );
  OR_GATE U13399 ( .I1(n13012), .I2(n13017), .O(n13015) );
  OR_GATE U13400 ( .I1(n13013), .I2(n13016), .O(n13014) );
  NAND_GATE U13401 ( .I1(n13016), .I2(n1005), .O(n13020) );
  NAND3_GATE U13402 ( .I1(n13020), .I2(n13019), .I3(n13018), .O(n13021) );
  NAND_GATE U13403 ( .I1(n13160), .I2(n13154), .O(n13022) );
  NAND_GATE U13404 ( .I1(n13156), .I2(n13022), .O(n13023) );
  INV_GATE U13405 ( .I1(n13160), .O(n13155) );
  NAND_GATE U13406 ( .I1(n13155), .I2(n86), .O(n13153) );
  NAND_GATE U13407 ( .I1(n13023), .I2(n13153), .O(n13437) );
  NAND_GATE U13408 ( .I1(n13436), .I2(n13437), .O(n13025) );
  NAND_GATE U13409 ( .I1(B[3]), .I2(A[21]), .O(n13438) );
  INV_GATE U13410 ( .I1(n13438), .O(n13024) );
  NAND_GATE U13411 ( .I1(n13437), .I2(n13024), .O(n13433) );
  NAND_GATE U13412 ( .I1(n13146), .I2(n13148), .O(n13026) );
  NAND_GATE U13413 ( .I1(n13147), .I2(n13026), .O(n13027) );
  NAND_GATE U13414 ( .I1(n13142), .I2(n13027), .O(n13137) );
  NAND_GATE U13415 ( .I1(n13040), .I2(n13137), .O(n13133) );
  INV_GATE U13416 ( .I1(n13028), .O(n13029) );
  NAND_GATE U13417 ( .I1(n13029), .I2(n13033), .O(n13039) );
  NAND_GATE U13418 ( .I1(n13031), .I2(n13030), .O(n13037) );
  NAND_GATE U13419 ( .I1(n13037), .I2(n13036), .O(n13038) );
  NAND_GATE U13420 ( .I1(n13039), .I2(n13038), .O(n13136) );
  NAND_GATE U13421 ( .I1(n13137), .I2(n13136), .O(n13041) );
  NAND_GATE U13422 ( .I1(n13040), .I2(n13136), .O(n13132) );
  NAND3_GATE U13423 ( .I1(n13133), .I2(n13041), .I3(n13132), .O(n13454) );
  NAND_GATE U13424 ( .I1(n13453), .I2(n13456), .O(n13042) );
  NAND_GATE U13425 ( .I1(n13454), .I2(n13042), .O(n13043) );
  NAND_GATE U13426 ( .I1(n13449), .I2(n13043), .O(n13121) );
  INV_GATE U13427 ( .I1(n13044), .O(n13045) );
  NAND_GATE U13428 ( .I1(n13045), .I2(n13047), .O(n13053) );
  NAND3_GATE U13429 ( .I1(n13046), .I2(n13048), .I3(n489), .O(n13051) );
  NAND3_GATE U13430 ( .I1(n13051), .I2(n13050), .I3(n13049), .O(n13052) );
  NAND_GATE U13431 ( .I1(n13053), .I2(n13052), .O(n13122) );
  NAND_GATE U13432 ( .I1(n13121), .I2(n13122), .O(n13055) );
  NAND_GATE U13433 ( .I1(B[3]), .I2(A[25]), .O(n13128) );
  INV_GATE U13434 ( .I1(n13128), .O(n13117) );
  NAND_GATE U13435 ( .I1(n13117), .I2(n13122), .O(n13054) );
  NAND_GATE U13436 ( .I1(n13117), .I2(n13121), .O(n13118) );
  NAND3_GATE U13437 ( .I1(n13055), .I2(n13054), .I3(n13118), .O(n13469) );
  NAND_GATE U13438 ( .I1(n13471), .I2(n13473), .O(n13056) );
  NAND_GATE U13439 ( .I1(n13469), .I2(n13056), .O(n13057) );
  NAND_GATE U13440 ( .I1(n13466), .I2(n13057), .O(n13489) );
  NAND3_GATE U13441 ( .I1(n13058), .I2(n412), .I3(n13489), .O(n13059) );
  NAND_GATE U13442 ( .I1(n13494), .I2(n13489), .O(n13493) );
  NAND_GATE U13443 ( .I1(n13502), .I2(n13504), .O(n13061) );
  NAND_GATE U13444 ( .I1(n13511), .I2(n13061), .O(n13062) );
  NAND_GATE U13445 ( .I1(n13510), .I2(n13062), .O(n13113) );
  NAND_GATE U13446 ( .I1(n13108), .I2(n13113), .O(n13070) );
  NAND_GATE U13447 ( .I1(n399), .I2(n13100), .O(n13065) );
  NAND_GATE U13448 ( .I1(n13102), .I2(n13101), .O(n13064) );
  NAND_GATE U13449 ( .I1(n13065), .I2(n13064), .O(n13066) );
  NAND_GATE U13450 ( .I1(n13103), .I2(n13066), .O(n13099) );
  NAND_GATE U13451 ( .I1(n1016), .I2(n13099), .O(n13069) );
  NAND3_GATE U13452 ( .I1(n13067), .I2(n13099), .I3(n13113), .O(n13068) );
  NAND_GATE U13453 ( .I1(n13518), .I2(n13516), .O(n13071) );
  NAND_GATE U13454 ( .I1(n13523), .I2(n13071), .O(n13072) );
  AND4_GATE U13455 ( .I1(n13077), .I2(n13076), .I3(n13075), .I4(n13074), .O(
        n13090) );
  NAND_GATE U13456 ( .I1(n716), .I2(n13080), .O(n13084) );
  NAND_GATE U13457 ( .I1(n13082), .I2(n13081), .O(n13083) );
  NAND_GATE U13458 ( .I1(n13084), .I2(n13083), .O(n13085) );
  NAND_GATE U13459 ( .I1(n13086), .I2(n13085), .O(n13087) );
  NAND_GATE U13460 ( .I1(n13088), .I2(n13087), .O(n13089) );
  NAND_GATE U13461 ( .I1(n13090), .I2(n13089), .O(n13091) );
  NAND_GATE U13462 ( .I1(n13092), .I2(n13091), .O(n13093) );
  NAND_GATE U13463 ( .I1(n613), .I2(n13093), .O(n13096) );
  INV_GATE U13464 ( .I1(n13093), .O(n14822) );
  NAND_GATE U13465 ( .I1(n13096), .I2(n13095), .O(\A1[33] ) );
  NAND_GATE U13466 ( .I1(n13097), .I2(n604), .O(n13098) );
  NAND_GATE U13467 ( .I1(n13094), .I2(n13098), .O(n13527) );
  NAND_GATE U13468 ( .I1(n1404), .I2(A[30]), .O(n13921) );
  NAND3_GATE U13469 ( .I1(n1016), .I2(n637), .I3(n13099), .O(n13110) );
  NAND3_GATE U13470 ( .I1(n13103), .I2(n13102), .I3(n13101), .O(n13105) );
  NAND3_GATE U13471 ( .I1(n13065), .I2(n13105), .I3(n13104), .O(n13106) );
  NAND_GATE U13472 ( .I1(n13107), .I2(n13106), .O(n13111) );
  NAND3_GATE U13473 ( .I1(n13108), .I2(n13113), .I3(n13112), .O(n13109) );
  NAND_GATE U13474 ( .I1(n13110), .I2(n13109), .O(n13925) );
  NAND_GATE U13475 ( .I1(n637), .I2(n13111), .O(n13116) );
  NAND_GATE U13476 ( .I1(n13113), .I2(n13112), .O(n13115) );
  NAND_GATE U13477 ( .I1(n1404), .I2(A[26]), .O(n13555) );
  INV_GATE U13478 ( .I1(n13555), .O(n13551) );
  INV_GATE U13479 ( .I1(n13121), .O(n13123) );
  NAND3_GATE U13480 ( .I1(n13122), .I2(n13123), .I3(n13117), .O(n13130) );
  INV_GATE U13481 ( .I1(n13118), .O(n13119) );
  INV_GATE U13482 ( .I1(n13122), .O(n13120) );
  NAND_GATE U13483 ( .I1(n13119), .I2(n13120), .O(n13129) );
  AND_GATE U13484 ( .I1(n13130), .I2(n13129), .O(n13125) );
  NAND_GATE U13485 ( .I1(n13121), .I2(n13120), .O(n13127) );
  NAND_GATE U13486 ( .I1(n13123), .I2(n13122), .O(n13126) );
  NAND3_GATE U13487 ( .I1(n13128), .I2(n13127), .I3(n13126), .O(n13124) );
  NAND_GATE U13488 ( .I1(n13125), .I2(n13124), .O(n13550) );
  NAND4_GATE U13489 ( .I1(n13128), .I2(n13127), .I3(n13555), .I4(n13126), .O(
        n13464) );
  NAND_GATE U13490 ( .I1(n13130), .I2(n13129), .O(n13131) );
  NAND_GATE U13491 ( .I1(n13555), .I2(n13131), .O(n13463) );
  OR_GATE U13492 ( .I1(n13132), .I2(n13137), .O(n13135) );
  OR_GATE U13493 ( .I1(n13136), .I2(n13133), .O(n13134) );
  NAND_GATE U13494 ( .I1(n124), .I2(n13136), .O(n13140) );
  NAND3_GATE U13495 ( .I1(n13140), .I2(n13139), .I3(n13138), .O(n13141) );
  INV_GATE U13496 ( .I1(n13894), .O(n13897) );
  NAND_GATE U13497 ( .I1(n1404), .I2(A[24]), .O(n13961) );
  INV_GATE U13498 ( .I1(n13142), .O(n13143) );
  NAND_GATE U13499 ( .I1(n13143), .I2(n13147), .O(n13152) );
  NAND_GATE U13500 ( .I1(n13146), .I2(n1282), .O(n13144) );
  NAND_GATE U13501 ( .I1(n13145), .I2(n13144), .O(n13150) );
  NAND_GATE U13502 ( .I1(n13150), .I2(n13149), .O(n13151) );
  NAND_GATE U13503 ( .I1(n13152), .I2(n13151), .O(n13885) );
  NAND_GATE U13504 ( .I1(n70), .I2(n13154), .O(n13158) );
  NAND_GATE U13505 ( .I1(n13155), .I2(n13158), .O(n13161) );
  NAND_GATE U13506 ( .I1(n13156), .I2(n86), .O(n13157) );
  NAND_GATE U13507 ( .I1(n13158), .I2(n13157), .O(n13159) );
  INV_GATE U13508 ( .I1(n13163), .O(n13164) );
  NAND_GATE U13509 ( .I1(n13167), .I2(n13164), .O(n13175) );
  NAND_GATE U13510 ( .I1(n49), .I2(n13165), .O(n13169) );
  NAND_GATE U13511 ( .I1(n13166), .I2(n13169), .O(n13173) );
  NAND_GATE U13512 ( .I1(n13167), .I2(n136), .O(n13168) );
  NAND_GATE U13513 ( .I1(n13169), .I2(n13168), .O(n13170) );
  NAND_GATE U13514 ( .I1(n13171), .I2(n13170), .O(n13172) );
  NAND_GATE U13515 ( .I1(n13173), .I2(n13172), .O(n13174) );
  NAND_GATE U13516 ( .I1(n13175), .I2(n13174), .O(n13856) );
  OR_GATE U13517 ( .I1(n13176), .I2(n13178), .O(n13189) );
  NAND_GATE U13518 ( .I1(n13178), .I2(n13177), .O(n13183) );
  NAND_GATE U13519 ( .I1(n13179), .I2(n13183), .O(n13187) );
  NAND_GATE U13520 ( .I1(n13181), .I2(n13180), .O(n13182) );
  NAND_GATE U13521 ( .I1(n13183), .I2(n13182), .O(n13184) );
  NAND_GATE U13522 ( .I1(n13185), .I2(n13184), .O(n13186) );
  NAND_GATE U13523 ( .I1(n13187), .I2(n13186), .O(n13188) );
  NAND_GATE U13524 ( .I1(n13189), .I2(n13188), .O(n13841) );
  OR_GATE U13525 ( .I1(n13190), .I2(n13194), .O(n13193) );
  OR_GATE U13526 ( .I1(n13191), .I2(n13195), .O(n13192) );
  AND_GATE U13527 ( .I1(n13193), .I2(n13192), .O(n13200) );
  NAND_GATE U13528 ( .I1(n13194), .I2(n1062), .O(n13198) );
  NAND3_GATE U13529 ( .I1(n13198), .I2(n13197), .I3(n13196), .O(n13199) );
  NAND_GATE U13530 ( .I1(n13200), .I2(n13199), .O(n13612) );
  INV_GATE U13531 ( .I1(n13612), .O(n13615) );
  OR_GATE U13532 ( .I1(n13201), .I2(n13203), .O(n13214) );
  NAND_GATE U13533 ( .I1(n13203), .I2(n13202), .O(n13208) );
  NAND_GATE U13534 ( .I1(n13204), .I2(n13208), .O(n13212) );
  NAND_GATE U13535 ( .I1(n13206), .I2(n13205), .O(n13207) );
  NAND_GATE U13536 ( .I1(n13208), .I2(n13207), .O(n13209) );
  NAND_GATE U13537 ( .I1(n13210), .I2(n13209), .O(n13211) );
  NAND_GATE U13538 ( .I1(n13212), .I2(n13211), .O(n13213) );
  NAND_GATE U13539 ( .I1(n13214), .I2(n13213), .O(n13628) );
  OR_GATE U13540 ( .I1(n13215), .I2(n13219), .O(n13218) );
  OR_GATE U13541 ( .I1(n13216), .I2(n13220), .O(n13217) );
  AND_GATE U13542 ( .I1(n13218), .I2(n13217), .O(n13225) );
  NAND_GATE U13543 ( .I1(n13219), .I2(n1072), .O(n13223) );
  NAND3_GATE U13544 ( .I1(n13223), .I2(n13222), .I3(n13221), .O(n13224) );
  NAND_GATE U13545 ( .I1(n13225), .I2(n13224), .O(n13637) );
  INV_GATE U13546 ( .I1(n13637), .O(n13640) );
  OR_GATE U13547 ( .I1(n13226), .I2(n13228), .O(n13239) );
  NAND_GATE U13548 ( .I1(n13228), .I2(n13227), .O(n13233) );
  NAND_GATE U13549 ( .I1(n13229), .I2(n13233), .O(n13237) );
  NAND_GATE U13550 ( .I1(n13231), .I2(n13230), .O(n13232) );
  NAND_GATE U13551 ( .I1(n13233), .I2(n13232), .O(n13234) );
  NAND_GATE U13552 ( .I1(n13235), .I2(n13234), .O(n13236) );
  NAND_GATE U13553 ( .I1(n13237), .I2(n13236), .O(n13238) );
  NAND_GATE U13554 ( .I1(n13239), .I2(n13238), .O(n13653) );
  OR_GATE U13555 ( .I1(n13240), .I2(n13244), .O(n13243) );
  OR_GATE U13556 ( .I1(n13241), .I2(n13245), .O(n13242) );
  AND_GATE U13557 ( .I1(n13243), .I2(n13242), .O(n13250) );
  NAND_GATE U13558 ( .I1(n13244), .I2(n1078), .O(n13248) );
  NAND3_GATE U13559 ( .I1(n13248), .I2(n13247), .I3(n13246), .O(n13249) );
  NAND_GATE U13560 ( .I1(n13250), .I2(n13249), .O(n13662) );
  INV_GATE U13561 ( .I1(n13662), .O(n13665) );
  OR_GATE U13562 ( .I1(n13251), .I2(n13253), .O(n13264) );
  NAND_GATE U13563 ( .I1(n13253), .I2(n13252), .O(n13258) );
  NAND_GATE U13564 ( .I1(n13254), .I2(n13258), .O(n13262) );
  NAND_GATE U13565 ( .I1(n13256), .I2(n13255), .O(n13257) );
  NAND_GATE U13566 ( .I1(n13258), .I2(n13257), .O(n13259) );
  NAND_GATE U13567 ( .I1(n13260), .I2(n13259), .O(n13261) );
  NAND_GATE U13568 ( .I1(n13262), .I2(n13261), .O(n13263) );
  NAND_GATE U13569 ( .I1(n13264), .I2(n13263), .O(n13678) );
  OR_GATE U13570 ( .I1(n13265), .I2(n13269), .O(n13268) );
  OR_GATE U13571 ( .I1(n13266), .I2(n13270), .O(n13267) );
  AND_GATE U13572 ( .I1(n13268), .I2(n13267), .O(n13275) );
  NAND_GATE U13573 ( .I1(n13269), .I2(n1085), .O(n13273) );
  NAND3_GATE U13574 ( .I1(n13273), .I2(n13272), .I3(n13271), .O(n13274) );
  NAND_GATE U13575 ( .I1(n13275), .I2(n13274), .O(n13687) );
  INV_GATE U13576 ( .I1(n13687), .O(n13690) );
  OR_GATE U13577 ( .I1(n13276), .I2(n13278), .O(n13289) );
  NAND_GATE U13578 ( .I1(n13278), .I2(n13277), .O(n13283) );
  NAND_GATE U13579 ( .I1(n13279), .I2(n13283), .O(n13287) );
  NAND_GATE U13580 ( .I1(n13281), .I2(n13280), .O(n13282) );
  NAND_GATE U13581 ( .I1(n13283), .I2(n13282), .O(n13284) );
  NAND_GATE U13582 ( .I1(n13285), .I2(n13284), .O(n13286) );
  NAND_GATE U13583 ( .I1(n13287), .I2(n13286), .O(n13288) );
  NAND_GATE U13584 ( .I1(n13289), .I2(n13288), .O(n13703) );
  OR_GATE U13585 ( .I1(n13290), .I2(n13294), .O(n13293) );
  OR_GATE U13586 ( .I1(n13291), .I2(n13295), .O(n13292) );
  AND_GATE U13587 ( .I1(n13293), .I2(n13292), .O(n13300) );
  NAND_GATE U13588 ( .I1(n13294), .I2(n1090), .O(n13298) );
  NAND3_GATE U13589 ( .I1(n13298), .I2(n13297), .I3(n13296), .O(n13299) );
  NAND_GATE U13590 ( .I1(n13300), .I2(n13299), .O(n13712) );
  INV_GATE U13591 ( .I1(n13712), .O(n13715) );
  OR_GATE U13592 ( .I1(n13301), .I2(n13303), .O(n13314) );
  NAND_GATE U13593 ( .I1(n13303), .I2(n13302), .O(n13308) );
  NAND_GATE U13594 ( .I1(n13304), .I2(n13308), .O(n13312) );
  NAND_GATE U13595 ( .I1(n13306), .I2(n13305), .O(n13307) );
  NAND_GATE U13596 ( .I1(n13308), .I2(n13307), .O(n13309) );
  NAND_GATE U13597 ( .I1(n13310), .I2(n13309), .O(n13311) );
  NAND_GATE U13598 ( .I1(n13312), .I2(n13311), .O(n13313) );
  NAND_GATE U13599 ( .I1(n13314), .I2(n13313), .O(n13728) );
  OR_GATE U13600 ( .I1(n13315), .I2(n13319), .O(n13318) );
  OR_GATE U13601 ( .I1(n13316), .I2(n13320), .O(n13317) );
  AND_GATE U13602 ( .I1(n13318), .I2(n13317), .O(n13325) );
  NAND_GATE U13603 ( .I1(n13319), .I2(n1193), .O(n13323) );
  NAND3_GATE U13604 ( .I1(n13323), .I2(n13322), .I3(n13321), .O(n13324) );
  NAND_GATE U13605 ( .I1(n13325), .I2(n13324), .O(n13737) );
  INV_GATE U13606 ( .I1(n13737), .O(n13740) );
  OR_GATE U13607 ( .I1(n13326), .I2(n13328), .O(n13339) );
  NAND_GATE U13608 ( .I1(n13328), .I2(n13327), .O(n13333) );
  NAND_GATE U13609 ( .I1(n13329), .I2(n13333), .O(n13337) );
  NAND_GATE U13610 ( .I1(n13331), .I2(n13330), .O(n13332) );
  NAND_GATE U13611 ( .I1(n13333), .I2(n13332), .O(n13334) );
  NAND_GATE U13612 ( .I1(n13335), .I2(n13334), .O(n13336) );
  NAND_GATE U13613 ( .I1(n13337), .I2(n13336), .O(n13338) );
  NAND_GATE U13614 ( .I1(n13339), .I2(n13338), .O(n13753) );
  OR_GATE U13615 ( .I1(n13340), .I2(n13344), .O(n13343) );
  OR_GATE U13616 ( .I1(n13341), .I2(n13345), .O(n13342) );
  AND_GATE U13617 ( .I1(n13343), .I2(n13342), .O(n13350) );
  NAND_GATE U13618 ( .I1(n13344), .I2(n1249), .O(n13348) );
  NAND3_GATE U13619 ( .I1(n13348), .I2(n13347), .I3(n13346), .O(n13349) );
  NAND_GATE U13620 ( .I1(n13350), .I2(n13349), .O(n13762) );
  INV_GATE U13621 ( .I1(n13762), .O(n13765) );
  INV_GATE U13622 ( .I1(n13351), .O(n13352) );
  NAND_GATE U13623 ( .I1(n13356), .I2(n13352), .O(n13364) );
  NAND_GATE U13624 ( .I1(n13354), .I2(n13358), .O(n13362) );
  NAND_GATE U13625 ( .I1(n13356), .I2(n13355), .O(n13357) );
  NAND_GATE U13626 ( .I1(n13358), .I2(n13357), .O(n13359) );
  NAND_GATE U13627 ( .I1(n13360), .I2(n13359), .O(n13361) );
  NAND_GATE U13628 ( .I1(n13362), .I2(n13361), .O(n13363) );
  NAND_GATE U13629 ( .I1(n13364), .I2(n13363), .O(n13778) );
  NAND_GATE U13630 ( .I1(n1407), .I2(A[0]), .O(n13365) );
  NAND_GATE U13631 ( .I1(n14241), .I2(n13365), .O(n13366) );
  NAND_GATE U13632 ( .I1(B[4]), .I2(n13366), .O(n13370) );
  NAND_GATE U13633 ( .I1(n1408), .I2(A[1]), .O(n13367) );
  NAND_GATE U13634 ( .I1(n724), .I2(n13367), .O(n13368) );
  NAND_GATE U13635 ( .I1(B[3]), .I2(n13368), .O(n13369) );
  NAND_GATE U13636 ( .I1(n13370), .I2(n13369), .O(n13790) );
  NAND_GATE U13637 ( .I1(n1404), .I2(A[2]), .O(n13794) );
  NAND3_GATE U13638 ( .I1(n1404), .I2(B[3]), .I3(n1254), .O(n13787) );
  NAND_GATE U13639 ( .I1(n13794), .I2(n13787), .O(n13371) );
  NAND_GATE U13640 ( .I1(n13790), .I2(n13371), .O(n13372) );
  INV_GATE U13641 ( .I1(n13794), .O(n13788) );
  INV_GATE U13642 ( .I1(n13787), .O(n13789) );
  NAND_GATE U13643 ( .I1(n13788), .I2(n13789), .O(n13785) );
  NAND_GATE U13644 ( .I1(n13372), .I2(n13785), .O(n13779) );
  NAND_GATE U13645 ( .I1(n13778), .I2(n13779), .O(n13374) );
  NAND_GATE U13646 ( .I1(n1404), .I2(A[3]), .O(n13780) );
  INV_GATE U13647 ( .I1(n13780), .O(n13373) );
  NAND_GATE U13648 ( .I1(n13778), .I2(n13373), .O(n13775) );
  NAND_GATE U13649 ( .I1(n13779), .I2(n13373), .O(n13774) );
  NAND3_GATE U13650 ( .I1(n13374), .I2(n13775), .I3(n13774), .O(n13764) );
  INV_GATE U13651 ( .I1(n13764), .O(n13761) );
  NAND_GATE U13652 ( .I1(n1404), .I2(A[4]), .O(n13769) );
  NAND_GATE U13653 ( .I1(n13761), .I2(n13769), .O(n13375) );
  NAND_GATE U13654 ( .I1(n13765), .I2(n13375), .O(n13376) );
  INV_GATE U13655 ( .I1(n13769), .O(n13763) );
  NAND_GATE U13656 ( .I1(n13764), .I2(n13763), .O(n13760) );
  NAND_GATE U13657 ( .I1(n13376), .I2(n13760), .O(n13754) );
  NAND_GATE U13658 ( .I1(n13753), .I2(n13754), .O(n13378) );
  NAND_GATE U13659 ( .I1(n1404), .I2(A[5]), .O(n13755) );
  INV_GATE U13660 ( .I1(n13755), .O(n13377) );
  NAND_GATE U13661 ( .I1(n13753), .I2(n13377), .O(n13750) );
  NAND_GATE U13662 ( .I1(n13754), .I2(n13377), .O(n13749) );
  NAND3_GATE U13663 ( .I1(n13378), .I2(n13750), .I3(n13749), .O(n13739) );
  INV_GATE U13664 ( .I1(n13739), .O(n13736) );
  NAND_GATE U13665 ( .I1(n1404), .I2(A[6]), .O(n13744) );
  NAND_GATE U13666 ( .I1(n13736), .I2(n13744), .O(n13379) );
  NAND_GATE U13667 ( .I1(n13740), .I2(n13379), .O(n13380) );
  INV_GATE U13668 ( .I1(n13744), .O(n13738) );
  NAND_GATE U13669 ( .I1(n13739), .I2(n13738), .O(n13735) );
  NAND_GATE U13670 ( .I1(n13380), .I2(n13735), .O(n13729) );
  NAND_GATE U13671 ( .I1(n13728), .I2(n13729), .O(n13382) );
  NAND_GATE U13672 ( .I1(n1405), .I2(A[7]), .O(n13730) );
  INV_GATE U13673 ( .I1(n13730), .O(n13381) );
  NAND_GATE U13674 ( .I1(n13728), .I2(n13381), .O(n13725) );
  NAND_GATE U13675 ( .I1(n13729), .I2(n13381), .O(n13724) );
  NAND3_GATE U13676 ( .I1(n13382), .I2(n13725), .I3(n13724), .O(n13714) );
  INV_GATE U13677 ( .I1(n13714), .O(n13711) );
  NAND_GATE U13678 ( .I1(n1405), .I2(A[8]), .O(n13719) );
  NAND_GATE U13679 ( .I1(n13711), .I2(n13719), .O(n13383) );
  NAND_GATE U13680 ( .I1(n13715), .I2(n13383), .O(n13384) );
  INV_GATE U13681 ( .I1(n13719), .O(n13713) );
  NAND_GATE U13682 ( .I1(n13714), .I2(n13713), .O(n13710) );
  NAND_GATE U13683 ( .I1(n13384), .I2(n13710), .O(n13704) );
  NAND_GATE U13684 ( .I1(n13703), .I2(n13704), .O(n13386) );
  NAND_GATE U13685 ( .I1(n1405), .I2(A[9]), .O(n13705) );
  INV_GATE U13686 ( .I1(n13705), .O(n13385) );
  NAND_GATE U13687 ( .I1(n13703), .I2(n13385), .O(n13700) );
  NAND_GATE U13688 ( .I1(n13704), .I2(n13385), .O(n13699) );
  NAND3_GATE U13689 ( .I1(n13386), .I2(n13700), .I3(n13699), .O(n13689) );
  INV_GATE U13690 ( .I1(n13689), .O(n13686) );
  NAND_GATE U13691 ( .I1(n1405), .I2(A[10]), .O(n13694) );
  NAND_GATE U13692 ( .I1(n13686), .I2(n13694), .O(n13387) );
  NAND_GATE U13693 ( .I1(n13690), .I2(n13387), .O(n13388) );
  INV_GATE U13694 ( .I1(n13694), .O(n13688) );
  NAND_GATE U13695 ( .I1(n13689), .I2(n13688), .O(n13685) );
  NAND_GATE U13696 ( .I1(n13388), .I2(n13685), .O(n13679) );
  NAND_GATE U13697 ( .I1(n13678), .I2(n13679), .O(n13390) );
  NAND_GATE U13698 ( .I1(n1405), .I2(A[11]), .O(n13680) );
  INV_GATE U13699 ( .I1(n13680), .O(n13389) );
  NAND_GATE U13700 ( .I1(n13678), .I2(n13389), .O(n13675) );
  NAND_GATE U13701 ( .I1(n13679), .I2(n13389), .O(n13674) );
  NAND3_GATE U13702 ( .I1(n13390), .I2(n13675), .I3(n13674), .O(n13664) );
  INV_GATE U13703 ( .I1(n13664), .O(n13661) );
  NAND_GATE U13704 ( .I1(n1405), .I2(A[12]), .O(n13669) );
  NAND_GATE U13705 ( .I1(n13661), .I2(n13669), .O(n13391) );
  NAND_GATE U13706 ( .I1(n13665), .I2(n13391), .O(n13392) );
  INV_GATE U13707 ( .I1(n13669), .O(n13663) );
  NAND_GATE U13708 ( .I1(n13664), .I2(n13663), .O(n13660) );
  NAND_GATE U13709 ( .I1(n13392), .I2(n13660), .O(n13654) );
  NAND_GATE U13710 ( .I1(n13653), .I2(n13654), .O(n13394) );
  NAND_GATE U13711 ( .I1(n1405), .I2(A[13]), .O(n13655) );
  INV_GATE U13712 ( .I1(n13655), .O(n13393) );
  NAND_GATE U13713 ( .I1(n13653), .I2(n13393), .O(n13650) );
  NAND_GATE U13714 ( .I1(n13654), .I2(n13393), .O(n13649) );
  NAND3_GATE U13715 ( .I1(n13394), .I2(n13650), .I3(n13649), .O(n13639) );
  INV_GATE U13716 ( .I1(n13639), .O(n13636) );
  NAND_GATE U13717 ( .I1(n1405), .I2(A[14]), .O(n13644) );
  NAND_GATE U13718 ( .I1(n13636), .I2(n13644), .O(n13395) );
  NAND_GATE U13719 ( .I1(n13640), .I2(n13395), .O(n13396) );
  INV_GATE U13720 ( .I1(n13644), .O(n13638) );
  NAND_GATE U13721 ( .I1(n13639), .I2(n13638), .O(n13635) );
  NAND_GATE U13722 ( .I1(n13396), .I2(n13635), .O(n13629) );
  NAND_GATE U13723 ( .I1(n13628), .I2(n13629), .O(n13398) );
  NAND_GATE U13724 ( .I1(n1405), .I2(A[15]), .O(n13630) );
  INV_GATE U13725 ( .I1(n13630), .O(n13397) );
  NAND_GATE U13726 ( .I1(n13628), .I2(n13397), .O(n13625) );
  NAND_GATE U13727 ( .I1(n13629), .I2(n13397), .O(n13624) );
  NAND3_GATE U13728 ( .I1(n13398), .I2(n13625), .I3(n13624), .O(n13614) );
  INV_GATE U13729 ( .I1(n13614), .O(n13611) );
  NAND_GATE U13730 ( .I1(n1405), .I2(A[16]), .O(n13619) );
  NAND_GATE U13731 ( .I1(n13611), .I2(n13619), .O(n13399) );
  NAND_GATE U13732 ( .I1(n13615), .I2(n13399), .O(n13400) );
  INV_GATE U13733 ( .I1(n13619), .O(n13613) );
  NAND_GATE U13734 ( .I1(n13614), .I2(n13613), .O(n13610) );
  NAND_GATE U13735 ( .I1(n13400), .I2(n13610), .O(n13842) );
  NAND_GATE U13736 ( .I1(n13841), .I2(n13842), .O(n13402) );
  NAND_GATE U13737 ( .I1(n1405), .I2(A[17]), .O(n13843) );
  INV_GATE U13738 ( .I1(n13843), .O(n13401) );
  NAND_GATE U13739 ( .I1(n13842), .I2(n13401), .O(n13838) );
  NAND_GATE U13740 ( .I1(n13841), .I2(n13401), .O(n13837) );
  NAND3_GATE U13741 ( .I1(n13402), .I2(n13838), .I3(n13837), .O(n13601) );
  NAND_GATE U13742 ( .I1(n1405), .I2(A[18]), .O(n13605) );
  OR_GATE U13743 ( .I1(n13403), .I2(n13408), .O(n13406) );
  OR_GATE U13744 ( .I1(n13404), .I2(n13407), .O(n13405) );
  AND_GATE U13745 ( .I1(n13406), .I2(n13405), .O(n13413) );
  NAND_GATE U13746 ( .I1(n13407), .I2(n1041), .O(n13411) );
  NAND3_GATE U13747 ( .I1(n13411), .I2(n13410), .I3(n13409), .O(n13412) );
  NAND_GATE U13748 ( .I1(n13413), .I2(n13412), .O(n13597) );
  NAND_GATE U13749 ( .I1(n13605), .I2(n13597), .O(n13414) );
  NAND_GATE U13750 ( .I1(n13601), .I2(n13414), .O(n13415) );
  INV_GATE U13751 ( .I1(n13605), .O(n13599) );
  INV_GATE U13752 ( .I1(n13597), .O(n13600) );
  NAND_GATE U13753 ( .I1(n13599), .I2(n13600), .O(n13595) );
  NAND_GATE U13754 ( .I1(n13415), .I2(n13595), .O(n13857) );
  NAND_GATE U13755 ( .I1(n13856), .I2(n13857), .O(n13417) );
  NAND_GATE U13756 ( .I1(n1405), .I2(A[19]), .O(n13858) );
  INV_GATE U13757 ( .I1(n13858), .O(n13416) );
  NAND_GATE U13758 ( .I1(n13857), .I2(n13416), .O(n13853) );
  NAND_GATE U13759 ( .I1(n13856), .I2(n13416), .O(n13852) );
  NAND3_GATE U13760 ( .I1(n13417), .I2(n13853), .I3(n13852), .O(n13586) );
  NAND_GATE U13761 ( .I1(n1405), .I2(A[20]), .O(n13590) );
  OR_GATE U13762 ( .I1(n13418), .I2(n13423), .O(n13421) );
  OR_GATE U13763 ( .I1(n13419), .I2(n13422), .O(n13420) );
  NAND_GATE U13764 ( .I1(n13422), .I2(n1011), .O(n13426) );
  NAND3_GATE U13765 ( .I1(n13426), .I2(n13425), .I3(n13424), .O(n13427) );
  NAND_GATE U13766 ( .I1(n13590), .I2(n13582), .O(n13428) );
  NAND_GATE U13767 ( .I1(n13586), .I2(n13428), .O(n13429) );
  INV_GATE U13768 ( .I1(n13590), .O(n13584) );
  INV_GATE U13769 ( .I1(n13582), .O(n13585) );
  NAND_GATE U13770 ( .I1(n13584), .I2(n13585), .O(n13580) );
  NAND_GATE U13771 ( .I1(n13429), .I2(n13580), .O(n13872) );
  NAND_GATE U13772 ( .I1(n13871), .I2(n13872), .O(n13431) );
  NAND_GATE U13773 ( .I1(n1405), .I2(A[21]), .O(n13873) );
  INV_GATE U13774 ( .I1(n13873), .O(n13430) );
  NAND_GATE U13775 ( .I1(n13872), .I2(n13430), .O(n13868) );
  NAND_GATE U13776 ( .I1(n13871), .I2(n13430), .O(n13867) );
  NAND3_GATE U13777 ( .I1(n13431), .I2(n13868), .I3(n13867), .O(n13573) );
  NAND_GATE U13778 ( .I1(n1405), .I2(A[22]), .O(n13575) );
  OR_GATE U13779 ( .I1(n13432), .I2(n13437), .O(n13435) );
  OR_GATE U13780 ( .I1(n13433), .I2(n13436), .O(n13434) );
  AND_GATE U13781 ( .I1(n13435), .I2(n13434), .O(n13442) );
  NAND_GATE U13782 ( .I1(n13436), .I2(n1031), .O(n13440) );
  NAND3_GATE U13783 ( .I1(n13440), .I2(n13439), .I3(n13438), .O(n13441) );
  NAND_GATE U13784 ( .I1(n13442), .I2(n13441), .O(n13571) );
  NAND_GATE U13785 ( .I1(n13575), .I2(n13571), .O(n13443) );
  NAND_GATE U13786 ( .I1(n13573), .I2(n13443), .O(n13444) );
  INV_GATE U13787 ( .I1(n13571), .O(n13572) );
  NAND_GATE U13788 ( .I1(n493), .I2(n13572), .O(n13569) );
  NAND_GATE U13789 ( .I1(n13444), .I2(n13569), .O(n13886) );
  NAND_GATE U13790 ( .I1(n13885), .I2(n13886), .O(n13446) );
  NAND_GATE U13791 ( .I1(n1405), .I2(A[23]), .O(n13887) );
  INV_GATE U13792 ( .I1(n13887), .O(n13445) );
  NAND_GATE U13793 ( .I1(n13886), .I2(n13445), .O(n13882) );
  NAND_GATE U13794 ( .I1(n13885), .I2(n13445), .O(n13881) );
  NAND3_GATE U13795 ( .I1(n13446), .I2(n13882), .I3(n13881), .O(n13896) );
  NAND_GATE U13796 ( .I1(n13894), .I2(n13961), .O(n13447) );
  NAND_GATE U13797 ( .I1(n13896), .I2(n13447), .O(n13448) );
  NAND_GATE U13798 ( .I1(n13895), .I2(n13448), .O(n13562) );
  INV_GATE U13799 ( .I1(n13449), .O(n13450) );
  NAND_GATE U13800 ( .I1(n13450), .I2(n13454), .O(n13460) );
  NAND_GATE U13801 ( .I1(n13452), .I2(n13451), .O(n13458) );
  NAND_GATE U13802 ( .I1(n13458), .I2(n13457), .O(n13459) );
  NAND_GATE U13803 ( .I1(n13460), .I2(n13459), .O(n13565) );
  NAND_GATE U13804 ( .I1(n13562), .I2(n13565), .O(n13462) );
  NAND_GATE U13805 ( .I1(n1405), .I2(A[25]), .O(n13559) );
  INV_GATE U13806 ( .I1(n13559), .O(n13461) );
  NAND_GATE U13807 ( .I1(n13461), .I2(n13565), .O(n13563) );
  NAND_GATE U13808 ( .I1(n13461), .I2(n13562), .O(n13564) );
  NAND3_GATE U13809 ( .I1(n13462), .I2(n13563), .I3(n13564), .O(n13553) );
  NAND3_GATE U13810 ( .I1(n13464), .I2(n13463), .I3(n13553), .O(n13465) );
  NAND_GATE U13811 ( .I1(n13549), .I2(n13465), .O(n13540) );
  NAND_GATE U13812 ( .I1(n13471), .I2(n13472), .O(n13467) );
  NAND_GATE U13813 ( .I1(n13468), .I2(n13467), .O(n13476) );
  NAND_GATE U13814 ( .I1(n13470), .I2(n13469), .O(n13475) );
  NAND3_GATE U13815 ( .I1(n13473), .I2(n13472), .I3(n13471), .O(n13474) );
  NAND3_GATE U13816 ( .I1(n13476), .I2(n13475), .I3(n13474), .O(n13477) );
  NAND_GATE U13817 ( .I1(n13478), .I2(n13477), .O(n13545) );
  NAND_GATE U13818 ( .I1(n13540), .I2(n13545), .O(n13481) );
  NAND_GATE U13819 ( .I1(n1405), .I2(A[27]), .O(n13548) );
  INV_GATE U13820 ( .I1(n13548), .O(n13539) );
  NAND_GATE U13821 ( .I1(n13539), .I2(n13545), .O(n13480) );
  NAND_GATE U13822 ( .I1(n13539), .I2(n13540), .O(n13479) );
  NAND3_GATE U13823 ( .I1(n13481), .I2(n13480), .I3(n13479), .O(n13914) );
  NAND_GATE U13824 ( .I1(n1405), .I2(A[28]), .O(n14355) );
  NAND_GATE U13825 ( .I1(n13483), .I2(n13482), .O(n13486) );
  NAND3_GATE U13826 ( .I1(n13486), .I2(n13485), .I3(n13484), .O(n13487) );
  NAND_GATE U13827 ( .I1(n13488), .I2(n13487), .O(n13495) );
  NAND_GATE U13828 ( .I1(n641), .I2(n13495), .O(n13491) );
  NAND3_GATE U13829 ( .I1(n13492), .I2(n13491), .I3(n13490), .O(n13498) );
  OR_GATE U13830 ( .I1(n13495), .I2(n13493), .O(n13497) );
  NAND3_GATE U13831 ( .I1(n641), .I2(n13495), .I3(n13494), .O(n13496) );
  NAND3_GATE U13832 ( .I1(n13498), .I2(n13497), .I3(n13496), .O(n13912) );
  NAND_GATE U13833 ( .I1(n14355), .I2(n13912), .O(n13499) );
  NAND_GATE U13834 ( .I1(n13914), .I2(n13499), .O(n13501) );
  INV_GATE U13835 ( .I1(n14355), .O(n13911) );
  NAND_GATE U13836 ( .I1(n13911), .I2(n573), .O(n13500) );
  NAND_GATE U13837 ( .I1(n13501), .I2(n13500), .O(n13530) );
  NAND3_GATE U13838 ( .I1(n13504), .I2(n615), .I3(n13502), .O(n13509) );
  NAND_GATE U13839 ( .I1(n13503), .I2(n13511), .O(n13508) );
  NAND_GATE U13840 ( .I1(n13504), .I2(n615), .O(n13505) );
  NAND_GATE U13841 ( .I1(n13506), .I2(n13505), .O(n13507) );
  NAND3_GATE U13842 ( .I1(n13509), .I2(n13508), .I3(n13507), .O(n13514) );
  INV_GATE U13843 ( .I1(n13510), .O(n13512) );
  NAND_GATE U13844 ( .I1(n13512), .I2(n13511), .O(n13513) );
  NAND_GATE U13845 ( .I1(n13514), .I2(n13513), .O(n13535) );
  NAND_GATE U13846 ( .I1(n13530), .I2(n13535), .O(n13923) );
  NAND_GATE U13847 ( .I1(n1405), .I2(A[29]), .O(n13533) );
  INV_GATE U13848 ( .I1(n13533), .O(n13534) );
  NAND_GATE U13849 ( .I1(n13534), .I2(n13535), .O(n13924) );
  NAND_GATE U13850 ( .I1(n13534), .I2(n13530), .O(n13926) );
  NAND3_GATE U13851 ( .I1(n13923), .I2(n13924), .I3(n13926), .O(n13930) );
  NAND_GATE U13852 ( .I1(n13921), .I2(n13922), .O(n13515) );
  NAND3_GATE U13853 ( .I1(n13516), .I2(n1387), .I3(n13518), .O(n13521) );
  NAND_GATE U13854 ( .I1(n13517), .I2(n13523), .O(n13520) );
  NAND3_GATE U13855 ( .I1(n13521), .I2(n13520), .I3(n13519), .O(n13526) );
  INV_GATE U13856 ( .I1(n13522), .O(n13524) );
  NAND_GATE U13857 ( .I1(n13524), .I2(n13523), .O(n13525) );
  NAND_GATE U13858 ( .I1(n13526), .I2(n13525), .O(n13931) );
  NAND_GATE U13859 ( .I1(n13932), .I2(n13931), .O(n13934) );
  NAND_GATE U13860 ( .I1(n13527), .I2(n614), .O(n13528) );
  NAND_GATE U13861 ( .I1(n13529), .I2(n13528), .O(\A1[32] ) );
  NAND_GATE U13862 ( .I1(n642), .I2(n13535), .O(n13532) );
  NAND3_GATE U13863 ( .I1(n13533), .I2(n13532), .I3(n13531), .O(n13538) );
  OR_GATE U13864 ( .I1(n13535), .I2(n13926), .O(n13537) );
  NAND3_GATE U13865 ( .I1(n642), .I2(n13535), .I3(n13534), .O(n13536) );
  NAND3_GATE U13866 ( .I1(n13538), .I2(n13537), .I3(n13536), .O(n13940) );
  NAND_GATE U13867 ( .I1(B[1]), .I2(A[30]), .O(n13941) );
  INV_GATE U13868 ( .I1(n13941), .O(n13943) );
  NAND_GATE U13869 ( .I1(n1403), .I2(A[31]), .O(n14371) );
  NAND_GATE U13870 ( .I1(B[1]), .I2(A[29]), .O(n14363) );
  INV_GATE U13871 ( .I1(n14363), .O(n13916) );
  NAND_GATE U13872 ( .I1(n13544), .I2(n1046), .O(n13543) );
  NAND_GATE U13873 ( .I1(n13545), .I2(n1023), .O(n13542) );
  NAND_GATE U13874 ( .I1(n13540), .I2(n13544), .O(n13547) );
  NAND3_GATE U13875 ( .I1(n13548), .I2(n13547), .I3(n13546), .O(n13541) );
  NAND3_GATE U13876 ( .I1(n13543), .I2(n13542), .I3(n13541), .O(n14339) );
  INV_GATE U13877 ( .I1(n14339), .O(n14337) );
  NAND_GATE U13878 ( .I1(B[1]), .I2(A[28]), .O(n14338) );
  INV_GATE U13879 ( .I1(n14338), .O(n14341) );
  NAND3_GATE U13880 ( .I1(n1046), .I2(n13544), .I3(n14338), .O(n13908) );
  NAND3_GATE U13881 ( .I1(n1023), .I2(n13545), .I3(n14338), .O(n13907) );
  NAND4_GATE U13882 ( .I1(n13548), .I2(n13547), .I3(n13546), .I4(n14338), .O(
        n13906) );
  NAND3_GATE U13883 ( .I1(n13552), .I2(n13554), .I3(n13551), .O(n13557) );
  NAND_GATE U13884 ( .I1(n13558), .I2(n13565), .O(n13561) );
  NAND3_GATE U13885 ( .I1(n13561), .I2(n13560), .I3(n13559), .O(n13568) );
  OR_GATE U13886 ( .I1(n13563), .I2(n13562), .O(n13567) );
  OR_GATE U13887 ( .I1(n13565), .I2(n13564), .O(n13566) );
  NAND3_GATE U13888 ( .I1(n13568), .I2(n13567), .I3(n13566), .O(n14326) );
  INV_GATE U13889 ( .I1(n14326), .O(n14328) );
  NAND_GATE U13890 ( .I1(B[1]), .I2(A[26]), .O(n14329) );
  INV_GATE U13891 ( .I1(n14329), .O(n14324) );
  NAND_GATE U13892 ( .I1(n14328), .I2(n14324), .O(n14322) );
  NAND_GATE U13893 ( .I1(B[1]), .I2(A[25]), .O(n13971) );
  INV_GATE U13894 ( .I1(n13971), .O(n13899) );
  INV_GATE U13895 ( .I1(n13569), .O(n13570) );
  NAND_GATE U13896 ( .I1(n13573), .I2(n13570), .O(n13579) );
  NAND_GATE U13897 ( .I1(n493), .I2(n13574), .O(n13577) );
  NAND_GATE U13898 ( .I1(n13577), .I2(n13576), .O(n13578) );
  NAND_GATE U13899 ( .I1(n13579), .I2(n13578), .O(n14295) );
  INV_GATE U13900 ( .I1(n13580), .O(n13581) );
  NAND_GATE U13901 ( .I1(n13586), .I2(n13581), .O(n13594) );
  INV_GATE U13902 ( .I1(n13586), .O(n13583) );
  NAND_GATE U13903 ( .I1(n13583), .I2(n13582), .O(n13588) );
  NAND_GATE U13904 ( .I1(n13584), .I2(n13588), .O(n13592) );
  NAND_GATE U13905 ( .I1(n13588), .I2(n13587), .O(n13589) );
  NAND_GATE U13906 ( .I1(n13590), .I2(n13589), .O(n13591) );
  NAND_GATE U13907 ( .I1(n13592), .I2(n13591), .O(n13593) );
  NAND_GATE U13908 ( .I1(n13594), .I2(n13593), .O(n13992) );
  INV_GATE U13909 ( .I1(n13595), .O(n13596) );
  NAND_GATE U13910 ( .I1(n13601), .I2(n13596), .O(n13609) );
  INV_GATE U13911 ( .I1(n13601), .O(n13598) );
  NAND_GATE U13912 ( .I1(n13598), .I2(n13597), .O(n13603) );
  NAND_GATE U13913 ( .I1(n13599), .I2(n13603), .O(n13607) );
  NAND_GATE U13914 ( .I1(n13601), .I2(n13600), .O(n13602) );
  NAND_GATE U13915 ( .I1(n13603), .I2(n13602), .O(n13604) );
  NAND_GATE U13916 ( .I1(n13605), .I2(n13604), .O(n13606) );
  NAND_GATE U13917 ( .I1(n13607), .I2(n13606), .O(n13608) );
  NAND_GATE U13918 ( .I1(n13609), .I2(n13608), .O(n14018) );
  OR_GATE U13919 ( .I1(n13610), .I2(n13612), .O(n13623) );
  NAND_GATE U13920 ( .I1(n13612), .I2(n13611), .O(n13617) );
  NAND_GATE U13921 ( .I1(n13613), .I2(n13617), .O(n13621) );
  NAND_GATE U13922 ( .I1(n13615), .I2(n13614), .O(n13616) );
  NAND_GATE U13923 ( .I1(n13617), .I2(n13616), .O(n13618) );
  NAND_GATE U13924 ( .I1(n13619), .I2(n13618), .O(n13620) );
  NAND_GATE U13925 ( .I1(n13621), .I2(n13620), .O(n13622) );
  NAND_GATE U13926 ( .I1(n13623), .I2(n13622), .O(n14044) );
  OR_GATE U13927 ( .I1(n13624), .I2(n13628), .O(n13627) );
  OR_GATE U13928 ( .I1(n13625), .I2(n13629), .O(n13626) );
  AND_GATE U13929 ( .I1(n13627), .I2(n13626), .O(n13634) );
  NAND_GATE U13930 ( .I1(n13628), .I2(n1068), .O(n13632) );
  NAND3_GATE U13931 ( .I1(n13632), .I2(n13631), .I3(n13630), .O(n13633) );
  NAND_GATE U13932 ( .I1(n13634), .I2(n13633), .O(n14053) );
  INV_GATE U13933 ( .I1(n14053), .O(n14056) );
  OR_GATE U13934 ( .I1(n13635), .I2(n13637), .O(n13648) );
  NAND_GATE U13935 ( .I1(n13637), .I2(n13636), .O(n13642) );
  NAND_GATE U13936 ( .I1(n13638), .I2(n13642), .O(n13646) );
  NAND_GATE U13937 ( .I1(n13640), .I2(n13639), .O(n13641) );
  NAND_GATE U13938 ( .I1(n13642), .I2(n13641), .O(n13643) );
  NAND_GATE U13939 ( .I1(n13644), .I2(n13643), .O(n13645) );
  NAND_GATE U13940 ( .I1(n13646), .I2(n13645), .O(n13647) );
  NAND_GATE U13941 ( .I1(n13648), .I2(n13647), .O(n14069) );
  OR_GATE U13942 ( .I1(n13649), .I2(n13653), .O(n13652) );
  OR_GATE U13943 ( .I1(n13650), .I2(n13654), .O(n13651) );
  AND_GATE U13944 ( .I1(n13652), .I2(n13651), .O(n13659) );
  NAND_GATE U13945 ( .I1(n13653), .I2(n1077), .O(n13657) );
  NAND3_GATE U13946 ( .I1(n13657), .I2(n13656), .I3(n13655), .O(n13658) );
  NAND_GATE U13947 ( .I1(n13659), .I2(n13658), .O(n14078) );
  INV_GATE U13948 ( .I1(n14078), .O(n14081) );
  OR_GATE U13949 ( .I1(n13660), .I2(n13662), .O(n13673) );
  NAND_GATE U13950 ( .I1(n13662), .I2(n13661), .O(n13667) );
  NAND_GATE U13951 ( .I1(n13663), .I2(n13667), .O(n13671) );
  NAND_GATE U13952 ( .I1(n13665), .I2(n13664), .O(n13666) );
  NAND_GATE U13953 ( .I1(n13667), .I2(n13666), .O(n13668) );
  NAND_GATE U13954 ( .I1(n13669), .I2(n13668), .O(n13670) );
  NAND_GATE U13955 ( .I1(n13671), .I2(n13670), .O(n13672) );
  NAND_GATE U13956 ( .I1(n13673), .I2(n13672), .O(n14094) );
  OR_GATE U13957 ( .I1(n13674), .I2(n13678), .O(n13677) );
  OR_GATE U13958 ( .I1(n13675), .I2(n13679), .O(n13676) );
  AND_GATE U13959 ( .I1(n13677), .I2(n13676), .O(n13684) );
  NAND_GATE U13960 ( .I1(n13678), .I2(n1084), .O(n13682) );
  NAND3_GATE U13961 ( .I1(n13682), .I2(n13681), .I3(n13680), .O(n13683) );
  NAND_GATE U13962 ( .I1(n13684), .I2(n13683), .O(n14103) );
  INV_GATE U13963 ( .I1(n14103), .O(n14106) );
  OR_GATE U13964 ( .I1(n13685), .I2(n13687), .O(n13698) );
  NAND_GATE U13965 ( .I1(n13687), .I2(n13686), .O(n13692) );
  NAND_GATE U13966 ( .I1(n13688), .I2(n13692), .O(n13696) );
  NAND_GATE U13967 ( .I1(n13690), .I2(n13689), .O(n13691) );
  NAND_GATE U13968 ( .I1(n13692), .I2(n13691), .O(n13693) );
  NAND_GATE U13969 ( .I1(n13694), .I2(n13693), .O(n13695) );
  NAND_GATE U13970 ( .I1(n13696), .I2(n13695), .O(n13697) );
  NAND_GATE U13971 ( .I1(n13698), .I2(n13697), .O(n14119) );
  OR_GATE U13972 ( .I1(n13699), .I2(n13703), .O(n13702) );
  OR_GATE U13973 ( .I1(n13700), .I2(n13704), .O(n13701) );
  AND_GATE U13974 ( .I1(n13702), .I2(n13701), .O(n13709) );
  NAND_GATE U13975 ( .I1(n13703), .I2(n1089), .O(n13707) );
  NAND3_GATE U13976 ( .I1(n13707), .I2(n13706), .I3(n13705), .O(n13708) );
  NAND_GATE U13977 ( .I1(n13709), .I2(n13708), .O(n14128) );
  INV_GATE U13978 ( .I1(n14128), .O(n14131) );
  OR_GATE U13979 ( .I1(n13710), .I2(n13712), .O(n13723) );
  NAND_GATE U13980 ( .I1(n13712), .I2(n13711), .O(n13717) );
  NAND_GATE U13981 ( .I1(n13713), .I2(n13717), .O(n13721) );
  NAND_GATE U13982 ( .I1(n13715), .I2(n13714), .O(n13716) );
  NAND_GATE U13983 ( .I1(n13717), .I2(n13716), .O(n13718) );
  NAND_GATE U13984 ( .I1(n13719), .I2(n13718), .O(n13720) );
  NAND_GATE U13985 ( .I1(n13721), .I2(n13720), .O(n13722) );
  NAND_GATE U13986 ( .I1(n13723), .I2(n13722), .O(n14144) );
  OR_GATE U13987 ( .I1(n13724), .I2(n13728), .O(n13727) );
  OR_GATE U13988 ( .I1(n13725), .I2(n13729), .O(n13726) );
  AND_GATE U13989 ( .I1(n13727), .I2(n13726), .O(n13734) );
  NAND_GATE U13990 ( .I1(n13728), .I2(n1092), .O(n13732) );
  NAND3_GATE U13991 ( .I1(n13732), .I2(n13731), .I3(n13730), .O(n13733) );
  NAND_GATE U13992 ( .I1(n13734), .I2(n13733), .O(n14153) );
  INV_GATE U13993 ( .I1(n14153), .O(n14156) );
  OR_GATE U13994 ( .I1(n13735), .I2(n13737), .O(n13748) );
  NAND_GATE U13995 ( .I1(n13737), .I2(n13736), .O(n13742) );
  NAND_GATE U13996 ( .I1(n13738), .I2(n13742), .O(n13746) );
  NAND_GATE U13997 ( .I1(n13740), .I2(n13739), .O(n13741) );
  NAND_GATE U13998 ( .I1(n13742), .I2(n13741), .O(n13743) );
  NAND_GATE U13999 ( .I1(n13744), .I2(n13743), .O(n13745) );
  NAND_GATE U14000 ( .I1(n13746), .I2(n13745), .O(n13747) );
  NAND_GATE U14001 ( .I1(n13748), .I2(n13747), .O(n14169) );
  OR_GATE U14002 ( .I1(n13749), .I2(n13753), .O(n13752) );
  OR_GATE U14003 ( .I1(n13750), .I2(n13754), .O(n13751) );
  AND_GATE U14004 ( .I1(n13752), .I2(n13751), .O(n13759) );
  NAND_GATE U14005 ( .I1(n13753), .I2(n1195), .O(n13757) );
  NAND3_GATE U14006 ( .I1(n13757), .I2(n13756), .I3(n13755), .O(n13758) );
  NAND_GATE U14007 ( .I1(n13759), .I2(n13758), .O(n14178) );
  INV_GATE U14008 ( .I1(n14178), .O(n14181) );
  OR_GATE U14009 ( .I1(n13760), .I2(n13762), .O(n13773) );
  NAND_GATE U14010 ( .I1(n13762), .I2(n13761), .O(n13767) );
  NAND_GATE U14011 ( .I1(n13763), .I2(n13767), .O(n13771) );
  NAND_GATE U14012 ( .I1(n13765), .I2(n13764), .O(n13766) );
  NAND_GATE U14013 ( .I1(n13767), .I2(n13766), .O(n13768) );
  NAND_GATE U14014 ( .I1(n13769), .I2(n13768), .O(n13770) );
  NAND_GATE U14015 ( .I1(n13771), .I2(n13770), .O(n13772) );
  NAND_GATE U14016 ( .I1(n13773), .I2(n13772), .O(n14194) );
  OR_GATE U14017 ( .I1(n13774), .I2(n13778), .O(n13777) );
  OR_GATE U14018 ( .I1(n13775), .I2(n13779), .O(n13776) );
  AND_GATE U14019 ( .I1(n13777), .I2(n13776), .O(n13784) );
  NAND_GATE U14020 ( .I1(n13778), .I2(n1250), .O(n13782) );
  NAND3_GATE U14021 ( .I1(n13782), .I2(n13781), .I3(n13780), .O(n13783) );
  NAND_GATE U14022 ( .I1(n13784), .I2(n13783), .O(n14203) );
  INV_GATE U14023 ( .I1(n14203), .O(n14206) );
  INV_GATE U14024 ( .I1(n13785), .O(n13786) );
  NAND_GATE U14025 ( .I1(n13790), .I2(n13786), .O(n13798) );
  NAND_GATE U14026 ( .I1(n13788), .I2(n13792), .O(n13796) );
  NAND_GATE U14027 ( .I1(n13790), .I2(n13789), .O(n13791) );
  NAND_GATE U14028 ( .I1(n13792), .I2(n13791), .O(n13793) );
  NAND_GATE U14029 ( .I1(n13794), .I2(n13793), .O(n13795) );
  NAND_GATE U14030 ( .I1(n13796), .I2(n13795), .O(n13797) );
  NAND_GATE U14031 ( .I1(n13798), .I2(n13797), .O(n14219) );
  NAND_GATE U14032 ( .I1(n1406), .I2(A[0]), .O(n13799) );
  NAND_GATE U14033 ( .I1(n14241), .I2(n13799), .O(n13800) );
  NAND_GATE U14034 ( .I1(B[3]), .I2(n13800), .O(n13804) );
  NAND_GATE U14035 ( .I1(n1407), .I2(A[1]), .O(n13801) );
  NAND_GATE U14036 ( .I1(n724), .I2(n13801), .O(n13802) );
  NAND_GATE U14037 ( .I1(n1405), .I2(n13802), .O(n13803) );
  NAND_GATE U14038 ( .I1(n13804), .I2(n13803), .O(n14231) );
  NAND_GATE U14039 ( .I1(B[1]), .I2(A[2]), .O(n14235) );
  NAND3_GATE U14040 ( .I1(B[1]), .I2(n1405), .I3(n1254), .O(n14228) );
  NAND_GATE U14041 ( .I1(n14235), .I2(n14228), .O(n13805) );
  NAND_GATE U14042 ( .I1(n14231), .I2(n13805), .O(n13806) );
  INV_GATE U14043 ( .I1(n14235), .O(n14229) );
  INV_GATE U14044 ( .I1(n14228), .O(n14230) );
  NAND_GATE U14045 ( .I1(n14229), .I2(n14230), .O(n14226) );
  NAND_GATE U14046 ( .I1(n13806), .I2(n14226), .O(n14220) );
  NAND_GATE U14047 ( .I1(n14219), .I2(n14220), .O(n13808) );
  NAND_GATE U14048 ( .I1(B[1]), .I2(A[3]), .O(n14221) );
  INV_GATE U14049 ( .I1(n14221), .O(n13807) );
  NAND_GATE U14050 ( .I1(n14219), .I2(n13807), .O(n14216) );
  NAND_GATE U14051 ( .I1(n14220), .I2(n13807), .O(n14215) );
  NAND3_GATE U14052 ( .I1(n13808), .I2(n14216), .I3(n14215), .O(n14205) );
  INV_GATE U14053 ( .I1(n14205), .O(n14202) );
  NAND_GATE U14054 ( .I1(B[1]), .I2(A[4]), .O(n14210) );
  NAND_GATE U14055 ( .I1(n14202), .I2(n14210), .O(n13809) );
  NAND_GATE U14056 ( .I1(n14206), .I2(n13809), .O(n13810) );
  INV_GATE U14057 ( .I1(n14210), .O(n14204) );
  NAND_GATE U14058 ( .I1(n14205), .I2(n14204), .O(n14201) );
  NAND_GATE U14059 ( .I1(n13810), .I2(n14201), .O(n14195) );
  NAND_GATE U14060 ( .I1(n14194), .I2(n14195), .O(n13812) );
  NAND_GATE U14061 ( .I1(B[1]), .I2(A[5]), .O(n14196) );
  INV_GATE U14062 ( .I1(n14196), .O(n13811) );
  NAND_GATE U14063 ( .I1(n14194), .I2(n13811), .O(n14191) );
  NAND_GATE U14064 ( .I1(n14195), .I2(n13811), .O(n14190) );
  NAND3_GATE U14065 ( .I1(n13812), .I2(n14191), .I3(n14190), .O(n14180) );
  INV_GATE U14066 ( .I1(n14180), .O(n14177) );
  NAND_GATE U14067 ( .I1(B[1]), .I2(A[6]), .O(n14185) );
  NAND_GATE U14068 ( .I1(n14177), .I2(n14185), .O(n13813) );
  NAND_GATE U14069 ( .I1(n14181), .I2(n13813), .O(n13814) );
  INV_GATE U14070 ( .I1(n14185), .O(n14179) );
  NAND_GATE U14071 ( .I1(n14180), .I2(n14179), .O(n14176) );
  NAND_GATE U14072 ( .I1(n13814), .I2(n14176), .O(n14170) );
  NAND_GATE U14073 ( .I1(n14169), .I2(n14170), .O(n13816) );
  NAND_GATE U14074 ( .I1(B[1]), .I2(A[7]), .O(n14171) );
  INV_GATE U14075 ( .I1(n14171), .O(n13815) );
  NAND_GATE U14076 ( .I1(n14169), .I2(n13815), .O(n14166) );
  NAND_GATE U14077 ( .I1(n14170), .I2(n13815), .O(n14165) );
  NAND3_GATE U14078 ( .I1(n13816), .I2(n14166), .I3(n14165), .O(n14155) );
  INV_GATE U14079 ( .I1(n14155), .O(n14152) );
  NAND_GATE U14080 ( .I1(B[1]), .I2(A[8]), .O(n14160) );
  NAND_GATE U14081 ( .I1(n14152), .I2(n14160), .O(n13817) );
  NAND_GATE U14082 ( .I1(n14156), .I2(n13817), .O(n13818) );
  INV_GATE U14083 ( .I1(n14160), .O(n14154) );
  NAND_GATE U14084 ( .I1(n14155), .I2(n14154), .O(n14151) );
  NAND_GATE U14085 ( .I1(n13818), .I2(n14151), .O(n14145) );
  NAND_GATE U14086 ( .I1(n14144), .I2(n14145), .O(n13820) );
  NAND_GATE U14087 ( .I1(B[1]), .I2(A[9]), .O(n14146) );
  INV_GATE U14088 ( .I1(n14146), .O(n13819) );
  NAND_GATE U14089 ( .I1(n14144), .I2(n13819), .O(n14141) );
  NAND_GATE U14090 ( .I1(n14145), .I2(n13819), .O(n14140) );
  NAND3_GATE U14091 ( .I1(n13820), .I2(n14141), .I3(n14140), .O(n14130) );
  INV_GATE U14092 ( .I1(n14130), .O(n14127) );
  NAND_GATE U14093 ( .I1(B[1]), .I2(A[10]), .O(n14135) );
  NAND_GATE U14094 ( .I1(n14127), .I2(n14135), .O(n13821) );
  NAND_GATE U14095 ( .I1(n14131), .I2(n13821), .O(n13822) );
  INV_GATE U14096 ( .I1(n14135), .O(n14129) );
  NAND_GATE U14097 ( .I1(n14130), .I2(n14129), .O(n14126) );
  NAND_GATE U14098 ( .I1(n13822), .I2(n14126), .O(n14120) );
  NAND_GATE U14099 ( .I1(n14119), .I2(n14120), .O(n13824) );
  NAND_GATE U14100 ( .I1(B[1]), .I2(A[11]), .O(n14121) );
  INV_GATE U14101 ( .I1(n14121), .O(n13823) );
  NAND_GATE U14102 ( .I1(n14119), .I2(n13823), .O(n14116) );
  NAND_GATE U14103 ( .I1(n14120), .I2(n13823), .O(n14115) );
  NAND3_GATE U14104 ( .I1(n13824), .I2(n14116), .I3(n14115), .O(n14105) );
  INV_GATE U14105 ( .I1(n14105), .O(n14102) );
  NAND_GATE U14106 ( .I1(B[1]), .I2(A[12]), .O(n14110) );
  NAND_GATE U14107 ( .I1(n14102), .I2(n14110), .O(n13825) );
  NAND_GATE U14108 ( .I1(n14106), .I2(n13825), .O(n13826) );
  INV_GATE U14109 ( .I1(n14110), .O(n14104) );
  NAND_GATE U14110 ( .I1(n14105), .I2(n14104), .O(n14101) );
  NAND_GATE U14111 ( .I1(n13826), .I2(n14101), .O(n14095) );
  NAND_GATE U14112 ( .I1(n14094), .I2(n14095), .O(n13828) );
  NAND_GATE U14113 ( .I1(B[1]), .I2(A[13]), .O(n14096) );
  INV_GATE U14114 ( .I1(n14096), .O(n13827) );
  NAND_GATE U14115 ( .I1(n14094), .I2(n13827), .O(n14091) );
  NAND_GATE U14116 ( .I1(n14095), .I2(n13827), .O(n14090) );
  NAND3_GATE U14117 ( .I1(n13828), .I2(n14091), .I3(n14090), .O(n14080) );
  INV_GATE U14118 ( .I1(n14080), .O(n14077) );
  NAND_GATE U14119 ( .I1(B[1]), .I2(A[14]), .O(n14085) );
  NAND_GATE U14120 ( .I1(n14077), .I2(n14085), .O(n13829) );
  NAND_GATE U14121 ( .I1(n14081), .I2(n13829), .O(n13830) );
  INV_GATE U14122 ( .I1(n14085), .O(n14079) );
  NAND_GATE U14123 ( .I1(n14080), .I2(n14079), .O(n14076) );
  NAND_GATE U14124 ( .I1(n13830), .I2(n14076), .O(n14070) );
  NAND_GATE U14125 ( .I1(n14069), .I2(n14070), .O(n13832) );
  NAND_GATE U14126 ( .I1(B[1]), .I2(A[15]), .O(n14071) );
  INV_GATE U14127 ( .I1(n14071), .O(n13831) );
  NAND_GATE U14128 ( .I1(n14069), .I2(n13831), .O(n14066) );
  NAND_GATE U14129 ( .I1(n14070), .I2(n13831), .O(n14065) );
  NAND3_GATE U14130 ( .I1(n13832), .I2(n14066), .I3(n14065), .O(n14055) );
  INV_GATE U14131 ( .I1(n14055), .O(n14052) );
  NAND_GATE U14132 ( .I1(B[1]), .I2(A[16]), .O(n14060) );
  NAND_GATE U14133 ( .I1(n14052), .I2(n14060), .O(n13833) );
  NAND_GATE U14134 ( .I1(n14056), .I2(n13833), .O(n13834) );
  INV_GATE U14135 ( .I1(n14060), .O(n14054) );
  NAND_GATE U14136 ( .I1(n14055), .I2(n14054), .O(n14051) );
  NAND_GATE U14137 ( .I1(n13834), .I2(n14051), .O(n14045) );
  NAND_GATE U14138 ( .I1(n14044), .I2(n14045), .O(n13836) );
  NAND_GATE U14139 ( .I1(B[1]), .I2(A[17]), .O(n14046) );
  INV_GATE U14140 ( .I1(n14046), .O(n13835) );
  NAND_GATE U14141 ( .I1(n14045), .I2(n13835), .O(n14041) );
  NAND3_GATE U14142 ( .I1(n13836), .I2(n14041), .I3(n14040), .O(n14031) );
  NAND_GATE U14143 ( .I1(B[1]), .I2(A[18]), .O(n14035) );
  OR_GATE U14144 ( .I1(n13837), .I2(n13842), .O(n13840) );
  OR_GATE U14145 ( .I1(n13838), .I2(n13841), .O(n13839) );
  AND_GATE U14146 ( .I1(n13840), .I2(n13839), .O(n13847) );
  NAND_GATE U14147 ( .I1(n13841), .I2(n1055), .O(n13845) );
  NAND3_GATE U14148 ( .I1(n13845), .I2(n13844), .I3(n13843), .O(n13846) );
  NAND_GATE U14149 ( .I1(n13847), .I2(n13846), .O(n14027) );
  NAND_GATE U14150 ( .I1(n14035), .I2(n14027), .O(n13848) );
  NAND_GATE U14151 ( .I1(n14031), .I2(n13848), .O(n13849) );
  INV_GATE U14152 ( .I1(n14035), .O(n14029) );
  INV_GATE U14153 ( .I1(n14027), .O(n14030) );
  NAND_GATE U14154 ( .I1(n14029), .I2(n14030), .O(n14025) );
  NAND_GATE U14155 ( .I1(n13849), .I2(n14025), .O(n14019) );
  NAND_GATE U14156 ( .I1(n14018), .I2(n14019), .O(n13851) );
  NAND_GATE U14157 ( .I1(B[1]), .I2(A[19]), .O(n14020) );
  INV_GATE U14158 ( .I1(n14020), .O(n13850) );
  NAND_GATE U14159 ( .I1(n14019), .I2(n13850), .O(n14015) );
  NAND_GATE U14160 ( .I1(n14018), .I2(n13850), .O(n14014) );
  NAND3_GATE U14161 ( .I1(n13851), .I2(n14015), .I3(n14014), .O(n14005) );
  NAND_GATE U14162 ( .I1(B[1]), .I2(A[20]), .O(n14009) );
  OR_GATE U14163 ( .I1(n13852), .I2(n13857), .O(n13855) );
  OR_GATE U14164 ( .I1(n13853), .I2(n13856), .O(n13854) );
  AND_GATE U14165 ( .I1(n13855), .I2(n13854), .O(n13862) );
  NAND_GATE U14166 ( .I1(n13856), .I2(n1049), .O(n13860) );
  NAND3_GATE U14167 ( .I1(n13860), .I2(n13859), .I3(n13858), .O(n13861) );
  NAND_GATE U14168 ( .I1(n13862), .I2(n13861), .O(n14001) );
  NAND_GATE U14169 ( .I1(n14009), .I2(n14001), .O(n13863) );
  NAND_GATE U14170 ( .I1(n14005), .I2(n13863), .O(n13864) );
  INV_GATE U14171 ( .I1(n14009), .O(n14003) );
  INV_GATE U14172 ( .I1(n14001), .O(n14004) );
  NAND_GATE U14173 ( .I1(n14003), .I2(n14004), .O(n13999) );
  NAND_GATE U14174 ( .I1(n13864), .I2(n13999), .O(n13993) );
  NAND_GATE U14175 ( .I1(n13992), .I2(n13993), .O(n13866) );
  NAND_GATE U14176 ( .I1(B[1]), .I2(A[21]), .O(n13994) );
  INV_GATE U14177 ( .I1(n13994), .O(n13865) );
  NAND_GATE U14178 ( .I1(n13993), .I2(n13865), .O(n13989) );
  NAND_GATE U14179 ( .I1(n13992), .I2(n13865), .O(n13988) );
  NAND3_GATE U14180 ( .I1(n13866), .I2(n13989), .I3(n13988), .O(n13981) );
  NAND_GATE U14181 ( .I1(B[1]), .I2(A[22]), .O(n13983) );
  OR_GATE U14182 ( .I1(n13867), .I2(n13872), .O(n13870) );
  OR_GATE U14183 ( .I1(n13868), .I2(n13871), .O(n13869) );
  NAND_GATE U14184 ( .I1(n13871), .I2(n1009), .O(n13875) );
  NAND3_GATE U14185 ( .I1(n13875), .I2(n13874), .I3(n13873), .O(n13876) );
  NAND_GATE U14186 ( .I1(n13983), .I2(n13978), .O(n13877) );
  NAND_GATE U14187 ( .I1(n13981), .I2(n13877), .O(n13878) );
  INV_GATE U14188 ( .I1(n13983), .O(n13979) );
  INV_GATE U14189 ( .I1(n13978), .O(n13980) );
  NAND_GATE U14190 ( .I1(n13979), .I2(n13980), .O(n13976) );
  NAND_GATE U14191 ( .I1(n13878), .I2(n13976), .O(n14296) );
  NAND_GATE U14192 ( .I1(n14295), .I2(n14296), .O(n13880) );
  NAND_GATE U14193 ( .I1(B[1]), .I2(A[23]), .O(n14297) );
  INV_GATE U14194 ( .I1(n14297), .O(n13879) );
  NAND_GATE U14195 ( .I1(n14296), .I2(n13879), .O(n14292) );
  NAND_GATE U14196 ( .I1(n14295), .I2(n13879), .O(n14291) );
  NAND3_GATE U14197 ( .I1(n13880), .I2(n14292), .I3(n14291), .O(n14310) );
  NAND_GATE U14198 ( .I1(B[1]), .I2(A[24]), .O(n14313) );
  OR_GATE U14199 ( .I1(n13881), .I2(n13886), .O(n13884) );
  OR_GATE U14200 ( .I1(n13882), .I2(n13885), .O(n13883) );
  NAND_GATE U14201 ( .I1(n13885), .I2(n491), .O(n13889) );
  NAND3_GATE U14202 ( .I1(n13889), .I2(n13888), .I3(n13887), .O(n13890) );
  NAND_GATE U14203 ( .I1(n14313), .I2(n14307), .O(n13891) );
  NAND_GATE U14204 ( .I1(n14310), .I2(n13891), .O(n13892) );
  INV_GATE U14205 ( .I1(n14313), .O(n14306) );
  INV_GATE U14206 ( .I1(n14307), .O(n14309) );
  NAND_GATE U14207 ( .I1(n14306), .I2(n14309), .O(n14303) );
  NAND_GATE U14208 ( .I1(n13892), .I2(n14303), .O(n13970) );
  NAND_GATE U14209 ( .I1(n13899), .I2(n13970), .O(n13966) );
  INV_GATE U14210 ( .I1(n13896), .O(n13893) );
  NAND_GATE U14211 ( .I1(n13894), .I2(n13893), .O(n13898) );
  NAND_GATE U14212 ( .I1(n418), .I2(n13898), .O(n13963) );
  NAND3_GATE U14213 ( .I1(n13899), .I2(n13900), .I3(n13962), .O(n13960) );
  NAND3_GATE U14214 ( .I1(n13970), .I2(n13900), .I3(n13962), .O(n13901) );
  NAND3_GATE U14215 ( .I1(n13966), .I2(n13960), .I3(n13901), .O(n14327) );
  NAND_GATE U14216 ( .I1(n14326), .I2(n14329), .O(n13902) );
  NAND_GATE U14217 ( .I1(n14327), .I2(n13902), .O(n13903) );
  NAND_GATE U14218 ( .I1(n14322), .I2(n13903), .O(n13956) );
  NAND_GATE U14219 ( .I1(B[1]), .I2(A[27]), .O(n13952) );
  INV_GATE U14220 ( .I1(n13952), .O(n13904) );
  NAND_GATE U14221 ( .I1(n13904), .I2(n13956), .O(n13953) );
  NAND3_GATE U14222 ( .I1(n13905), .I2(n13953), .I3(n13955), .O(n14346) );
  NAND4_GATE U14223 ( .I1(n13908), .I2(n13907), .I3(n13906), .I4(n14346), .O(
        n13909) );
  NAND_GATE U14224 ( .I1(n14345), .I2(n13909), .O(n14362) );
  NAND_GATE U14225 ( .I1(n13916), .I2(n14362), .O(n14358) );
  INV_GATE U14226 ( .I1(n13914), .O(n13913) );
  NAND_GATE U14227 ( .I1(n13913), .I2(n13912), .O(n13910) );
  NAND_GATE U14228 ( .I1(n13911), .I2(n13910), .O(n14356) );
  NAND3_GATE U14229 ( .I1(n573), .I2(n13911), .I3(n13914), .O(n14357) );
  NAND_GATE U14230 ( .I1(n13914), .I2(n573), .O(n13915) );
  NAND_GATE U14231 ( .I1(n13910), .I2(n13915), .O(n14354) );
  NAND_GATE U14232 ( .I1(n14355), .I2(n14354), .O(n13918) );
  NAND3_GATE U14233 ( .I1(n13916), .I2(n13917), .I3(n13918), .O(n14353) );
  NAND3_GATE U14234 ( .I1(n13918), .I2(n13917), .I3(n14362), .O(n13919) );
  NAND3_GATE U14235 ( .I1(n14358), .I2(n14353), .I3(n13919), .O(n13942) );
  NAND_GATE U14236 ( .I1(n13940), .I2(n13941), .O(n13920) );
  NAND_GATE U14237 ( .I1(n13942), .I2(n13920), .O(n14370) );
  NAND3_GATE U14238 ( .I1(n14372), .I2(n14371), .I3(n14370), .O(n14825) );
  NAND3_GATE U14239 ( .I1(n13922), .I2(n1274), .I3(n13921), .O(n13928) );
  NAND3_GATE U14240 ( .I1(n13929), .I2(n13928), .I3(n13927), .O(n14369) );
  NAND_GATE U14241 ( .I1(n1399), .I2(n13930), .O(n14373) );
  NAND_GATE U14242 ( .I1(n14369), .I2(n14373), .O(n14824) );
  NAND_GATE U14243 ( .I1(n14825), .I2(n14824), .O(n14375) );
  OR_GATE U14244 ( .I1(n13932), .I2(n13931), .O(n13933) );
  NAND_GATE U14245 ( .I1(n13934), .I2(n13933), .O(n13935) );
  NAND_GATE U14246 ( .I1(n639), .I2(n13935), .O(n13937) );
  NAND_GATE U14247 ( .I1(n14375), .I2(n14823), .O(n13936) );
  NAND_GATE U14248 ( .I1(n13937), .I2(n13936), .O(\A1[31] ) );
  INV_GATE U14249 ( .I1(n14372), .O(n13938) );
  NAND_GATE U14250 ( .I1(n13938), .I2(n13942), .O(n13949) );
  NAND_GATE U14251 ( .I1(n13939), .I2(n13943), .O(n13947) );
  NAND_GATE U14252 ( .I1(n13939), .I2(n13942), .O(n13946) );
  NAND_GATE U14253 ( .I1(n13943), .I2(n13942), .O(n13944) );
  NAND4_GATE U14254 ( .I1(n13947), .I2(n13946), .I3(n13945), .I4(n13944), .O(
        n13948) );
  NAND_GATE U14255 ( .I1(n13949), .I2(n13948), .O(n14827) );
  NAND_GATE U14256 ( .I1(A[30]), .I2(n1401), .O(n14392) );
  NAND_GATE U14257 ( .I1(n13954), .I2(n13956), .O(n13950) );
  NAND3_GATE U14258 ( .I1(n13952), .I2(n13951), .I3(n13950), .O(n13959) );
  OR_GATE U14259 ( .I1(n13956), .I2(n13955), .O(n13957) );
  NAND_GATE U14260 ( .I1(A[28]), .I2(n1401), .O(n14416) );
  NAND_GATE U14261 ( .I1(A[27]), .I2(n1401), .O(n14425) );
  INV_GATE U14262 ( .I1(n14425), .O(n14422) );
  OR_GATE U14263 ( .I1(n13960), .I2(n13970), .O(n13968) );
  NAND_GATE U14264 ( .I1(n13963), .I2(n13962), .O(n13964) );
  NAND_GATE U14265 ( .I1(n13965), .I2(n13964), .O(n13969) );
  OR_GATE U14266 ( .I1(n13969), .I2(n13966), .O(n13967) );
  AND_GATE U14267 ( .I1(n13968), .I2(n13967), .O(n13975) );
  NAND_GATE U14268 ( .I1(n1004), .I2(n13969), .O(n13973) );
  NAND3_GATE U14269 ( .I1(n13973), .I2(n13972), .I3(n13971), .O(n13974) );
  NAND_GATE U14270 ( .I1(n13975), .I2(n13974), .O(n14439) );
  NAND_GATE U14271 ( .I1(A[25]), .I2(n1401), .O(n14447) );
  NAND_GATE U14272 ( .I1(A[24]), .I2(n1401), .O(n14460) );
  INV_GATE U14273 ( .I1(n14460), .O(n14455) );
  INV_GATE U14274 ( .I1(n13976), .O(n13977) );
  NAND_GATE U14275 ( .I1(n13981), .I2(n13977), .O(n13987) );
  NAND_GATE U14276 ( .I1(n13979), .I2(n13982), .O(n13985) );
  NAND_GATE U14277 ( .I1(n13985), .I2(n13984), .O(n13986) );
  NAND_GATE U14278 ( .I1(n13987), .I2(n13986), .O(n14479) );
  OR_GATE U14279 ( .I1(n13989), .I2(n13992), .O(n13990) );
  AND_GATE U14280 ( .I1(n13991), .I2(n13990), .O(n13998) );
  NAND_GATE U14281 ( .I1(n13992), .I2(n1050), .O(n13996) );
  NAND3_GATE U14282 ( .I1(n13996), .I2(n13995), .I3(n13994), .O(n13997) );
  NAND_GATE U14283 ( .I1(n13998), .I2(n13997), .O(n14490) );
  INV_GATE U14284 ( .I1(n14490), .O(n14483) );
  INV_GATE U14285 ( .I1(n13999), .O(n14000) );
  NAND_GATE U14286 ( .I1(n14005), .I2(n14000), .O(n14013) );
  INV_GATE U14287 ( .I1(n14005), .O(n14002) );
  NAND_GATE U14288 ( .I1(n14002), .I2(n14001), .O(n14007) );
  NAND_GATE U14289 ( .I1(n14003), .I2(n14007), .O(n14011) );
  NAND_GATE U14290 ( .I1(n14007), .I2(n14006), .O(n14008) );
  NAND_GATE U14291 ( .I1(n14009), .I2(n14008), .O(n14010) );
  NAND_GATE U14292 ( .I1(n14011), .I2(n14010), .O(n14012) );
  NAND_GATE U14293 ( .I1(n14013), .I2(n14012), .O(n14505) );
  OR_GATE U14294 ( .I1(n14014), .I2(n14019), .O(n14017) );
  OR_GATE U14295 ( .I1(n14015), .I2(n14018), .O(n14016) );
  AND_GATE U14296 ( .I1(n14017), .I2(n14016), .O(n14024) );
  NAND_GATE U14297 ( .I1(n14018), .I2(n1045), .O(n14022) );
  NAND3_GATE U14298 ( .I1(n14022), .I2(n14021), .I3(n14020), .O(n14023) );
  NAND_GATE U14299 ( .I1(n14024), .I2(n14023), .O(n14517) );
  INV_GATE U14300 ( .I1(n14517), .O(n14510) );
  INV_GATE U14301 ( .I1(n14025), .O(n14026) );
  NAND_GATE U14302 ( .I1(n14031), .I2(n14026), .O(n14039) );
  INV_GATE U14303 ( .I1(n14031), .O(n14028) );
  NAND_GATE U14304 ( .I1(n14028), .I2(n14027), .O(n14033) );
  NAND_GATE U14305 ( .I1(n14029), .I2(n14033), .O(n14037) );
  NAND_GATE U14306 ( .I1(n14031), .I2(n14030), .O(n14032) );
  NAND_GATE U14307 ( .I1(n14033), .I2(n14032), .O(n14034) );
  NAND_GATE U14308 ( .I1(n14035), .I2(n14034), .O(n14036) );
  NAND_GATE U14309 ( .I1(n14037), .I2(n14036), .O(n14038) );
  NAND_GATE U14310 ( .I1(n14039), .I2(n14038), .O(n14533) );
  OR_GATE U14311 ( .I1(n14040), .I2(n14045), .O(n14043) );
  OR_GATE U14312 ( .I1(n14041), .I2(n14044), .O(n14042) );
  AND_GATE U14313 ( .I1(n14043), .I2(n14042), .O(n14050) );
  NAND_GATE U14314 ( .I1(n14044), .I2(n1063), .O(n14048) );
  NAND3_GATE U14315 ( .I1(n14048), .I2(n14047), .I3(n14046), .O(n14049) );
  NAND_GATE U14316 ( .I1(n14050), .I2(n14049), .O(n14546) );
  INV_GATE U14317 ( .I1(n14546), .O(n14539) );
  OR_GATE U14318 ( .I1(n14051), .I2(n14053), .O(n14064) );
  NAND_GATE U14319 ( .I1(n14053), .I2(n14052), .O(n14058) );
  NAND_GATE U14320 ( .I1(n14054), .I2(n14058), .O(n14062) );
  NAND_GATE U14321 ( .I1(n14056), .I2(n14055), .O(n14057) );
  NAND_GATE U14322 ( .I1(n14058), .I2(n14057), .O(n14059) );
  NAND_GATE U14323 ( .I1(n14060), .I2(n14059), .O(n14061) );
  NAND_GATE U14324 ( .I1(n14062), .I2(n14061), .O(n14063) );
  NAND_GATE U14325 ( .I1(n14064), .I2(n14063), .O(n14562) );
  OR_GATE U14326 ( .I1(n14065), .I2(n14069), .O(n14068) );
  OR_GATE U14327 ( .I1(n14066), .I2(n14070), .O(n14067) );
  AND_GATE U14328 ( .I1(n14068), .I2(n14067), .O(n14075) );
  NAND_GATE U14329 ( .I1(n14069), .I2(n1073), .O(n14073) );
  NAND3_GATE U14330 ( .I1(n14073), .I2(n14072), .I3(n14071), .O(n14074) );
  NAND_GATE U14331 ( .I1(n14075), .I2(n14074), .O(n14575) );
  INV_GATE U14332 ( .I1(n14575), .O(n14568) );
  OR_GATE U14333 ( .I1(n14076), .I2(n14078), .O(n14089) );
  NAND_GATE U14334 ( .I1(n14078), .I2(n14077), .O(n14083) );
  NAND_GATE U14335 ( .I1(n14079), .I2(n14083), .O(n14087) );
  NAND_GATE U14336 ( .I1(n14081), .I2(n14080), .O(n14082) );
  NAND_GATE U14337 ( .I1(n14083), .I2(n14082), .O(n14084) );
  NAND_GATE U14338 ( .I1(n14085), .I2(n14084), .O(n14086) );
  NAND_GATE U14339 ( .I1(n14087), .I2(n14086), .O(n14088) );
  NAND_GATE U14340 ( .I1(n14089), .I2(n14088), .O(n14591) );
  OR_GATE U14341 ( .I1(n14090), .I2(n14094), .O(n14093) );
  OR_GATE U14342 ( .I1(n14091), .I2(n14095), .O(n14092) );
  AND_GATE U14343 ( .I1(n14093), .I2(n14092), .O(n14100) );
  NAND_GATE U14344 ( .I1(n14094), .I2(n1081), .O(n14098) );
  NAND3_GATE U14345 ( .I1(n14098), .I2(n14097), .I3(n14096), .O(n14099) );
  NAND_GATE U14346 ( .I1(n14100), .I2(n14099), .O(n14604) );
  INV_GATE U14347 ( .I1(n14604), .O(n14597) );
  OR_GATE U14348 ( .I1(n14101), .I2(n14103), .O(n14114) );
  NAND_GATE U14349 ( .I1(n14103), .I2(n14102), .O(n14108) );
  NAND_GATE U14350 ( .I1(n14104), .I2(n14108), .O(n14112) );
  NAND_GATE U14351 ( .I1(n14106), .I2(n14105), .O(n14107) );
  NAND_GATE U14352 ( .I1(n14108), .I2(n14107), .O(n14109) );
  NAND_GATE U14353 ( .I1(n14110), .I2(n14109), .O(n14111) );
  NAND_GATE U14354 ( .I1(n14112), .I2(n14111), .O(n14113) );
  NAND_GATE U14355 ( .I1(n14114), .I2(n14113), .O(n14620) );
  OR_GATE U14356 ( .I1(n14115), .I2(n14119), .O(n14118) );
  OR_GATE U14357 ( .I1(n14116), .I2(n14120), .O(n14117) );
  AND_GATE U14358 ( .I1(n14118), .I2(n14117), .O(n14125) );
  NAND_GATE U14359 ( .I1(n14119), .I2(n1087), .O(n14123) );
  NAND3_GATE U14360 ( .I1(n14123), .I2(n14122), .I3(n14121), .O(n14124) );
  NAND_GATE U14361 ( .I1(n14125), .I2(n14124), .O(n14633) );
  INV_GATE U14362 ( .I1(n14633), .O(n14626) );
  OR_GATE U14363 ( .I1(n14126), .I2(n14128), .O(n14139) );
  NAND_GATE U14364 ( .I1(n14128), .I2(n14127), .O(n14133) );
  NAND_GATE U14365 ( .I1(n14129), .I2(n14133), .O(n14137) );
  NAND_GATE U14366 ( .I1(n14131), .I2(n14130), .O(n14132) );
  NAND_GATE U14367 ( .I1(n14133), .I2(n14132), .O(n14134) );
  NAND_GATE U14368 ( .I1(n14135), .I2(n14134), .O(n14136) );
  NAND_GATE U14369 ( .I1(n14137), .I2(n14136), .O(n14138) );
  NAND_GATE U14370 ( .I1(n14139), .I2(n14138), .O(n14649) );
  OR_GATE U14371 ( .I1(n14140), .I2(n14144), .O(n14143) );
  OR_GATE U14372 ( .I1(n14141), .I2(n14145), .O(n14142) );
  AND_GATE U14373 ( .I1(n14143), .I2(n14142), .O(n14150) );
  NAND_GATE U14374 ( .I1(n14144), .I2(n1091), .O(n14148) );
  NAND3_GATE U14375 ( .I1(n14148), .I2(n14147), .I3(n14146), .O(n14149) );
  NAND_GATE U14376 ( .I1(n14150), .I2(n14149), .O(n14662) );
  INV_GATE U14377 ( .I1(n14662), .O(n14655) );
  OR_GATE U14378 ( .I1(n14151), .I2(n14153), .O(n14164) );
  NAND_GATE U14379 ( .I1(n14153), .I2(n14152), .O(n14158) );
  NAND_GATE U14380 ( .I1(n14154), .I2(n14158), .O(n14162) );
  NAND_GATE U14381 ( .I1(n14156), .I2(n14155), .O(n14157) );
  NAND_GATE U14382 ( .I1(n14158), .I2(n14157), .O(n14159) );
  NAND_GATE U14383 ( .I1(n14160), .I2(n14159), .O(n14161) );
  NAND_GATE U14384 ( .I1(n14162), .I2(n14161), .O(n14163) );
  NAND_GATE U14385 ( .I1(n14164), .I2(n14163), .O(n14678) );
  OR_GATE U14386 ( .I1(n14165), .I2(n14169), .O(n14168) );
  OR_GATE U14387 ( .I1(n14166), .I2(n14170), .O(n14167) );
  AND_GATE U14388 ( .I1(n14168), .I2(n14167), .O(n14175) );
  NAND_GATE U14389 ( .I1(n14169), .I2(n1093), .O(n14173) );
  NAND3_GATE U14390 ( .I1(n14173), .I2(n14172), .I3(n14171), .O(n14174) );
  NAND_GATE U14391 ( .I1(n14175), .I2(n14174), .O(n14691) );
  INV_GATE U14392 ( .I1(n14691), .O(n14684) );
  OR_GATE U14393 ( .I1(n14176), .I2(n14178), .O(n14189) );
  NAND_GATE U14394 ( .I1(n14178), .I2(n14177), .O(n14183) );
  NAND_GATE U14395 ( .I1(n14179), .I2(n14183), .O(n14187) );
  NAND_GATE U14396 ( .I1(n14181), .I2(n14180), .O(n14182) );
  NAND_GATE U14397 ( .I1(n14183), .I2(n14182), .O(n14184) );
  NAND_GATE U14398 ( .I1(n14185), .I2(n14184), .O(n14186) );
  NAND_GATE U14399 ( .I1(n14187), .I2(n14186), .O(n14188) );
  NAND_GATE U14400 ( .I1(n14189), .I2(n14188), .O(n14707) );
  OR_GATE U14401 ( .I1(n14190), .I2(n14194), .O(n14193) );
  OR_GATE U14402 ( .I1(n14191), .I2(n14195), .O(n14192) );
  AND_GATE U14403 ( .I1(n14193), .I2(n14192), .O(n14200) );
  NAND_GATE U14404 ( .I1(n14194), .I2(n1196), .O(n14198) );
  NAND3_GATE U14405 ( .I1(n14198), .I2(n14197), .I3(n14196), .O(n14199) );
  NAND_GATE U14406 ( .I1(n14200), .I2(n14199), .O(n14720) );
  INV_GATE U14407 ( .I1(n14720), .O(n14713) );
  OR_GATE U14408 ( .I1(n14201), .I2(n14203), .O(n14214) );
  NAND_GATE U14409 ( .I1(n14203), .I2(n14202), .O(n14208) );
  NAND_GATE U14410 ( .I1(n14204), .I2(n14208), .O(n14212) );
  NAND_GATE U14411 ( .I1(n14206), .I2(n14205), .O(n14207) );
  NAND_GATE U14412 ( .I1(n14208), .I2(n14207), .O(n14209) );
  NAND_GATE U14413 ( .I1(n14210), .I2(n14209), .O(n14211) );
  NAND_GATE U14414 ( .I1(n14212), .I2(n14211), .O(n14213) );
  NAND_GATE U14415 ( .I1(n14214), .I2(n14213), .O(n14736) );
  OR_GATE U14416 ( .I1(n14215), .I2(n14219), .O(n14218) );
  OR_GATE U14417 ( .I1(n14216), .I2(n14220), .O(n14217) );
  AND_GATE U14418 ( .I1(n14218), .I2(n14217), .O(n14225) );
  NAND_GATE U14419 ( .I1(n14219), .I2(n1251), .O(n14223) );
  NAND3_GATE U14420 ( .I1(n14223), .I2(n14222), .I3(n14221), .O(n14224) );
  NAND_GATE U14421 ( .I1(n14225), .I2(n14224), .O(n14749) );
  INV_GATE U14422 ( .I1(n14749), .O(n14742) );
  INV_GATE U14423 ( .I1(n14226), .O(n14227) );
  NAND_GATE U14424 ( .I1(n14231), .I2(n14227), .O(n14239) );
  NAND_GATE U14425 ( .I1(n14229), .I2(n14233), .O(n14237) );
  NAND_GATE U14426 ( .I1(n14231), .I2(n14230), .O(n14232) );
  NAND_GATE U14427 ( .I1(n14233), .I2(n14232), .O(n14234) );
  NAND_GATE U14428 ( .I1(n14235), .I2(n14234), .O(n14236) );
  NAND_GATE U14429 ( .I1(n14237), .I2(n14236), .O(n14238) );
  NAND_GATE U14430 ( .I1(n14239), .I2(n14238), .O(n14765) );
  NAND3_GATE U14431 ( .I1(B[1]), .I2(B[0]), .I3(n1254), .O(n14778) );
  INV_GATE U14432 ( .I1(n14778), .O(n14771) );
  NAND_GATE U14433 ( .I1(n1403), .I2(A[0]), .O(n14240) );
  NAND_GATE U14434 ( .I1(n14241), .I2(n14240), .O(n14242) );
  NAND_GATE U14435 ( .I1(n1405), .I2(n14242), .O(n14246) );
  NAND_GATE U14436 ( .I1(n1406), .I2(A[1]), .O(n14243) );
  NAND_GATE U14437 ( .I1(n724), .I2(n14243), .O(n14244) );
  NAND_GATE U14438 ( .I1(B[1]), .I2(n14244), .O(n14245) );
  NAND_GATE U14439 ( .I1(n14246), .I2(n14245), .O(n14770) );
  INV_GATE U14440 ( .I1(n14770), .O(n14768) );
  NAND_GATE U14441 ( .I1(A[2]), .I2(B[0]), .O(n14775) );
  NAND_GATE U14442 ( .I1(n14768), .I2(n14775), .O(n14247) );
  NAND_GATE U14443 ( .I1(n14771), .I2(n14247), .O(n14248) );
  INV_GATE U14444 ( .I1(n14775), .O(n14769) );
  NAND_GATE U14445 ( .I1(n14770), .I2(n14769), .O(n14779) );
  NAND_GATE U14446 ( .I1(n14248), .I2(n14779), .O(n14755) );
  INV_GATE U14447 ( .I1(n14755), .O(n14757) );
  NAND_GATE U14448 ( .I1(A[3]), .I2(n1401), .O(n14760) );
  NAND_GATE U14449 ( .I1(n14757), .I2(n14760), .O(n14249) );
  NAND_GATE U14450 ( .I1(n14765), .I2(n14249), .O(n14250) );
  INV_GATE U14451 ( .I1(n14760), .O(n14754) );
  NAND_GATE U14452 ( .I1(n14755), .I2(n14754), .O(n14763) );
  NAND_GATE U14453 ( .I1(n14250), .I2(n14763), .O(n14741) );
  INV_GATE U14454 ( .I1(n14741), .O(n14739) );
  NAND_GATE U14455 ( .I1(A[4]), .I2(n1401), .O(n14746) );
  NAND_GATE U14456 ( .I1(n14739), .I2(n14746), .O(n14251) );
  NAND_GATE U14457 ( .I1(n14742), .I2(n14251), .O(n14252) );
  INV_GATE U14458 ( .I1(n14746), .O(n14740) );
  NAND_GATE U14459 ( .I1(n14741), .I2(n14740), .O(n14750) );
  NAND_GATE U14460 ( .I1(n14252), .I2(n14750), .O(n14726) );
  INV_GATE U14461 ( .I1(n14726), .O(n14728) );
  NAND_GATE U14462 ( .I1(A[5]), .I2(n1401), .O(n14731) );
  NAND_GATE U14463 ( .I1(n14728), .I2(n14731), .O(n14253) );
  NAND_GATE U14464 ( .I1(n14736), .I2(n14253), .O(n14254) );
  INV_GATE U14465 ( .I1(n14731), .O(n14725) );
  NAND_GATE U14466 ( .I1(n14726), .I2(n14725), .O(n14734) );
  NAND_GATE U14467 ( .I1(n14254), .I2(n14734), .O(n14712) );
  INV_GATE U14468 ( .I1(n14712), .O(n14710) );
  NAND_GATE U14469 ( .I1(A[6]), .I2(n1401), .O(n14717) );
  NAND_GATE U14470 ( .I1(n14710), .I2(n14717), .O(n14255) );
  NAND_GATE U14471 ( .I1(n14713), .I2(n14255), .O(n14256) );
  INV_GATE U14472 ( .I1(n14717), .O(n14711) );
  NAND_GATE U14473 ( .I1(n14712), .I2(n14711), .O(n14721) );
  NAND_GATE U14474 ( .I1(n14256), .I2(n14721), .O(n14697) );
  INV_GATE U14475 ( .I1(n14697), .O(n14699) );
  NAND_GATE U14476 ( .I1(A[7]), .I2(n1401), .O(n14702) );
  NAND_GATE U14477 ( .I1(n14699), .I2(n14702), .O(n14257) );
  NAND_GATE U14478 ( .I1(n14707), .I2(n14257), .O(n14258) );
  INV_GATE U14479 ( .I1(n14702), .O(n14696) );
  NAND_GATE U14480 ( .I1(n14697), .I2(n14696), .O(n14705) );
  NAND_GATE U14481 ( .I1(n14258), .I2(n14705), .O(n14683) );
  INV_GATE U14482 ( .I1(n14683), .O(n14681) );
  NAND_GATE U14483 ( .I1(A[8]), .I2(n1401), .O(n14688) );
  NAND_GATE U14484 ( .I1(n14681), .I2(n14688), .O(n14259) );
  NAND_GATE U14485 ( .I1(n14684), .I2(n14259), .O(n14260) );
  INV_GATE U14486 ( .I1(n14688), .O(n14682) );
  NAND_GATE U14487 ( .I1(n14683), .I2(n14682), .O(n14692) );
  NAND_GATE U14488 ( .I1(n14260), .I2(n14692), .O(n14668) );
  INV_GATE U14489 ( .I1(n14668), .O(n14670) );
  NAND_GATE U14490 ( .I1(A[9]), .I2(n1401), .O(n14673) );
  NAND_GATE U14491 ( .I1(n14670), .I2(n14673), .O(n14261) );
  NAND_GATE U14492 ( .I1(n14678), .I2(n14261), .O(n14262) );
  INV_GATE U14493 ( .I1(n14673), .O(n14667) );
  NAND_GATE U14494 ( .I1(n14668), .I2(n14667), .O(n14676) );
  NAND_GATE U14495 ( .I1(n14262), .I2(n14676), .O(n14654) );
  INV_GATE U14496 ( .I1(n14654), .O(n14652) );
  NAND_GATE U14497 ( .I1(A[10]), .I2(n1401), .O(n14659) );
  NAND_GATE U14498 ( .I1(n14652), .I2(n14659), .O(n14263) );
  NAND_GATE U14499 ( .I1(n14655), .I2(n14263), .O(n14264) );
  INV_GATE U14500 ( .I1(n14659), .O(n14653) );
  NAND_GATE U14501 ( .I1(n14654), .I2(n14653), .O(n14663) );
  NAND_GATE U14502 ( .I1(n14264), .I2(n14663), .O(n14639) );
  INV_GATE U14503 ( .I1(n14639), .O(n14641) );
  NAND_GATE U14504 ( .I1(A[11]), .I2(n1401), .O(n14644) );
  NAND_GATE U14505 ( .I1(n14641), .I2(n14644), .O(n14265) );
  NAND_GATE U14506 ( .I1(n14649), .I2(n14265), .O(n14266) );
  INV_GATE U14507 ( .I1(n14644), .O(n14638) );
  NAND_GATE U14508 ( .I1(n14639), .I2(n14638), .O(n14647) );
  NAND_GATE U14509 ( .I1(n14266), .I2(n14647), .O(n14625) );
  INV_GATE U14510 ( .I1(n14625), .O(n14623) );
  NAND_GATE U14511 ( .I1(A[12]), .I2(n1401), .O(n14630) );
  NAND_GATE U14512 ( .I1(n14623), .I2(n14630), .O(n14267) );
  NAND_GATE U14513 ( .I1(n14626), .I2(n14267), .O(n14268) );
  INV_GATE U14514 ( .I1(n14630), .O(n14624) );
  NAND_GATE U14515 ( .I1(n14625), .I2(n14624), .O(n14634) );
  NAND_GATE U14516 ( .I1(n14268), .I2(n14634), .O(n14610) );
  INV_GATE U14517 ( .I1(n14610), .O(n14612) );
  NAND_GATE U14518 ( .I1(A[13]), .I2(n1401), .O(n14615) );
  NAND_GATE U14519 ( .I1(n14612), .I2(n14615), .O(n14269) );
  NAND_GATE U14520 ( .I1(n14620), .I2(n14269), .O(n14270) );
  INV_GATE U14521 ( .I1(n14615), .O(n14609) );
  NAND_GATE U14522 ( .I1(n14610), .I2(n14609), .O(n14618) );
  NAND_GATE U14523 ( .I1(n14270), .I2(n14618), .O(n14596) );
  INV_GATE U14524 ( .I1(n14596), .O(n14594) );
  NAND_GATE U14525 ( .I1(A[14]), .I2(n1401), .O(n14601) );
  NAND_GATE U14526 ( .I1(n14594), .I2(n14601), .O(n14271) );
  NAND_GATE U14527 ( .I1(n14597), .I2(n14271), .O(n14272) );
  INV_GATE U14528 ( .I1(n14601), .O(n14595) );
  NAND_GATE U14529 ( .I1(n14596), .I2(n14595), .O(n14605) );
  NAND_GATE U14530 ( .I1(n14272), .I2(n14605), .O(n14581) );
  INV_GATE U14531 ( .I1(n14581), .O(n14583) );
  NAND_GATE U14532 ( .I1(A[15]), .I2(n1401), .O(n14586) );
  NAND_GATE U14533 ( .I1(n14583), .I2(n14586), .O(n14273) );
  NAND_GATE U14534 ( .I1(n14591), .I2(n14273), .O(n14274) );
  INV_GATE U14535 ( .I1(n14586), .O(n14580) );
  NAND_GATE U14536 ( .I1(n14581), .I2(n14580), .O(n14589) );
  NAND_GATE U14537 ( .I1(n14274), .I2(n14589), .O(n14567) );
  INV_GATE U14538 ( .I1(n14567), .O(n14565) );
  NAND_GATE U14539 ( .I1(A[16]), .I2(n1401), .O(n14572) );
  NAND_GATE U14540 ( .I1(n14565), .I2(n14572), .O(n14275) );
  NAND_GATE U14541 ( .I1(n14568), .I2(n14275), .O(n14276) );
  INV_GATE U14542 ( .I1(n14572), .O(n14566) );
  NAND_GATE U14543 ( .I1(n14567), .I2(n14566), .O(n14576) );
  NAND_GATE U14544 ( .I1(n14276), .I2(n14576), .O(n14552) );
  NAND_GATE U14545 ( .I1(A[17]), .I2(n1401), .O(n14557) );
  NAND_GATE U14546 ( .I1(n14554), .I2(n14557), .O(n14277) );
  NAND_GATE U14547 ( .I1(n14562), .I2(n14277), .O(n14278) );
  INV_GATE U14548 ( .I1(n14557), .O(n14551) );
  NAND_GATE U14549 ( .I1(n14552), .I2(n14551), .O(n14560) );
  NAND_GATE U14550 ( .I1(n14278), .I2(n14560), .O(n14538) );
  INV_GATE U14551 ( .I1(n14538), .O(n14536) );
  NAND_GATE U14552 ( .I1(A[18]), .I2(n1401), .O(n14543) );
  NAND_GATE U14553 ( .I1(n14539), .I2(n14279), .O(n14280) );
  INV_GATE U14554 ( .I1(n14543), .O(n14537) );
  NAND_GATE U14555 ( .I1(n14538), .I2(n14537), .O(n14547) );
  NAND_GATE U14556 ( .I1(n14280), .I2(n14547), .O(n14523) );
  NAND_GATE U14557 ( .I1(A[19]), .I2(n1401), .O(n14528) );
  NAND_GATE U14558 ( .I1(n14525), .I2(n14528), .O(n14281) );
  NAND_GATE U14559 ( .I1(n14533), .I2(n14281), .O(n14282) );
  INV_GATE U14560 ( .I1(n14528), .O(n14522) );
  NAND_GATE U14561 ( .I1(n14523), .I2(n14522), .O(n14531) );
  NAND_GATE U14562 ( .I1(A[20]), .I2(n1401), .O(n14514) );
  NAND_GATE U14563 ( .I1(n791), .I2(n14514), .O(n14283) );
  NAND_GATE U14564 ( .I1(n14510), .I2(n14283), .O(n14284) );
  INV_GATE U14565 ( .I1(n14514), .O(n14508) );
  NAND_GATE U14566 ( .I1(n14509), .I2(n14508), .O(n14518) );
  NAND_GATE U14567 ( .I1(n14284), .I2(n14518), .O(n14496) );
  NAND_GATE U14568 ( .I1(A[21]), .I2(n1401), .O(n14500) );
  NAND_GATE U14569 ( .I1(n14497), .I2(n14500), .O(n14285) );
  NAND_GATE U14570 ( .I1(n14505), .I2(n14285), .O(n14286) );
  INV_GATE U14571 ( .I1(n14500), .O(n14495) );
  NAND_GATE U14572 ( .I1(n14496), .I2(n14495), .O(n14503) );
  NAND_GATE U14573 ( .I1(A[22]), .I2(n1401), .O(n14487) );
  NAND_GATE U14574 ( .I1(n37), .I2(n14286), .O(n14287) );
  NAND_GATE U14575 ( .I1(n14483), .I2(n14287), .O(n14288) );
  INV_GATE U14576 ( .I1(n14487), .O(n14482) );
  NAND_GATE U14577 ( .I1(n14288), .I2(n14491), .O(n14469) );
  INV_GATE U14578 ( .I1(n14469), .O(n14471) );
  NAND_GATE U14579 ( .I1(A[23]), .I2(n1401), .O(n14474) );
  NAND_GATE U14580 ( .I1(n1369), .I2(n14288), .O(n14289) );
  NAND_GATE U14581 ( .I1(n14479), .I2(n14289), .O(n14290) );
  INV_GATE U14582 ( .I1(n14474), .O(n14468) );
  NAND_GATE U14583 ( .I1(n14469), .I2(n14468), .O(n14477) );
  NAND_GATE U14584 ( .I1(n14455), .I2(n440), .O(n14463) );
  OR_GATE U14585 ( .I1(n14291), .I2(n14296), .O(n14294) );
  OR_GATE U14586 ( .I1(n14292), .I2(n14295), .O(n14293) );
  NAND_GATE U14587 ( .I1(n14295), .I2(n1033), .O(n14299) );
  NAND3_GATE U14588 ( .I1(n14299), .I2(n14298), .I3(n14297), .O(n14300) );
  INV_GATE U14589 ( .I1(n14464), .O(n14456) );
  NAND_GATE U14590 ( .I1(n14290), .I2(n439), .O(n14301) );
  NAND_GATE U14591 ( .I1(n14456), .I2(n14301), .O(n14302) );
  NAND_GATE U14592 ( .I1(n14463), .I2(n14302), .O(n14444) );
  INV_GATE U14593 ( .I1(n14303), .O(n14304) );
  NAND_GATE U14594 ( .I1(n14310), .I2(n14304), .O(n14317) );
  NAND_GATE U14595 ( .I1(n14308), .I2(n14307), .O(n14305) );
  NAND_GATE U14596 ( .I1(n14306), .I2(n14305), .O(n14315) );
  NAND_GATE U14597 ( .I1(n14310), .I2(n14309), .O(n14311) );
  NAND_GATE U14598 ( .I1(n14305), .I2(n14311), .O(n14312) );
  NAND_GATE U14599 ( .I1(n14313), .I2(n14312), .O(n14314) );
  NAND_GATE U14600 ( .I1(n14315), .I2(n14314), .O(n14316) );
  NAND_GATE U14601 ( .I1(n14317), .I2(n14316), .O(n14451) );
  NAND_GATE U14602 ( .I1(n14451), .I2(n14318), .O(n14319) );
  NAND_GATE U14603 ( .I1(A[26]), .I2(n1401), .O(n14436) );
  NAND_GATE U14604 ( .I1(n1353), .I2(n14319), .O(n14320) );
  NAND_GATE U14605 ( .I1(n484), .I2(n14320), .O(n14321) );
  NAND_GATE U14606 ( .I1(n1368), .I2(n448), .O(n14440) );
  NAND_GATE U14607 ( .I1(n14326), .I2(n14325), .O(n14323) );
  NAND_GATE U14608 ( .I1(n14324), .I2(n14323), .O(n14331) );
  NAND_GATE U14609 ( .I1(n14331), .I2(n14330), .O(n14332) );
  NAND_GATE U14610 ( .I1(n14333), .I2(n14332), .O(n14429) );
  NAND_GATE U14611 ( .I1(n14321), .I2(n682), .O(n14334) );
  NAND_GATE U14612 ( .I1(n14429), .I2(n14334), .O(n14336) );
  NAND3_GATE U14613 ( .I1(n14416), .I2(n14428), .I3(n14336), .O(n14335) );
  NAND_GATE U14614 ( .I1(n794), .I2(n14335), .O(n14351) );
  INV_GATE U14615 ( .I1(n14416), .O(n14411) );
  NAND_GATE U14616 ( .I1(n14428), .I2(n14336), .O(n14412) );
  NAND_GATE U14617 ( .I1(A[29]), .I2(n1401), .O(n14403) );
  NAND3_GATE U14618 ( .I1(n14351), .I2(n14418), .I3(n14403), .O(n14350) );
  NAND_GATE U14619 ( .I1(n14337), .I2(n14346), .O(n14344) );
  NAND3_GATE U14620 ( .I1(n14339), .I2(n684), .I3(n14338), .O(n14343) );
  NAND_GATE U14621 ( .I1(n14339), .I2(n684), .O(n14340) );
  NAND_GATE U14622 ( .I1(n14341), .I2(n14340), .O(n14342) );
  NAND3_GATE U14623 ( .I1(n14344), .I2(n14343), .I3(n14342), .O(n14349) );
  INV_GATE U14624 ( .I1(n14345), .O(n14347) );
  NAND_GATE U14625 ( .I1(n14347), .I2(n14346), .O(n14348) );
  NAND_GATE U14626 ( .I1(n14349), .I2(n14348), .O(n14408) );
  NAND_GATE U14627 ( .I1(n14350), .I2(n14408), .O(n14352) );
  INV_GATE U14628 ( .I1(n14403), .O(n14398) );
  NAND_GATE U14629 ( .I1(n14418), .I2(n14351), .O(n14399) );
  NAND_GATE U14630 ( .I1(n14398), .I2(n14399), .O(n14406) );
  NAND_GATE U14631 ( .I1(n626), .I2(n633), .O(n14394) );
  NAND_GATE U14632 ( .I1(A[31]), .I2(n1402), .O(n14380) );
  OR_GATE U14633 ( .I1(n14353), .I2(n14362), .O(n14360) );
  OR_GATE U14634 ( .I1(n14361), .I2(n14358), .O(n14359) );
  AND_GATE U14635 ( .I1(n14360), .I2(n14359), .O(n14367) );
  NAND_GATE U14636 ( .I1(n997), .I2(n14361), .O(n14365) );
  NAND3_GATE U14637 ( .I1(n14365), .I2(n14364), .I3(n14363), .O(n14366) );
  NAND_GATE U14638 ( .I1(n14367), .I2(n14366), .O(n14395) );
  NAND_GATE U14639 ( .I1(n14352), .I2(n632), .O(n14368) );
  NAND3_GATE U14640 ( .I1(n14394), .I2(n14380), .I3(n14379), .O(n14828) );
  NAND_GATE U14641 ( .I1(n14827), .I2(n14828), .O(n14382) );
  NAND5_GATE U14642 ( .I1(n14373), .I2(n14372), .I3(n14371), .I4(n14370), .I5(
        n14369), .O(n14374) );
  NAND_GATE U14643 ( .I1(n14375), .I2(n14374), .O(n14376) );
  NAND_GATE U14644 ( .I1(n14382), .I2(n14826), .O(n14377) );
  NAND_GATE U14645 ( .I1(n14378), .I2(n14377), .O(\A1[30] ) );
  AND3_GATE U14646 ( .I1(n14394), .I2(n14380), .I3(n14379), .O(n14831) );
  NAND_GATE U14647 ( .I1(n14830), .I2(n14831), .O(n14381) );
  NAND_GATE U14648 ( .I1(n14382), .I2(n14381), .O(n14385) );
  INV_GATE U14649 ( .I1(n14385), .O(n14383) );
  NAND_GATE U14650 ( .I1(n14384), .I2(n14383), .O(n14388) );
  NAND_GATE U14651 ( .I1(n14386), .I2(n14385), .O(n14387) );
  AND_GATE U14652 ( .I1(n14388), .I2(n14387), .O(\A1[29] ) );
  NAND_GATE U14653 ( .I1(n936), .I2(n14395), .O(n14390) );
  NAND_GATE U14654 ( .I1(n626), .I2(n14390), .O(n14393) );
  NAND_GATE U14655 ( .I1(n14390), .I2(n14389), .O(n14391) );
  OR_GATE U14656 ( .I1(n14395), .I2(n14394), .O(n14396) );
  INV_GATE U14657 ( .I1(n14399), .O(n14400) );
  NAND_GATE U14658 ( .I1(n135), .I2(n14400), .O(n14397) );
  NAND_GATE U14659 ( .I1(n14398), .I2(n14397), .O(n14405) );
  NAND_GATE U14660 ( .I1(n135), .I2(n14399), .O(n14402) );
  NAND_GATE U14661 ( .I1(n14408), .I2(n14400), .O(n14401) );
  NAND3_GATE U14662 ( .I1(n14403), .I2(n14402), .I3(n14401), .O(n14404) );
  NAND_GATE U14663 ( .I1(n14405), .I2(n14404), .O(n14410) );
  INV_GATE U14664 ( .I1(n14406), .O(n14407) );
  NAND_GATE U14665 ( .I1(n14408), .I2(n14407), .O(n14409) );
  NAND_GATE U14666 ( .I1(n14410), .I2(n14409), .O(\A1[27] ) );
  NAND_GATE U14667 ( .I1(n14411), .I2(n14414), .O(n14417) );
  NAND_GATE U14668 ( .I1(n14412), .I2(n794), .O(n14413) );
  NAND_GATE U14669 ( .I1(n14414), .I2(n14413), .O(n14415) );
  OR_GATE U14670 ( .I1(n14419), .I2(n14418), .O(n14420) );
  NAND_GATE U14671 ( .I1(n14422), .I2(n14421), .O(n14427) );
  NAND_GATE U14672 ( .I1(n683), .I2(n128), .O(n14424) );
  NAND3_GATE U14673 ( .I1(n14425), .I2(n14424), .I3(n14423), .O(n14426) );
  NAND_GATE U14674 ( .I1(n14427), .I2(n14426), .O(n14432) );
  INV_GATE U14675 ( .I1(n14428), .O(n14430) );
  NAND_GATE U14676 ( .I1(n14430), .I2(n14429), .O(n14431) );
  NAND_GATE U14677 ( .I1(n14432), .I2(n14431), .O(\A1[25] ) );
  NAND_GATE U14678 ( .I1(n14439), .I2(n1388), .O(n14434) );
  NAND_GATE U14679 ( .I1(n448), .I2(n14434), .O(n14438) );
  NAND_GATE U14680 ( .I1(n484), .I2(n1368), .O(n14433) );
  NAND_GATE U14681 ( .I1(n14434), .I2(n14433), .O(n14435) );
  NAND_GATE U14682 ( .I1(n14436), .I2(n14435), .O(n14437) );
  NAND_GATE U14683 ( .I1(n14438), .I2(n14437), .O(n14442) );
  OR_GATE U14684 ( .I1(n14440), .I2(n14439), .O(n14441) );
  NAND_GATE U14685 ( .I1(n14442), .I2(n14441), .O(\A1[24] ) );
  NAND_GATE U14686 ( .I1(n445), .I2(n560), .O(n14443) );
  NAND_GATE U14687 ( .I1(n529), .I2(n14443), .O(n14449) );
  NAND_GATE U14688 ( .I1(n14444), .I2(n560), .O(n14446) );
  NAND_GATE U14689 ( .I1(n445), .I2(n14451), .O(n14445) );
  NAND3_GATE U14690 ( .I1(n14447), .I2(n14446), .I3(n14445), .O(n14448) );
  NAND_GATE U14691 ( .I1(n14449), .I2(n14448), .O(n14454) );
  INV_GATE U14692 ( .I1(n14450), .O(n14452) );
  NAND_GATE U14693 ( .I1(n14452), .I2(n14451), .O(n14453) );
  NAND_GATE U14694 ( .I1(n14454), .I2(n14453), .O(\A1[23] ) );
  NAND_GATE U14695 ( .I1(n141), .I2(n14464), .O(n14458) );
  NAND_GATE U14696 ( .I1(n14455), .I2(n14458), .O(n14462) );
  NAND_GATE U14697 ( .I1(n440), .I2(n14456), .O(n14457) );
  NAND_GATE U14698 ( .I1(n14458), .I2(n14457), .O(n14459) );
  NAND_GATE U14699 ( .I1(n14460), .I2(n14459), .O(n14461) );
  NAND_GATE U14700 ( .I1(n14462), .I2(n14461), .O(n14466) );
  OR_GATE U14701 ( .I1(n14464), .I2(n14463), .O(n14465) );
  NAND_GATE U14702 ( .I1(n14466), .I2(n14465), .O(\A1[22] ) );
  INV_GATE U14703 ( .I1(n14479), .O(n14470) );
  NAND_GATE U14704 ( .I1(n14470), .I2(n14471), .O(n14467) );
  NAND_GATE U14705 ( .I1(n14468), .I2(n14467), .O(n14476) );
  NAND_GATE U14706 ( .I1(n14470), .I2(n14469), .O(n14473) );
  NAND_GATE U14707 ( .I1(n14479), .I2(n14471), .O(n14472) );
  NAND3_GATE U14708 ( .I1(n14474), .I2(n14473), .I3(n14472), .O(n14475) );
  NAND_GATE U14709 ( .I1(n14476), .I2(n14475), .O(n14481) );
  INV_GATE U14710 ( .I1(n14477), .O(n14478) );
  NAND_GATE U14711 ( .I1(n14479), .I2(n14478), .O(n14480) );
  NAND_GATE U14712 ( .I1(n14481), .I2(n14480), .O(\A1[21] ) );
  NAND_GATE U14713 ( .I1(n14490), .I2(n1270), .O(n14485) );
  NAND_GATE U14714 ( .I1(n14482), .I2(n14485), .O(n14489) );
  NAND_GATE U14715 ( .I1(n14483), .I2(n36), .O(n14484) );
  NAND_GATE U14716 ( .I1(n14485), .I2(n14484), .O(n14486) );
  NAND_GATE U14717 ( .I1(n14487), .I2(n14486), .O(n14488) );
  NAND_GATE U14718 ( .I1(n14489), .I2(n14488), .O(n14493) );
  OR_GATE U14719 ( .I1(n14491), .I2(n14490), .O(n14492) );
  NAND_GATE U14720 ( .I1(n14493), .I2(n14492), .O(\A1[20] ) );
  NAND_GATE U14721 ( .I1(n437), .I2(n14497), .O(n14494) );
  NAND_GATE U14722 ( .I1(n14495), .I2(n14494), .O(n14502) );
  NAND_GATE U14723 ( .I1(n437), .I2(n14496), .O(n14499) );
  NAND_GATE U14724 ( .I1(n14505), .I2(n14497), .O(n14498) );
  NAND3_GATE U14725 ( .I1(n14500), .I2(n14499), .I3(n14498), .O(n14501) );
  NAND_GATE U14726 ( .I1(n14502), .I2(n14501), .O(n14507) );
  INV_GATE U14727 ( .I1(n14503), .O(n14504) );
  NAND_GATE U14728 ( .I1(n14505), .I2(n14504), .O(n14506) );
  NAND_GATE U14729 ( .I1(n14507), .I2(n14506), .O(\A1[19] ) );
  NAND_GATE U14730 ( .I1(n14517), .I2(n791), .O(n14512) );
  NAND_GATE U14731 ( .I1(n14508), .I2(n14512), .O(n14516) );
  NAND_GATE U14732 ( .I1(n14510), .I2(n14509), .O(n14511) );
  NAND_GATE U14733 ( .I1(n14512), .I2(n14511), .O(n14513) );
  NAND_GATE U14734 ( .I1(n14514), .I2(n14513), .O(n14515) );
  NAND_GATE U14735 ( .I1(n14516), .I2(n14515), .O(n14520) );
  OR_GATE U14736 ( .I1(n14518), .I2(n14517), .O(n14519) );
  NAND_GATE U14737 ( .I1(n14520), .I2(n14519), .O(\A1[18] ) );
  INV_GATE U14738 ( .I1(n14533), .O(n14524) );
  NAND_GATE U14739 ( .I1(n14524), .I2(n14525), .O(n14521) );
  NAND_GATE U14740 ( .I1(n14522), .I2(n14521), .O(n14530) );
  NAND_GATE U14741 ( .I1(n14524), .I2(n14523), .O(n14527) );
  NAND_GATE U14742 ( .I1(n14533), .I2(n14525), .O(n14526) );
  NAND3_GATE U14743 ( .I1(n14528), .I2(n14527), .I3(n14526), .O(n14529) );
  NAND_GATE U14744 ( .I1(n14530), .I2(n14529), .O(n14535) );
  INV_GATE U14745 ( .I1(n14531), .O(n14532) );
  NAND_GATE U14746 ( .I1(n14533), .I2(n14532), .O(n14534) );
  NAND_GATE U14747 ( .I1(n14535), .I2(n14534), .O(\A1[17] ) );
  NAND_GATE U14748 ( .I1(n14546), .I2(n14536), .O(n14541) );
  NAND_GATE U14749 ( .I1(n14537), .I2(n14541), .O(n14545) );
  NAND_GATE U14750 ( .I1(n14539), .I2(n14538), .O(n14540) );
  NAND_GATE U14751 ( .I1(n14541), .I2(n14540), .O(n14542) );
  NAND_GATE U14752 ( .I1(n14543), .I2(n14542), .O(n14544) );
  NAND_GATE U14753 ( .I1(n14545), .I2(n14544), .O(n14549) );
  OR_GATE U14754 ( .I1(n14547), .I2(n14546), .O(n14548) );
  NAND_GATE U14755 ( .I1(n14549), .I2(n14548), .O(\A1[16] ) );
  INV_GATE U14756 ( .I1(n14562), .O(n14553) );
  NAND_GATE U14757 ( .I1(n14553), .I2(n14554), .O(n14550) );
  NAND_GATE U14758 ( .I1(n14551), .I2(n14550), .O(n14559) );
  NAND_GATE U14759 ( .I1(n14553), .I2(n14552), .O(n14556) );
  NAND_GATE U14760 ( .I1(n14562), .I2(n14554), .O(n14555) );
  NAND3_GATE U14761 ( .I1(n14557), .I2(n14556), .I3(n14555), .O(n14558) );
  NAND_GATE U14762 ( .I1(n14559), .I2(n14558), .O(n14564) );
  INV_GATE U14763 ( .I1(n14560), .O(n14561) );
  NAND_GATE U14764 ( .I1(n14562), .I2(n14561), .O(n14563) );
  NAND_GATE U14765 ( .I1(n14564), .I2(n14563), .O(\A1[15] ) );
  NAND_GATE U14766 ( .I1(n14575), .I2(n14565), .O(n14570) );
  NAND_GATE U14767 ( .I1(n14566), .I2(n14570), .O(n14574) );
  NAND_GATE U14768 ( .I1(n14568), .I2(n14567), .O(n14569) );
  NAND_GATE U14769 ( .I1(n14570), .I2(n14569), .O(n14571) );
  NAND_GATE U14770 ( .I1(n14572), .I2(n14571), .O(n14573) );
  NAND_GATE U14771 ( .I1(n14574), .I2(n14573), .O(n14578) );
  OR_GATE U14772 ( .I1(n14576), .I2(n14575), .O(n14577) );
  NAND_GATE U14773 ( .I1(n14578), .I2(n14577), .O(\A1[14] ) );
  INV_GATE U14774 ( .I1(n14591), .O(n14582) );
  NAND_GATE U14775 ( .I1(n14582), .I2(n14583), .O(n14579) );
  NAND_GATE U14776 ( .I1(n14580), .I2(n14579), .O(n14588) );
  NAND_GATE U14777 ( .I1(n14582), .I2(n14581), .O(n14585) );
  NAND_GATE U14778 ( .I1(n14591), .I2(n14583), .O(n14584) );
  NAND3_GATE U14779 ( .I1(n14586), .I2(n14585), .I3(n14584), .O(n14587) );
  NAND_GATE U14780 ( .I1(n14588), .I2(n14587), .O(n14593) );
  INV_GATE U14781 ( .I1(n14589), .O(n14590) );
  NAND_GATE U14782 ( .I1(n14591), .I2(n14590), .O(n14592) );
  NAND_GATE U14783 ( .I1(n14593), .I2(n14592), .O(\A1[13] ) );
  NAND_GATE U14784 ( .I1(n14604), .I2(n14594), .O(n14599) );
  NAND_GATE U14785 ( .I1(n14595), .I2(n14599), .O(n14603) );
  NAND_GATE U14786 ( .I1(n14597), .I2(n14596), .O(n14598) );
  NAND_GATE U14787 ( .I1(n14599), .I2(n14598), .O(n14600) );
  NAND_GATE U14788 ( .I1(n14601), .I2(n14600), .O(n14602) );
  NAND_GATE U14789 ( .I1(n14603), .I2(n14602), .O(n14607) );
  OR_GATE U14790 ( .I1(n14605), .I2(n14604), .O(n14606) );
  NAND_GATE U14791 ( .I1(n14607), .I2(n14606), .O(\A1[12] ) );
  INV_GATE U14792 ( .I1(n14620), .O(n14611) );
  NAND_GATE U14793 ( .I1(n14611), .I2(n14612), .O(n14608) );
  NAND_GATE U14794 ( .I1(n14609), .I2(n14608), .O(n14617) );
  NAND_GATE U14795 ( .I1(n14611), .I2(n14610), .O(n14614) );
  NAND_GATE U14796 ( .I1(n14620), .I2(n14612), .O(n14613) );
  NAND3_GATE U14797 ( .I1(n14615), .I2(n14614), .I3(n14613), .O(n14616) );
  NAND_GATE U14798 ( .I1(n14617), .I2(n14616), .O(n14622) );
  INV_GATE U14799 ( .I1(n14618), .O(n14619) );
  NAND_GATE U14800 ( .I1(n14620), .I2(n14619), .O(n14621) );
  NAND_GATE U14801 ( .I1(n14622), .I2(n14621), .O(\A1[11] ) );
  NAND_GATE U14802 ( .I1(n14633), .I2(n14623), .O(n14628) );
  NAND_GATE U14803 ( .I1(n14624), .I2(n14628), .O(n14632) );
  NAND_GATE U14804 ( .I1(n14626), .I2(n14625), .O(n14627) );
  NAND_GATE U14805 ( .I1(n14628), .I2(n14627), .O(n14629) );
  NAND_GATE U14806 ( .I1(n14630), .I2(n14629), .O(n14631) );
  NAND_GATE U14807 ( .I1(n14632), .I2(n14631), .O(n14636) );
  OR_GATE U14808 ( .I1(n14634), .I2(n14633), .O(n14635) );
  NAND_GATE U14809 ( .I1(n14636), .I2(n14635), .O(\A1[10] ) );
  INV_GATE U14810 ( .I1(n14649), .O(n14640) );
  NAND_GATE U14811 ( .I1(n14640), .I2(n14641), .O(n14637) );
  NAND_GATE U14812 ( .I1(n14638), .I2(n14637), .O(n14646) );
  NAND_GATE U14813 ( .I1(n14640), .I2(n14639), .O(n14643) );
  NAND_GATE U14814 ( .I1(n14649), .I2(n14641), .O(n14642) );
  NAND3_GATE U14815 ( .I1(n14644), .I2(n14643), .I3(n14642), .O(n14645) );
  NAND_GATE U14816 ( .I1(n14646), .I2(n14645), .O(n14651) );
  INV_GATE U14817 ( .I1(n14647), .O(n14648) );
  NAND_GATE U14818 ( .I1(n14649), .I2(n14648), .O(n14650) );
  NAND_GATE U14819 ( .I1(n14651), .I2(n14650), .O(\A1[9] ) );
  NAND_GATE U14820 ( .I1(n14662), .I2(n14652), .O(n14657) );
  NAND_GATE U14821 ( .I1(n14653), .I2(n14657), .O(n14661) );
  NAND_GATE U14822 ( .I1(n14655), .I2(n14654), .O(n14656) );
  NAND_GATE U14823 ( .I1(n14657), .I2(n14656), .O(n14658) );
  NAND_GATE U14824 ( .I1(n14659), .I2(n14658), .O(n14660) );
  NAND_GATE U14825 ( .I1(n14661), .I2(n14660), .O(n14665) );
  OR_GATE U14826 ( .I1(n14663), .I2(n14662), .O(n14664) );
  NAND_GATE U14827 ( .I1(n14665), .I2(n14664), .O(\A1[8] ) );
  INV_GATE U14828 ( .I1(n14678), .O(n14669) );
  NAND_GATE U14829 ( .I1(n14669), .I2(n14670), .O(n14666) );
  NAND_GATE U14830 ( .I1(n14667), .I2(n14666), .O(n14675) );
  NAND_GATE U14831 ( .I1(n14669), .I2(n14668), .O(n14672) );
  NAND_GATE U14832 ( .I1(n14678), .I2(n14670), .O(n14671) );
  NAND3_GATE U14833 ( .I1(n14673), .I2(n14672), .I3(n14671), .O(n14674) );
  NAND_GATE U14834 ( .I1(n14675), .I2(n14674), .O(n14680) );
  INV_GATE U14835 ( .I1(n14676), .O(n14677) );
  NAND_GATE U14836 ( .I1(n14678), .I2(n14677), .O(n14679) );
  NAND_GATE U14837 ( .I1(n14680), .I2(n14679), .O(\A1[7] ) );
  NAND_GATE U14838 ( .I1(n14691), .I2(n14681), .O(n14686) );
  NAND_GATE U14839 ( .I1(n14682), .I2(n14686), .O(n14690) );
  NAND_GATE U14840 ( .I1(n14684), .I2(n14683), .O(n14685) );
  NAND_GATE U14841 ( .I1(n14686), .I2(n14685), .O(n14687) );
  NAND_GATE U14842 ( .I1(n14688), .I2(n14687), .O(n14689) );
  NAND_GATE U14843 ( .I1(n14690), .I2(n14689), .O(n14694) );
  OR_GATE U14844 ( .I1(n14692), .I2(n14691), .O(n14693) );
  NAND_GATE U14845 ( .I1(n14694), .I2(n14693), .O(\A1[6] ) );
  INV_GATE U14846 ( .I1(n14707), .O(n14698) );
  NAND_GATE U14847 ( .I1(n14698), .I2(n14699), .O(n14695) );
  NAND_GATE U14848 ( .I1(n14696), .I2(n14695), .O(n14704) );
  NAND_GATE U14849 ( .I1(n14698), .I2(n14697), .O(n14701) );
  NAND_GATE U14850 ( .I1(n14707), .I2(n14699), .O(n14700) );
  NAND3_GATE U14851 ( .I1(n14702), .I2(n14701), .I3(n14700), .O(n14703) );
  NAND_GATE U14852 ( .I1(n14704), .I2(n14703), .O(n14709) );
  INV_GATE U14853 ( .I1(n14705), .O(n14706) );
  NAND_GATE U14854 ( .I1(n14707), .I2(n14706), .O(n14708) );
  NAND_GATE U14855 ( .I1(n14709), .I2(n14708), .O(\A1[5] ) );
  NAND_GATE U14856 ( .I1(n14720), .I2(n14710), .O(n14715) );
  NAND_GATE U14857 ( .I1(n14711), .I2(n14715), .O(n14719) );
  NAND_GATE U14858 ( .I1(n14713), .I2(n14712), .O(n14714) );
  NAND_GATE U14859 ( .I1(n14715), .I2(n14714), .O(n14716) );
  NAND_GATE U14860 ( .I1(n14717), .I2(n14716), .O(n14718) );
  NAND_GATE U14861 ( .I1(n14719), .I2(n14718), .O(n14723) );
  OR_GATE U14862 ( .I1(n14721), .I2(n14720), .O(n14722) );
  NAND_GATE U14863 ( .I1(n14723), .I2(n14722), .O(\A1[4] ) );
  INV_GATE U14864 ( .I1(n14736), .O(n14727) );
  NAND_GATE U14865 ( .I1(n14727), .I2(n14728), .O(n14724) );
  NAND_GATE U14866 ( .I1(n14725), .I2(n14724), .O(n14733) );
  NAND_GATE U14867 ( .I1(n14727), .I2(n14726), .O(n14730) );
  NAND_GATE U14868 ( .I1(n14736), .I2(n14728), .O(n14729) );
  NAND3_GATE U14869 ( .I1(n14731), .I2(n14730), .I3(n14729), .O(n14732) );
  NAND_GATE U14870 ( .I1(n14733), .I2(n14732), .O(n14738) );
  INV_GATE U14871 ( .I1(n14734), .O(n14735) );
  NAND_GATE U14872 ( .I1(n14736), .I2(n14735), .O(n14737) );
  NAND_GATE U14873 ( .I1(n14738), .I2(n14737), .O(\A1[3] ) );
  NAND_GATE U14874 ( .I1(n14749), .I2(n14739), .O(n14744) );
  NAND_GATE U14875 ( .I1(n14740), .I2(n14744), .O(n14748) );
  NAND_GATE U14876 ( .I1(n14742), .I2(n14741), .O(n14743) );
  NAND_GATE U14877 ( .I1(n14744), .I2(n14743), .O(n14745) );
  NAND_GATE U14878 ( .I1(n14746), .I2(n14745), .O(n14747) );
  NAND_GATE U14879 ( .I1(n14748), .I2(n14747), .O(n14752) );
  OR_GATE U14880 ( .I1(n14750), .I2(n14749), .O(n14751) );
  NAND_GATE U14881 ( .I1(n14752), .I2(n14751), .O(\A1[2] ) );
  INV_GATE U14882 ( .I1(n14765), .O(n14756) );
  NAND_GATE U14883 ( .I1(n14756), .I2(n14757), .O(n14753) );
  NAND_GATE U14884 ( .I1(n14754), .I2(n14753), .O(n14762) );
  NAND_GATE U14885 ( .I1(n14756), .I2(n14755), .O(n14759) );
  NAND_GATE U14886 ( .I1(n14765), .I2(n14757), .O(n14758) );
  NAND3_GATE U14887 ( .I1(n14760), .I2(n14759), .I3(n14758), .O(n14761) );
  NAND_GATE U14888 ( .I1(n14762), .I2(n14761), .O(n14767) );
  INV_GATE U14889 ( .I1(n14763), .O(n14764) );
  NAND_GATE U14890 ( .I1(n14765), .I2(n14764), .O(n14766) );
  NAND_GATE U14891 ( .I1(n14767), .I2(n14766), .O(\A1[1] ) );
  NAND_GATE U14892 ( .I1(n14778), .I2(n14768), .O(n14773) );
  NAND_GATE U14893 ( .I1(n14769), .I2(n14773), .O(n14777) );
  NAND_GATE U14894 ( .I1(n14771), .I2(n14770), .O(n14772) );
  NAND_GATE U14895 ( .I1(n14773), .I2(n14772), .O(n14774) );
  NAND_GATE U14896 ( .I1(n14775), .I2(n14774), .O(n14776) );
  NAND_GATE U14897 ( .I1(n14777), .I2(n14776), .O(n14781) );
  OR_GATE U14898 ( .I1(n14779), .I2(n14778), .O(n14780) );
  NAND_GATE U14899 ( .I1(n14781), .I2(n14780), .O(\A1[0] ) );
  AND3_GATE U14900 ( .I1(A[31]), .I2(n346), .I3(n1474), .O(\A2[61] ) );
  INV_GATE U14901 ( .I1(n14782), .O(n14835) );
  INV_GATE U14902 ( .I1(n14783), .O(n14836) );
  AND_GATE U14903 ( .I1(n14785), .I2(n14784), .O(\A2[58] ) );
  AND_GATE U14904 ( .I1(n14787), .I2(n14786), .O(\A2[57] ) );
  AND_GATE U14905 ( .I1(n14789), .I2(n14788), .O(\A2[56] ) );
  AND_GATE U14906 ( .I1(n14791), .I2(n14790), .O(\A2[55] ) );
  AND_GATE U14907 ( .I1(n14793), .I2(n14792), .O(\A2[54] ) );
  AND_GATE U14908 ( .I1(n14795), .I2(n14794), .O(\A2[53] ) );
  AND_GATE U14909 ( .I1(n14797), .I2(n14796), .O(\A2[52] ) );
  AND_GATE U14910 ( .I1(n14799), .I2(n14798), .O(\A2[51] ) );
  AND_GATE U14911 ( .I1(n14801), .I2(n14800), .O(\A2[50] ) );
  AND_GATE U14912 ( .I1(n14803), .I2(n14802), .O(\A2[49] ) );
  AND3_GATE U14913 ( .I1(n14806), .I2(n14805), .I3(n14804), .O(\A2[48] ) );
  AND_GATE U14914 ( .I1(n14808), .I2(n14807), .O(\A2[47] ) );
  AND_GATE U14915 ( .I1(n14810), .I2(n14809), .O(\A2[46] ) );
  AND_GATE U14916 ( .I1(n14812), .I2(n14811), .O(\A2[45] ) );
  AND_GATE U14917 ( .I1(n14815), .I2(n14814), .O(\A2[43] ) );
  AND_GATE U14918 ( .I1(n14817), .I2(n14816), .O(\A2[42] ) );
  AND_GATE U14919 ( .I1(n14818), .I2(n830), .O(\A2[41] ) );
  AND_GATE U14920 ( .I1(n1320), .I2(n14819), .O(\A2[39] ) );
  AND_GATE U14921 ( .I1(n1263), .I2(n1390), .O(\A2[38] ) );
  AND_GATE U14922 ( .I1(n14821), .I2(n14820), .O(\A2[36] ) );
  AND_GATE U14923 ( .I1(n613), .I2(n14822), .O(\A2[34] ) );
  AND3_GATE U14924 ( .I1(n14825), .I2(n14824), .I3(n14823), .O(\A2[32] ) );
  NAND3_GATE U14925 ( .I1(n14828), .I2(n14827), .I3(n14829), .O(n14833) );
  NAND3_GATE U14926 ( .I1(n14831), .I2(n14830), .I3(n14829), .O(n14832) );
  AND3_GATE U14927 ( .I1(n14833), .I2(n14832), .I3(\A1[61] ), .O(n14834) );
  NAND_GATE U14930 ( .I1(B[1]), .I2(A[0]), .O(n14839) );
  AND_GATE U14931 ( .I1(A[0]), .I2(n1401), .O(PRODUCT[0]) );
endmodule


module pps_pf_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_GATE U1 ( .I1(A[2]), .O(SUM[2]) );
  INV_GATE U2 ( .I1(n112), .O(n2) );
  INV_GATE U3 ( .I1(n32), .O(n3) );
  INV_GATE U4 ( .I1(A[3]), .O(n4) );
  INV_GATE U5 ( .I1(A[4]), .O(n5) );
  INV_GATE U6 ( .I1(A[5]), .O(n6) );
  INV_GATE U7 ( .I1(A[6]), .O(n7) );
  INV_GATE U8 ( .I1(A[7]), .O(n8) );
  INV_GATE U9 ( .I1(A[8]), .O(n9) );
  INV_GATE U10 ( .I1(A[11]), .O(n10) );
  INV_GATE U11 ( .I1(A[12]), .O(n11) );
  INV_GATE U12 ( .I1(A[13]), .O(n12) );
  INV_GATE U13 ( .I1(A[14]), .O(n13) );
  INV_GATE U14 ( .I1(A[15]), .O(n14) );
  INV_GATE U15 ( .I1(A[16]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[18]), .O(n17) );
  INV_GATE U18 ( .I1(A[19]), .O(n18) );
  INV_GATE U19 ( .I1(A[20]), .O(n19) );
  INV_GATE U20 ( .I1(A[21]), .O(n20) );
  INV_GATE U21 ( .I1(A[22]), .O(n21) );
  INV_GATE U22 ( .I1(A[23]), .O(n22) );
  INV_GATE U23 ( .I1(A[24]), .O(n23) );
  INV_GATE U24 ( .I1(A[25]), .O(n24) );
  INV_GATE U25 ( .I1(A[26]), .O(n25) );
  INV_GATE U26 ( .I1(A[27]), .O(n26) );
  INV_GATE U27 ( .I1(A[28]), .O(n27) );
  INV_GATE U28 ( .I1(A[29]), .O(n28) );
  INV_GATE U29 ( .I1(A[30]), .O(n29) );
  NAND_GATE U30 ( .I1(n30), .I2(n31), .O(SUM[9]) );
  NAND_GATE U31 ( .I1(A[9]), .I2(n3), .O(n31) );
  OR_GATE U32 ( .I1(n3), .I2(A[9]), .O(n30) );
  NAND_GATE U33 ( .I1(n33), .I2(n34), .O(SUM[8]) );
  OR_GATE U34 ( .I1(n9), .I2(n35), .O(n34) );
  NAND_GATE U35 ( .I1(n35), .I2(n9), .O(n33) );
  AND_GATE U36 ( .I1(A[7]), .I2(n36), .O(n35) );
  NAND_GATE U37 ( .I1(n37), .I2(n38), .O(SUM[7]) );
  OR_GATE U38 ( .I1(n8), .I2(n36), .O(n38) );
  NAND_GATE U39 ( .I1(n36), .I2(n8), .O(n37) );
  NAND_GATE U40 ( .I1(n39), .I2(n40), .O(SUM[6]) );
  OR_GATE U41 ( .I1(n7), .I2(n41), .O(n40) );
  NAND_GATE U42 ( .I1(n41), .I2(n7), .O(n39) );
  AND_GATE U43 ( .I1(A[5]), .I2(n42), .O(n41) );
  NAND_GATE U44 ( .I1(n43), .I2(n44), .O(SUM[5]) );
  OR_GATE U45 ( .I1(n6), .I2(n42), .O(n44) );
  NAND_GATE U46 ( .I1(n42), .I2(n6), .O(n43) );
  NAND_GATE U47 ( .I1(n45), .I2(n46), .O(SUM[4]) );
  OR_GATE U48 ( .I1(n5), .I2(n47), .O(n46) );
  NAND_GATE U49 ( .I1(n47), .I2(n5), .O(n45) );
  AND_GATE U50 ( .I1(A[3]), .I2(A[2]), .O(n47) );
  NAND_GATE U51 ( .I1(n48), .I2(n49), .O(SUM[3]) );
  NAND_GATE U52 ( .I1(A[3]), .I2(SUM[2]), .O(n49) );
  NAND_GATE U53 ( .I1(A[2]), .I2(n4), .O(n48) );
  NAND_GATE U54 ( .I1(n50), .I2(n51), .O(SUM[31]) );
  NAND_GATE U55 ( .I1(A[31]), .I2(n52), .O(n51) );
  OR_GATE U56 ( .I1(n52), .I2(A[31]), .O(n50) );
  NAND_GATE U57 ( .I1(A[30]), .I2(n53), .O(n52) );
  NAND_GATE U58 ( .I1(n54), .I2(n55), .O(SUM[30]) );
  OR_GATE U59 ( .I1(n29), .I2(n53), .O(n55) );
  NAND_GATE U60 ( .I1(n53), .I2(n29), .O(n54) );
  AND_GATE U61 ( .I1(A[29]), .I2(n56), .O(n53) );
  NAND_GATE U62 ( .I1(n57), .I2(n58), .O(SUM[29]) );
  OR_GATE U63 ( .I1(n28), .I2(n56), .O(n58) );
  NAND_GATE U64 ( .I1(n56), .I2(n28), .O(n57) );
  AND3_GATE U65 ( .I1(A[27]), .I2(n59), .I3(A[28]), .O(n56) );
  NAND_GATE U66 ( .I1(n60), .I2(n61), .O(SUM[28]) );
  OR_GATE U67 ( .I1(n27), .I2(n62), .O(n61) );
  NAND_GATE U68 ( .I1(n62), .I2(n27), .O(n60) );
  AND_GATE U69 ( .I1(A[27]), .I2(n59), .O(n62) );
  NAND_GATE U70 ( .I1(n63), .I2(n64), .O(SUM[27]) );
  OR_GATE U71 ( .I1(n26), .I2(n59), .O(n64) );
  NAND_GATE U72 ( .I1(n59), .I2(n26), .O(n63) );
  AND3_GATE U73 ( .I1(A[25]), .I2(n65), .I3(A[26]), .O(n59) );
  NAND_GATE U74 ( .I1(n66), .I2(n67), .O(SUM[26]) );
  OR_GATE U75 ( .I1(n25), .I2(n68), .O(n67) );
  NAND_GATE U76 ( .I1(n68), .I2(n25), .O(n66) );
  AND_GATE U77 ( .I1(A[25]), .I2(n65), .O(n68) );
  NAND_GATE U78 ( .I1(n69), .I2(n70), .O(SUM[25]) );
  OR_GATE U79 ( .I1(n24), .I2(n65), .O(n70) );
  NAND_GATE U80 ( .I1(n65), .I2(n24), .O(n69) );
  AND3_GATE U81 ( .I1(A[23]), .I2(n71), .I3(A[24]), .O(n65) );
  NAND_GATE U82 ( .I1(n72), .I2(n73), .O(SUM[24]) );
  OR_GATE U83 ( .I1(n23), .I2(n74), .O(n73) );
  NAND_GATE U84 ( .I1(n74), .I2(n23), .O(n72) );
  AND_GATE U85 ( .I1(A[23]), .I2(n71), .O(n74) );
  NAND_GATE U86 ( .I1(n75), .I2(n76), .O(SUM[23]) );
  OR_GATE U87 ( .I1(n22), .I2(n71), .O(n76) );
  NAND_GATE U88 ( .I1(n71), .I2(n22), .O(n75) );
  AND3_GATE U89 ( .I1(A[21]), .I2(n77), .I3(A[22]), .O(n71) );
  NAND_GATE U90 ( .I1(n78), .I2(n79), .O(SUM[22]) );
  OR_GATE U91 ( .I1(n21), .I2(n80), .O(n79) );
  NAND_GATE U92 ( .I1(n80), .I2(n21), .O(n78) );
  AND_GATE U93 ( .I1(A[21]), .I2(n77), .O(n80) );
  NAND_GATE U94 ( .I1(n81), .I2(n82), .O(SUM[21]) );
  OR_GATE U95 ( .I1(n20), .I2(n77), .O(n82) );
  NAND_GATE U96 ( .I1(n77), .I2(n20), .O(n81) );
  AND3_GATE U97 ( .I1(A[19]), .I2(n83), .I3(A[20]), .O(n77) );
  NAND_GATE U98 ( .I1(n84), .I2(n85), .O(SUM[20]) );
  OR_GATE U99 ( .I1(n19), .I2(n86), .O(n85) );
  NAND_GATE U100 ( .I1(n86), .I2(n19), .O(n84) );
  AND_GATE U101 ( .I1(A[19]), .I2(n83), .O(n86) );
  NAND_GATE U102 ( .I1(n87), .I2(n88), .O(SUM[19]) );
  OR_GATE U103 ( .I1(n18), .I2(n83), .O(n88) );
  NAND_GATE U104 ( .I1(n83), .I2(n18), .O(n87) );
  AND3_GATE U105 ( .I1(A[17]), .I2(n89), .I3(A[18]), .O(n83) );
  NAND_GATE U106 ( .I1(n90), .I2(n91), .O(SUM[18]) );
  OR_GATE U107 ( .I1(n17), .I2(n92), .O(n91) );
  NAND_GATE U108 ( .I1(n92), .I2(n17), .O(n90) );
  AND_GATE U109 ( .I1(A[17]), .I2(n89), .O(n92) );
  NAND_GATE U110 ( .I1(n93), .I2(n94), .O(SUM[17]) );
  OR_GATE U111 ( .I1(n16), .I2(n89), .O(n94) );
  NAND_GATE U112 ( .I1(n89), .I2(n16), .O(n93) );
  AND3_GATE U113 ( .I1(A[15]), .I2(n95), .I3(A[16]), .O(n89) );
  NAND_GATE U114 ( .I1(n96), .I2(n97), .O(SUM[16]) );
  OR_GATE U115 ( .I1(n15), .I2(n98), .O(n97) );
  NAND_GATE U116 ( .I1(n98), .I2(n15), .O(n96) );
  AND_GATE U117 ( .I1(A[15]), .I2(n95), .O(n98) );
  NAND_GATE U118 ( .I1(n99), .I2(n100), .O(SUM[15]) );
  OR_GATE U119 ( .I1(n14), .I2(n95), .O(n100) );
  NAND_GATE U120 ( .I1(n95), .I2(n14), .O(n99) );
  AND3_GATE U121 ( .I1(A[13]), .I2(n101), .I3(A[14]), .O(n95) );
  NAND_GATE U122 ( .I1(n102), .I2(n103), .O(SUM[14]) );
  OR_GATE U123 ( .I1(n13), .I2(n104), .O(n103) );
  NAND_GATE U124 ( .I1(n104), .I2(n13), .O(n102) );
  AND_GATE U125 ( .I1(A[13]), .I2(n101), .O(n104) );
  NAND_GATE U126 ( .I1(n105), .I2(n106), .O(SUM[13]) );
  OR_GATE U127 ( .I1(n12), .I2(n101), .O(n106) );
  NAND_GATE U128 ( .I1(n101), .I2(n12), .O(n105) );
  AND3_GATE U129 ( .I1(A[11]), .I2(n2), .I3(A[12]), .O(n101) );
  NAND_GATE U130 ( .I1(n107), .I2(n108), .O(SUM[12]) );
  OR_GATE U131 ( .I1(n11), .I2(n109), .O(n108) );
  NAND_GATE U132 ( .I1(n109), .I2(n11), .O(n107) );
  AND_GATE U133 ( .I1(A[11]), .I2(n2), .O(n109) );
  NAND_GATE U134 ( .I1(n110), .I2(n111), .O(SUM[11]) );
  NAND_GATE U135 ( .I1(A[11]), .I2(n112), .O(n111) );
  NAND_GATE U136 ( .I1(n2), .I2(n10), .O(n110) );
  NAND3_GATE U137 ( .I1(n32), .I2(A[9]), .I3(A[10]), .O(n112) );
  NAND_GATE U138 ( .I1(n113), .I2(n114), .O(SUM[10]) );
  NAND_GATE U139 ( .I1(A[10]), .I2(n115), .O(n114) );
  OR_GATE U140 ( .I1(n115), .I2(A[10]), .O(n113) );
  NAND_GATE U141 ( .I1(n32), .I2(A[9]), .O(n115) );
  AND3_GATE U142 ( .I1(A[7]), .I2(n36), .I3(A[8]), .O(n32) );
  AND3_GATE U143 ( .I1(A[5]), .I2(n42), .I3(A[6]), .O(n36) );
  AND3_GATE U144 ( .I1(A[3]), .I2(A[2]), .I3(A[4]), .O(n42) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398;

  AND_GATE U1 ( .I1(n161), .I2(n160), .O(n1) );
  NAND_GATE U2 ( .I1(n163), .I2(n4), .O(n2) );
  AND_GATE U3 ( .I1(n2), .I2(n3), .O(n158) );
  OR_GATE U4 ( .I1(n160), .I2(n161), .O(n3) );
  AND_GATE U5 ( .I1(B[30]), .I2(n5), .O(n4) );
  INV_GATE U6 ( .I1(n160), .O(n5) );
  AND_GATE U7 ( .I1(n266), .I2(n92), .O(n6) );
  NAND_GATE U8 ( .I1(n268), .I2(n9), .O(n7) );
  AND_GATE U9 ( .I1(n7), .I2(n8), .O(n257) );
  OR_GATE U10 ( .I1(n92), .I2(n266), .O(n8) );
  AND_GATE U11 ( .I1(B[19]), .I2(A[20]), .O(n9) );
  AND_GATE U12 ( .I1(n267), .I2(n12), .O(n10) );
  OR_GATE U13 ( .I1(n10), .I2(n11), .O(n13) );
  AND_GATE U14 ( .I1(n93), .I2(n92), .O(n11) );
  AND_GATE U15 ( .I1(n266), .I2(n93), .O(n12) );
  NAND_GATE U16 ( .I1(n259), .I2(n16), .O(n14) );
  AND_GATE U17 ( .I1(n14), .I2(n15), .O(n248) );
  OR_GATE U18 ( .I1(n93), .I2(n257), .O(n15) );
  AND_GATE U19 ( .I1(B[20]), .I2(A[21]), .O(n16) );
  AND_GATE U20 ( .I1(n248), .I2(n94), .O(n17) );
  NAND_GATE U21 ( .I1(n250), .I2(n20), .O(n18) );
  AND_GATE U22 ( .I1(n18), .I2(n19), .O(n239) );
  OR_GATE U23 ( .I1(n94), .I2(n248), .O(n19) );
  AND_GATE U24 ( .I1(B[21]), .I2(A[22]), .O(n20) );
  AND_GATE U25 ( .I1(n249), .I2(n23), .O(n21) );
  OR_GATE U26 ( .I1(n21), .I2(n22), .O(n24) );
  AND_GATE U27 ( .I1(n95), .I2(n94), .O(n22) );
  AND_GATE U28 ( .I1(n248), .I2(n95), .O(n23) );
  NAND_GATE U29 ( .I1(n241), .I2(n27), .O(n25) );
  AND_GATE U30 ( .I1(n25), .I2(n26), .O(n230) );
  OR_GATE U31 ( .I1(n95), .I2(n239), .O(n26) );
  AND_GATE U32 ( .I1(B[22]), .I2(A[23]), .O(n27) );
  AND_GATE U33 ( .I1(n230), .I2(n96), .O(n28) );
  NAND_GATE U34 ( .I1(n232), .I2(n31), .O(n29) );
  AND_GATE U35 ( .I1(n29), .I2(n30), .O(n221) );
  OR_GATE U36 ( .I1(n96), .I2(n230), .O(n30) );
  AND_GATE U37 ( .I1(B[23]), .I2(A[24]), .O(n31) );
  AND_GATE U38 ( .I1(n231), .I2(n34), .O(n32) );
  OR_GATE U39 ( .I1(n32), .I2(n33), .O(n35) );
  AND_GATE U40 ( .I1(n97), .I2(n96), .O(n33) );
  AND_GATE U41 ( .I1(n230), .I2(n97), .O(n34) );
  NAND_GATE U42 ( .I1(n223), .I2(n38), .O(n36) );
  AND_GATE U43 ( .I1(n36), .I2(n37), .O(n212) );
  OR_GATE U44 ( .I1(n97), .I2(n221), .O(n37) );
  AND_GATE U45 ( .I1(B[24]), .I2(A[25]), .O(n38) );
  AND_GATE U46 ( .I1(n213), .I2(n41), .O(n39) );
  OR_GATE U47 ( .I1(n39), .I2(n40), .O(n52) );
  AND_GATE U48 ( .I1(n49), .I2(n50), .O(n40) );
  AND_GATE U49 ( .I1(n212), .I2(n49), .O(n41) );
  AND_GATE U50 ( .I1(n212), .I2(n98), .O(n42) );
  NAND_GATE U51 ( .I1(n214), .I2(n45), .O(n43) );
  AND_GATE U52 ( .I1(n43), .I2(n44), .O(n203) );
  OR_GATE U53 ( .I1(n98), .I2(n212), .O(n44) );
  AND_GATE U54 ( .I1(B[25]), .I2(A[26]), .O(n45) );
  AND_GATE U55 ( .I1(n213), .I2(n48), .O(n46) );
  OR_GATE U56 ( .I1(n46), .I2(n47), .O(n55) );
  AND_GATE U57 ( .I1(n99), .I2(n98), .O(n47) );
  AND_GATE U58 ( .I1(n212), .I2(n99), .O(n48) );
  OR_GATE U59 ( .I1(n59), .I2(n100), .O(n49) );
  OR_GATE U60 ( .I1(n98), .I2(n59), .O(n50) );
  NAND_GATE U61 ( .I1(n205), .I2(n53), .O(n51) );
  AND_GATE U62 ( .I1(n51), .I2(n52), .O(n60) );
  AND_GATE U63 ( .I1(B[26]), .I2(n54), .O(n53) );
  INV_GATE U64 ( .I1(n59), .O(n54) );
  NAND_GATE U65 ( .I1(n205), .I2(n58), .O(n56) );
  AND_GATE U66 ( .I1(n56), .I2(n57), .O(n194) );
  OR_GATE U67 ( .I1(n99), .I2(n203), .O(n57) );
  AND_GATE U68 ( .I1(B[26]), .I2(A[27]), .O(n58) );
  AND_GATE U69 ( .I1(n100), .I2(n99), .O(n59) );
  NAND_GATE U70 ( .I1(n196), .I2(n63), .O(n61) );
  AND_GATE U71 ( .I1(n61), .I2(n62), .O(n185) );
  OR_GATE U72 ( .I1(n100), .I2(n194), .O(n62) );
  AND_GATE U73 ( .I1(B[27]), .I2(A[28]), .O(n63) );
  OR_GATE U74 ( .I1(n101), .I2(n102), .O(n64) );
  AND_GATE U75 ( .I1(n185), .I2(n101), .O(n65) );
  AND_GATE U76 ( .I1(n186), .I2(n68), .O(n66) );
  OR_GATE U77 ( .I1(n66), .I2(n67), .O(n72) );
  AND_GATE U78 ( .I1(n102), .I2(n101), .O(n67) );
  AND_GATE U79 ( .I1(n185), .I2(n102), .O(n68) );
  NAND_GATE U80 ( .I1(n172), .I2(n71), .O(n69) );
  AND_GATE U81 ( .I1(n69), .I2(n70), .O(n161) );
  OR_GATE U82 ( .I1(n173), .I2(n64), .O(n70) );
  AND_GATE U83 ( .I1(B[29]), .I2(A[30]), .O(n71) );
  INV_GATE U84 ( .I1(A[1]), .O(n73) );
  INV_GATE U85 ( .I1(A[2]), .O(n74) );
  INV_GATE U86 ( .I1(A[3]), .O(n75) );
  INV_GATE U87 ( .I1(A[4]), .O(n76) );
  INV_GATE U88 ( .I1(A[5]), .O(n77) );
  INV_GATE U89 ( .I1(A[6]), .O(n78) );
  INV_GATE U90 ( .I1(A[7]), .O(n79) );
  INV_GATE U91 ( .I1(A[8]), .O(n80) );
  INV_GATE U92 ( .I1(A[9]), .O(n81) );
  INV_GATE U93 ( .I1(A[10]), .O(n82) );
  INV_GATE U94 ( .I1(A[11]), .O(n83) );
  INV_GATE U95 ( .I1(A[12]), .O(n84) );
  INV_GATE U96 ( .I1(A[13]), .O(n85) );
  INV_GATE U97 ( .I1(A[14]), .O(n86) );
  INV_GATE U98 ( .I1(A[15]), .O(n87) );
  INV_GATE U99 ( .I1(A[16]), .O(n88) );
  INV_GATE U100 ( .I1(A[17]), .O(n89) );
  INV_GATE U101 ( .I1(A[18]), .O(n90) );
  INV_GATE U102 ( .I1(A[19]), .O(n91) );
  INV_GATE U103 ( .I1(A[20]), .O(n92) );
  INV_GATE U104 ( .I1(A[21]), .O(n93) );
  INV_GATE U105 ( .I1(A[22]), .O(n94) );
  INV_GATE U106 ( .I1(A[23]), .O(n95) );
  INV_GATE U107 ( .I1(A[24]), .O(n96) );
  INV_GATE U108 ( .I1(A[25]), .O(n97) );
  INV_GATE U109 ( .I1(A[26]), .O(n98) );
  INV_GATE U110 ( .I1(A[27]), .O(n99) );
  INV_GATE U111 ( .I1(A[28]), .O(n100) );
  INV_GATE U112 ( .I1(A[29]), .O(n101) );
  INV_GATE U113 ( .I1(A[30]), .O(n102) );
  INV_GATE U114 ( .I1(A[31]), .O(n103) );
  INV_GATE U115 ( .I1(A[32]), .O(n104) );
  INV_GATE U116 ( .I1(B[0]), .O(n105) );
  AND_GATE U117 ( .I1(n106), .I2(n107), .O(SUM[9]) );
  NAND_GATE U118 ( .I1(n108), .I2(n109), .O(n107) );
  OR_GATE U119 ( .I1(n108), .I2(n109), .O(n106) );
  AND_GATE U120 ( .I1(n110), .I2(n111), .O(n108) );
  NAND_GATE U121 ( .I1(B[9]), .I2(n81), .O(n111) );
  OR_GATE U122 ( .I1(n81), .I2(B[9]), .O(n110) );
  AND_GATE U123 ( .I1(n112), .I2(n113), .O(SUM[8]) );
  NAND_GATE U124 ( .I1(n114), .I2(n115), .O(n113) );
  OR_GATE U125 ( .I1(n114), .I2(n115), .O(n112) );
  AND_GATE U126 ( .I1(n116), .I2(n117), .O(n114) );
  NAND_GATE U127 ( .I1(B[8]), .I2(n80), .O(n117) );
  OR_GATE U128 ( .I1(n80), .I2(B[8]), .O(n116) );
  AND_GATE U129 ( .I1(n118), .I2(n119), .O(SUM[7]) );
  NAND_GATE U130 ( .I1(n120), .I2(n121), .O(n119) );
  OR_GATE U131 ( .I1(n120), .I2(n121), .O(n118) );
  AND_GATE U132 ( .I1(n122), .I2(n123), .O(n120) );
  NAND_GATE U133 ( .I1(B[7]), .I2(n79), .O(n123) );
  OR_GATE U134 ( .I1(n79), .I2(B[7]), .O(n122) );
  AND_GATE U135 ( .I1(n124), .I2(n125), .O(SUM[6]) );
  NAND_GATE U136 ( .I1(n126), .I2(n127), .O(n125) );
  OR_GATE U137 ( .I1(n126), .I2(n127), .O(n124) );
  AND_GATE U138 ( .I1(n128), .I2(n129), .O(n126) );
  NAND_GATE U139 ( .I1(B[6]), .I2(n78), .O(n129) );
  OR_GATE U140 ( .I1(n78), .I2(B[6]), .O(n128) );
  AND_GATE U141 ( .I1(n130), .I2(n131), .O(SUM[5]) );
  NAND_GATE U142 ( .I1(n132), .I2(n133), .O(n131) );
  OR_GATE U143 ( .I1(n132), .I2(n133), .O(n130) );
  AND_GATE U144 ( .I1(n134), .I2(n135), .O(n132) );
  NAND_GATE U145 ( .I1(B[5]), .I2(n77), .O(n135) );
  OR_GATE U146 ( .I1(n77), .I2(B[5]), .O(n134) );
  AND_GATE U147 ( .I1(n136), .I2(n137), .O(SUM[4]) );
  NAND_GATE U148 ( .I1(n138), .I2(n139), .O(n137) );
  OR_GATE U149 ( .I1(n138), .I2(n139), .O(n136) );
  AND_GATE U150 ( .I1(n140), .I2(n141), .O(n138) );
  NAND_GATE U151 ( .I1(B[4]), .I2(n76), .O(n141) );
  OR_GATE U152 ( .I1(n76), .I2(B[4]), .O(n140) );
  AND_GATE U153 ( .I1(n142), .I2(n143), .O(SUM[3]) );
  NAND_GATE U154 ( .I1(n144), .I2(n145), .O(n143) );
  OR_GATE U155 ( .I1(n144), .I2(n145), .O(n142) );
  AND_GATE U156 ( .I1(n146), .I2(n147), .O(n144) );
  NAND_GATE U157 ( .I1(B[3]), .I2(n75), .O(n147) );
  OR_GATE U158 ( .I1(n75), .I2(B[3]), .O(n146) );
  AND_GATE U159 ( .I1(n148), .I2(n149), .O(SUM[32]) );
  NAND_GATE U160 ( .I1(n150), .I2(n151), .O(n149) );
  OR_GATE U161 ( .I1(n151), .I2(n150), .O(n148) );
  AND_GATE U162 ( .I1(n152), .I2(n153), .O(n150) );
  NAND_GATE U163 ( .I1(B[31]), .I2(n154), .O(n153) );
  NAND_GATE U164 ( .I1(n155), .I2(n103), .O(n154) );
  OR_GATE U165 ( .I1(n103), .I2(n155), .O(n152) );
  AND_GATE U166 ( .I1(n156), .I2(n157), .O(n151) );
  NAND_GATE U167 ( .I1(B[32]), .I2(n104), .O(n157) );
  OR_GATE U168 ( .I1(n104), .I2(B[32]), .O(n156) );
  AND_GATE U169 ( .I1(n158), .I2(n159), .O(SUM[31]) );
  NAND_GATE U170 ( .I1(n162), .I2(n1), .O(n159) );
  AND_GATE U171 ( .I1(n161), .I2(n162), .O(n155) );
  NAND_GATE U172 ( .I1(B[30]), .I2(n163), .O(n162) );
  NAND_GATE U173 ( .I1(n72), .I2(n171), .O(n163) );
  AND_GATE U174 ( .I1(n165), .I2(n166), .O(n160) );
  NAND_GATE U175 ( .I1(B[31]), .I2(n103), .O(n166) );
  OR_GATE U176 ( .I1(n103), .I2(B[31]), .O(n165) );
  AND_GATE U177 ( .I1(n167), .I2(n168), .O(SUM[30]) );
  NAND_GATE U178 ( .I1(n169), .I2(n164), .O(n168) );
  OR_GATE U179 ( .I1(n169), .I2(n164), .O(n167) );
  AND_GATE U180 ( .I1(n170), .I2(n171), .O(n164) );
  NAND_GATE U181 ( .I1(B[29]), .I2(n172), .O(n171) );
  NAND_GATE U182 ( .I1(n65), .I2(n186), .O(n172) );
  OR_GATE U183 ( .I1(n101), .I2(n173), .O(n170) );
  AND_GATE U184 ( .I1(n174), .I2(n175), .O(n169) );
  NAND_GATE U185 ( .I1(B[30]), .I2(n102), .O(n175) );
  OR_GATE U186 ( .I1(n102), .I2(B[30]), .O(n174) );
  AND_GATE U187 ( .I1(n176), .I2(n177), .O(SUM[2]) );
  NAND_GATE U188 ( .I1(n178), .I2(n179), .O(n177) );
  OR_GATE U189 ( .I1(n178), .I2(n179), .O(n176) );
  AND_GATE U190 ( .I1(n180), .I2(n181), .O(n178) );
  NAND_GATE U191 ( .I1(B[2]), .I2(n74), .O(n181) );
  OR_GATE U192 ( .I1(n74), .I2(B[2]), .O(n180) );
  AND_GATE U193 ( .I1(n182), .I2(n183), .O(SUM[29]) );
  NAND_GATE U194 ( .I1(n184), .I2(n173), .O(n183) );
  OR_GATE U195 ( .I1(n184), .I2(n173), .O(n182) );
  AND_GATE U196 ( .I1(n185), .I2(n186), .O(n173) );
  NAND_GATE U197 ( .I1(B[28]), .I2(n187), .O(n186) );
  NAND_GATE U198 ( .I1(n60), .I2(n195), .O(n187) );
  AND_GATE U199 ( .I1(n189), .I2(n190), .O(n184) );
  NAND_GATE U200 ( .I1(B[29]), .I2(n101), .O(n190) );
  OR_GATE U201 ( .I1(n101), .I2(B[29]), .O(n189) );
  AND_GATE U202 ( .I1(n191), .I2(n192), .O(SUM[28]) );
  NAND_GATE U203 ( .I1(n193), .I2(n188), .O(n192) );
  OR_GATE U204 ( .I1(n193), .I2(n188), .O(n191) );
  AND_GATE U205 ( .I1(n194), .I2(n195), .O(n188) );
  NAND_GATE U206 ( .I1(B[27]), .I2(n196), .O(n195) );
  NAND_GATE U207 ( .I1(n55), .I2(n204), .O(n196) );
  AND_GATE U208 ( .I1(n198), .I2(n199), .O(n193) );
  NAND_GATE U209 ( .I1(B[28]), .I2(n100), .O(n199) );
  OR_GATE U210 ( .I1(n100), .I2(B[28]), .O(n198) );
  AND_GATE U211 ( .I1(n200), .I2(n201), .O(SUM[27]) );
  NAND_GATE U212 ( .I1(n202), .I2(n197), .O(n201) );
  OR_GATE U213 ( .I1(n202), .I2(n197), .O(n200) );
  AND_GATE U214 ( .I1(n203), .I2(n204), .O(n197) );
  NAND_GATE U215 ( .I1(B[26]), .I2(n205), .O(n204) );
  NAND_GATE U216 ( .I1(n42), .I2(n213), .O(n205) );
  AND_GATE U217 ( .I1(n207), .I2(n208), .O(n202) );
  NAND_GATE U218 ( .I1(B[27]), .I2(n99), .O(n208) );
  OR_GATE U219 ( .I1(n99), .I2(B[27]), .O(n207) );
  AND_GATE U220 ( .I1(n209), .I2(n210), .O(SUM[26]) );
  NAND_GATE U221 ( .I1(n211), .I2(n206), .O(n210) );
  OR_GATE U222 ( .I1(n211), .I2(n206), .O(n209) );
  AND_GATE U223 ( .I1(n212), .I2(n213), .O(n206) );
  NAND_GATE U224 ( .I1(B[25]), .I2(n214), .O(n213) );
  NAND_GATE U225 ( .I1(n35), .I2(n222), .O(n214) );
  AND_GATE U226 ( .I1(n216), .I2(n217), .O(n211) );
  NAND_GATE U227 ( .I1(B[26]), .I2(n98), .O(n217) );
  OR_GATE U228 ( .I1(n98), .I2(B[26]), .O(n216) );
  AND_GATE U229 ( .I1(n218), .I2(n219), .O(SUM[25]) );
  NAND_GATE U230 ( .I1(n220), .I2(n215), .O(n219) );
  OR_GATE U231 ( .I1(n220), .I2(n215), .O(n218) );
  AND_GATE U232 ( .I1(n221), .I2(n222), .O(n215) );
  NAND_GATE U233 ( .I1(B[24]), .I2(n223), .O(n222) );
  NAND_GATE U234 ( .I1(n28), .I2(n231), .O(n223) );
  AND_GATE U235 ( .I1(n225), .I2(n226), .O(n220) );
  NAND_GATE U236 ( .I1(B[25]), .I2(n97), .O(n226) );
  OR_GATE U237 ( .I1(n97), .I2(B[25]), .O(n225) );
  AND_GATE U238 ( .I1(n227), .I2(n228), .O(SUM[24]) );
  NAND_GATE U239 ( .I1(n229), .I2(n224), .O(n228) );
  OR_GATE U240 ( .I1(n229), .I2(n224), .O(n227) );
  AND_GATE U241 ( .I1(n230), .I2(n231), .O(n224) );
  NAND_GATE U242 ( .I1(B[23]), .I2(n232), .O(n231) );
  NAND_GATE U243 ( .I1(n24), .I2(n240), .O(n232) );
  AND_GATE U244 ( .I1(n234), .I2(n235), .O(n229) );
  NAND_GATE U245 ( .I1(B[24]), .I2(n96), .O(n235) );
  OR_GATE U246 ( .I1(n96), .I2(B[24]), .O(n234) );
  AND_GATE U247 ( .I1(n236), .I2(n237), .O(SUM[23]) );
  NAND_GATE U248 ( .I1(n238), .I2(n233), .O(n237) );
  OR_GATE U249 ( .I1(n238), .I2(n233), .O(n236) );
  AND_GATE U250 ( .I1(n239), .I2(n240), .O(n233) );
  NAND_GATE U251 ( .I1(B[22]), .I2(n241), .O(n240) );
  NAND_GATE U252 ( .I1(n17), .I2(n249), .O(n241) );
  AND_GATE U253 ( .I1(n243), .I2(n244), .O(n238) );
  NAND_GATE U254 ( .I1(B[23]), .I2(n95), .O(n244) );
  OR_GATE U255 ( .I1(n95), .I2(B[23]), .O(n243) );
  AND_GATE U256 ( .I1(n245), .I2(n246), .O(SUM[22]) );
  NAND_GATE U257 ( .I1(n247), .I2(n242), .O(n246) );
  OR_GATE U258 ( .I1(n247), .I2(n242), .O(n245) );
  AND_GATE U259 ( .I1(n248), .I2(n249), .O(n242) );
  NAND_GATE U260 ( .I1(B[21]), .I2(n250), .O(n249) );
  NAND_GATE U261 ( .I1(n13), .I2(n258), .O(n250) );
  AND_GATE U262 ( .I1(n252), .I2(n253), .O(n247) );
  NAND_GATE U263 ( .I1(B[22]), .I2(n94), .O(n253) );
  OR_GATE U264 ( .I1(n94), .I2(B[22]), .O(n252) );
  AND_GATE U265 ( .I1(n254), .I2(n255), .O(SUM[21]) );
  NAND_GATE U266 ( .I1(n256), .I2(n251), .O(n255) );
  OR_GATE U267 ( .I1(n256), .I2(n251), .O(n254) );
  AND_GATE U268 ( .I1(n257), .I2(n258), .O(n251) );
  NAND_GATE U269 ( .I1(B[20]), .I2(n259), .O(n258) );
  NAND_GATE U270 ( .I1(n6), .I2(n267), .O(n259) );
  AND_GATE U271 ( .I1(n261), .I2(n262), .O(n256) );
  NAND_GATE U272 ( .I1(B[21]), .I2(n93), .O(n262) );
  OR_GATE U273 ( .I1(n93), .I2(B[21]), .O(n261) );
  AND_GATE U274 ( .I1(n263), .I2(n264), .O(SUM[20]) );
  NAND_GATE U275 ( .I1(n265), .I2(n260), .O(n264) );
  OR_GATE U276 ( .I1(n265), .I2(n260), .O(n263) );
  AND_GATE U277 ( .I1(n266), .I2(n267), .O(n260) );
  NAND_GATE U278 ( .I1(B[19]), .I2(n268), .O(n267) );
  NAND_GATE U279 ( .I1(n269), .I2(n91), .O(n268) );
  OR_GATE U280 ( .I1(n91), .I2(n269), .O(n266) );
  AND_GATE U281 ( .I1(n270), .I2(n271), .O(n265) );
  NAND_GATE U282 ( .I1(B[20]), .I2(n92), .O(n271) );
  OR_GATE U283 ( .I1(n92), .I2(B[20]), .O(n270) );
  AND_GATE U284 ( .I1(n272), .I2(n273), .O(SUM[1]) );
  NAND_GATE U285 ( .I1(n274), .I2(n275), .O(n273) );
  OR_GATE U286 ( .I1(n274), .I2(n275), .O(n272) );
  AND_GATE U287 ( .I1(n276), .I2(n277), .O(n274) );
  NAND_GATE U288 ( .I1(B[1]), .I2(n73), .O(n277) );
  OR_GATE U289 ( .I1(n73), .I2(B[1]), .O(n276) );
  AND_GATE U290 ( .I1(n278), .I2(n279), .O(SUM[19]) );
  NAND_GATE U291 ( .I1(n280), .I2(n269), .O(n279) );
  OR_GATE U292 ( .I1(n280), .I2(n269), .O(n278) );
  AND_GATE U293 ( .I1(n281), .I2(n282), .O(n269) );
  NAND_GATE U294 ( .I1(B[18]), .I2(n283), .O(n282) );
  NAND_GATE U295 ( .I1(n284), .I2(n90), .O(n283) );
  OR_GATE U296 ( .I1(n90), .I2(n284), .O(n281) );
  AND_GATE U297 ( .I1(n285), .I2(n286), .O(n280) );
  NAND_GATE U298 ( .I1(B[19]), .I2(n91), .O(n286) );
  OR_GATE U299 ( .I1(n91), .I2(B[19]), .O(n285) );
  AND_GATE U300 ( .I1(n287), .I2(n288), .O(SUM[18]) );
  NAND_GATE U301 ( .I1(n289), .I2(n284), .O(n288) );
  OR_GATE U302 ( .I1(n289), .I2(n284), .O(n287) );
  AND_GATE U303 ( .I1(n290), .I2(n291), .O(n284) );
  NAND_GATE U304 ( .I1(B[17]), .I2(n292), .O(n291) );
  NAND_GATE U305 ( .I1(n293), .I2(n89), .O(n292) );
  OR_GATE U306 ( .I1(n89), .I2(n293), .O(n290) );
  AND_GATE U307 ( .I1(n294), .I2(n295), .O(n289) );
  NAND_GATE U308 ( .I1(B[18]), .I2(n90), .O(n295) );
  OR_GATE U309 ( .I1(n90), .I2(B[18]), .O(n294) );
  AND_GATE U310 ( .I1(n296), .I2(n297), .O(SUM[17]) );
  NAND_GATE U311 ( .I1(n298), .I2(n293), .O(n297) );
  OR_GATE U312 ( .I1(n298), .I2(n293), .O(n296) );
  AND_GATE U313 ( .I1(n299), .I2(n300), .O(n293) );
  NAND_GATE U314 ( .I1(B[16]), .I2(n301), .O(n300) );
  NAND_GATE U315 ( .I1(n302), .I2(n88), .O(n301) );
  OR_GATE U316 ( .I1(n88), .I2(n302), .O(n299) );
  AND_GATE U317 ( .I1(n303), .I2(n304), .O(n298) );
  NAND_GATE U318 ( .I1(B[17]), .I2(n89), .O(n304) );
  OR_GATE U319 ( .I1(n89), .I2(B[17]), .O(n303) );
  AND_GATE U320 ( .I1(n305), .I2(n306), .O(SUM[16]) );
  NAND_GATE U321 ( .I1(n307), .I2(n302), .O(n306) );
  OR_GATE U322 ( .I1(n307), .I2(n302), .O(n305) );
  AND_GATE U323 ( .I1(n308), .I2(n309), .O(n302) );
  NAND_GATE U324 ( .I1(B[15]), .I2(n310), .O(n309) );
  NAND_GATE U325 ( .I1(n311), .I2(n87), .O(n310) );
  OR_GATE U326 ( .I1(n87), .I2(n311), .O(n308) );
  AND_GATE U327 ( .I1(n312), .I2(n313), .O(n307) );
  NAND_GATE U328 ( .I1(B[16]), .I2(n88), .O(n313) );
  OR_GATE U329 ( .I1(n88), .I2(B[16]), .O(n312) );
  AND_GATE U330 ( .I1(n314), .I2(n315), .O(SUM[15]) );
  NAND_GATE U331 ( .I1(n316), .I2(n311), .O(n315) );
  OR_GATE U332 ( .I1(n316), .I2(n311), .O(n314) );
  AND_GATE U333 ( .I1(n317), .I2(n318), .O(n311) );
  NAND_GATE U334 ( .I1(B[14]), .I2(n319), .O(n318) );
  NAND_GATE U335 ( .I1(n320), .I2(n86), .O(n319) );
  OR_GATE U336 ( .I1(n86), .I2(n320), .O(n317) );
  AND_GATE U337 ( .I1(n321), .I2(n322), .O(n316) );
  NAND_GATE U338 ( .I1(B[15]), .I2(n87), .O(n322) );
  OR_GATE U339 ( .I1(n87), .I2(B[15]), .O(n321) );
  AND_GATE U340 ( .I1(n323), .I2(n324), .O(SUM[14]) );
  NAND_GATE U341 ( .I1(n325), .I2(n320), .O(n324) );
  OR_GATE U342 ( .I1(n325), .I2(n320), .O(n323) );
  AND_GATE U343 ( .I1(n326), .I2(n327), .O(n320) );
  NAND_GATE U344 ( .I1(B[13]), .I2(n328), .O(n327) );
  NAND_GATE U345 ( .I1(n329), .I2(n85), .O(n328) );
  OR_GATE U346 ( .I1(n85), .I2(n329), .O(n326) );
  AND_GATE U347 ( .I1(n330), .I2(n331), .O(n325) );
  NAND_GATE U348 ( .I1(B[14]), .I2(n86), .O(n331) );
  OR_GATE U349 ( .I1(n86), .I2(B[14]), .O(n330) );
  AND_GATE U350 ( .I1(n332), .I2(n333), .O(SUM[13]) );
  NAND_GATE U351 ( .I1(n334), .I2(n329), .O(n333) );
  OR_GATE U352 ( .I1(n334), .I2(n329), .O(n332) );
  AND_GATE U353 ( .I1(n335), .I2(n336), .O(n329) );
  NAND_GATE U354 ( .I1(B[12]), .I2(n337), .O(n336) );
  NAND_GATE U355 ( .I1(n338), .I2(n84), .O(n337) );
  OR_GATE U356 ( .I1(n84), .I2(n338), .O(n335) );
  AND_GATE U357 ( .I1(n339), .I2(n340), .O(n334) );
  NAND_GATE U358 ( .I1(B[13]), .I2(n85), .O(n340) );
  OR_GATE U359 ( .I1(n85), .I2(B[13]), .O(n339) );
  AND_GATE U360 ( .I1(n341), .I2(n342), .O(SUM[12]) );
  NAND_GATE U361 ( .I1(n343), .I2(n338), .O(n342) );
  OR_GATE U362 ( .I1(n343), .I2(n338), .O(n341) );
  AND_GATE U363 ( .I1(n344), .I2(n345), .O(n338) );
  NAND_GATE U364 ( .I1(B[11]), .I2(n346), .O(n345) );
  NAND_GATE U365 ( .I1(n347), .I2(n83), .O(n346) );
  OR_GATE U366 ( .I1(n83), .I2(n347), .O(n344) );
  AND_GATE U367 ( .I1(n348), .I2(n349), .O(n343) );
  NAND_GATE U368 ( .I1(B[12]), .I2(n84), .O(n349) );
  OR_GATE U369 ( .I1(n84), .I2(B[12]), .O(n348) );
  AND_GATE U370 ( .I1(n350), .I2(n351), .O(SUM[11]) );
  NAND_GATE U371 ( .I1(n352), .I2(n347), .O(n351) );
  OR_GATE U372 ( .I1(n352), .I2(n347), .O(n350) );
  AND_GATE U373 ( .I1(n353), .I2(n354), .O(n347) );
  NAND_GATE U374 ( .I1(B[10]), .I2(n355), .O(n354) );
  NAND_GATE U375 ( .I1(n356), .I2(n82), .O(n355) );
  OR_GATE U376 ( .I1(n82), .I2(n356), .O(n353) );
  AND_GATE U377 ( .I1(n357), .I2(n358), .O(n352) );
  NAND_GATE U378 ( .I1(B[11]), .I2(n83), .O(n358) );
  OR_GATE U379 ( .I1(n83), .I2(B[11]), .O(n357) );
  AND_GATE U380 ( .I1(n359), .I2(n360), .O(SUM[10]) );
  NAND_GATE U381 ( .I1(n361), .I2(n356), .O(n360) );
  OR_GATE U382 ( .I1(n361), .I2(n356), .O(n359) );
  AND_GATE U383 ( .I1(n362), .I2(n363), .O(n356) );
  NAND_GATE U384 ( .I1(B[9]), .I2(n364), .O(n363) );
  NAND_GATE U385 ( .I1(n109), .I2(n81), .O(n364) );
  OR_GATE U386 ( .I1(n81), .I2(n109), .O(n362) );
  AND_GATE U387 ( .I1(n365), .I2(n366), .O(n109) );
  NAND_GATE U388 ( .I1(B[8]), .I2(n367), .O(n366) );
  NAND_GATE U389 ( .I1(n115), .I2(n80), .O(n367) );
  OR_GATE U390 ( .I1(n80), .I2(n115), .O(n365) );
  AND_GATE U391 ( .I1(n368), .I2(n369), .O(n115) );
  NAND_GATE U392 ( .I1(B[7]), .I2(n370), .O(n369) );
  NAND_GATE U393 ( .I1(n121), .I2(n79), .O(n370) );
  OR_GATE U394 ( .I1(n79), .I2(n121), .O(n368) );
  AND_GATE U395 ( .I1(n371), .I2(n372), .O(n121) );
  NAND_GATE U396 ( .I1(B[6]), .I2(n373), .O(n372) );
  NAND_GATE U397 ( .I1(n127), .I2(n78), .O(n373) );
  OR_GATE U398 ( .I1(n78), .I2(n127), .O(n371) );
  AND_GATE U399 ( .I1(n374), .I2(n375), .O(n127) );
  NAND_GATE U400 ( .I1(B[5]), .I2(n376), .O(n375) );
  NAND_GATE U401 ( .I1(n133), .I2(n77), .O(n376) );
  OR_GATE U402 ( .I1(n77), .I2(n133), .O(n374) );
  AND_GATE U403 ( .I1(n377), .I2(n378), .O(n133) );
  NAND_GATE U404 ( .I1(B[4]), .I2(n379), .O(n378) );
  NAND_GATE U405 ( .I1(n139), .I2(n76), .O(n379) );
  OR_GATE U406 ( .I1(n76), .I2(n139), .O(n377) );
  AND_GATE U407 ( .I1(n380), .I2(n381), .O(n139) );
  NAND_GATE U408 ( .I1(B[3]), .I2(n382), .O(n381) );
  NAND_GATE U409 ( .I1(n145), .I2(n75), .O(n382) );
  OR_GATE U410 ( .I1(n75), .I2(n145), .O(n380) );
  AND_GATE U411 ( .I1(n383), .I2(n384), .O(n145) );
  NAND_GATE U412 ( .I1(B[2]), .I2(n385), .O(n384) );
  NAND_GATE U413 ( .I1(n179), .I2(n74), .O(n385) );
  OR_GATE U414 ( .I1(n74), .I2(n179), .O(n383) );
  AND_GATE U415 ( .I1(n386), .I2(n387), .O(n179) );
  NAND_GATE U416 ( .I1(B[1]), .I2(n388), .O(n387) );
  NAND_GATE U417 ( .I1(n275), .I2(n73), .O(n388) );
  OR_GATE U418 ( .I1(n73), .I2(n275), .O(n386) );
  AND_GATE U419 ( .I1(n389), .I2(n390), .O(n275) );
  NAND_GATE U420 ( .I1(CI), .I2(n391), .O(n390) );
  OR_GATE U421 ( .I1(A[0]), .I2(B[0]), .O(n391) );
  NAND_GATE U422 ( .I1(B[0]), .I2(A[0]), .O(n389) );
  AND_GATE U423 ( .I1(n392), .I2(n393), .O(n361) );
  NAND_GATE U424 ( .I1(B[10]), .I2(n82), .O(n393) );
  OR_GATE U425 ( .I1(n82), .I2(B[10]), .O(n392) );
  NAND_GATE U426 ( .I1(n394), .I2(n395), .O(SUM[0]) );
  NAND_GATE U427 ( .I1(n396), .I2(A[0]), .O(n395) );
  OR_GATE U428 ( .I1(n396), .I2(A[0]), .O(n394) );
  AND_GATE U429 ( .I1(n397), .I2(n398), .O(n396) );
  NAND_GATE U430 ( .I1(CI), .I2(n105), .O(n398) );
  OR_GATE U431 ( .I1(n105), .I2(CI), .O(n397) );
endmodule


module pps_ex_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_GATE U1 ( .I1(A[30]), .O(n1) );
  INV_GATE U2 ( .I1(A[29]), .O(n2) );
  INV_GATE U3 ( .I1(A[28]), .O(n3) );
  INV_GATE U4 ( .I1(A[27]), .O(n4) );
  INV_GATE U5 ( .I1(A[26]), .O(n5) );
  INV_GATE U6 ( .I1(A[25]), .O(n6) );
  INV_GATE U7 ( .I1(A[24]), .O(n7) );
  INV_GATE U8 ( .I1(A[23]), .O(n8) );
  INV_GATE U9 ( .I1(A[22]), .O(n9) );
  INV_GATE U10 ( .I1(A[21]), .O(n10) );
  INV_GATE U11 ( .I1(A[20]), .O(n11) );
  INV_GATE U12 ( .I1(A[19]), .O(n12) );
  INV_GATE U13 ( .I1(A[18]), .O(n13) );
  INV_GATE U14 ( .I1(A[17]), .O(n14) );
  INV_GATE U15 ( .I1(A[16]), .O(n15) );
  INV_GATE U16 ( .I1(A[15]), .O(n16) );
  INV_GATE U17 ( .I1(A[14]), .O(n17) );
  INV_GATE U18 ( .I1(A[13]), .O(n18) );
  INV_GATE U19 ( .I1(A[12]), .O(n19) );
  INV_GATE U20 ( .I1(A[11]), .O(n20) );
  INV_GATE U21 ( .I1(n112), .O(n21) );
  INV_GATE U22 ( .I1(A[8]), .O(n22) );
  INV_GATE U23 ( .I1(n32), .O(n23) );
  INV_GATE U24 ( .I1(A[7]), .O(n24) );
  INV_GATE U25 ( .I1(A[6]), .O(n25) );
  INV_GATE U26 ( .I1(A[5]), .O(n26) );
  INV_GATE U27 ( .I1(A[4]), .O(n27) );
  INV_GATE U28 ( .I1(A[3]), .O(n28) );
  INV_GATE U29 ( .I1(A[2]), .O(SUM[2]) );
  NAND_GATE U30 ( .I1(n30), .I2(n31), .O(SUM[9]) );
  NAND_GATE U31 ( .I1(A[9]), .I2(n23), .O(n31) );
  OR_GATE U32 ( .I1(n23), .I2(A[9]), .O(n30) );
  NAND_GATE U33 ( .I1(n33), .I2(n34), .O(SUM[8]) );
  OR_GATE U34 ( .I1(n22), .I2(n35), .O(n34) );
  NAND_GATE U35 ( .I1(n35), .I2(n22), .O(n33) );
  AND_GATE U36 ( .I1(A[7]), .I2(n36), .O(n35) );
  NAND_GATE U37 ( .I1(n37), .I2(n38), .O(SUM[7]) );
  OR_GATE U38 ( .I1(n24), .I2(n36), .O(n38) );
  NAND_GATE U39 ( .I1(n36), .I2(n24), .O(n37) );
  NAND_GATE U40 ( .I1(n39), .I2(n40), .O(SUM[6]) );
  OR_GATE U41 ( .I1(n25), .I2(n41), .O(n40) );
  NAND_GATE U42 ( .I1(n41), .I2(n25), .O(n39) );
  AND_GATE U43 ( .I1(A[5]), .I2(n42), .O(n41) );
  NAND_GATE U44 ( .I1(n43), .I2(n44), .O(SUM[5]) );
  OR_GATE U45 ( .I1(n26), .I2(n42), .O(n44) );
  NAND_GATE U46 ( .I1(n42), .I2(n26), .O(n43) );
  NAND_GATE U47 ( .I1(n45), .I2(n46), .O(SUM[4]) );
  OR_GATE U48 ( .I1(n27), .I2(n47), .O(n46) );
  NAND_GATE U49 ( .I1(n47), .I2(n27), .O(n45) );
  AND_GATE U50 ( .I1(A[3]), .I2(A[2]), .O(n47) );
  NAND_GATE U51 ( .I1(n48), .I2(n49), .O(SUM[3]) );
  NAND_GATE U52 ( .I1(A[3]), .I2(SUM[2]), .O(n49) );
  NAND_GATE U53 ( .I1(A[2]), .I2(n28), .O(n48) );
  NAND_GATE U54 ( .I1(n50), .I2(n51), .O(SUM[31]) );
  NAND_GATE U55 ( .I1(A[31]), .I2(n52), .O(n51) );
  OR_GATE U56 ( .I1(n52), .I2(A[31]), .O(n50) );
  NAND_GATE U57 ( .I1(A[30]), .I2(n53), .O(n52) );
  NAND_GATE U58 ( .I1(n54), .I2(n55), .O(SUM[30]) );
  OR_GATE U59 ( .I1(n1), .I2(n53), .O(n55) );
  NAND_GATE U60 ( .I1(n53), .I2(n1), .O(n54) );
  AND_GATE U61 ( .I1(A[29]), .I2(n56), .O(n53) );
  NAND_GATE U62 ( .I1(n57), .I2(n58), .O(SUM[29]) );
  OR_GATE U63 ( .I1(n2), .I2(n56), .O(n58) );
  NAND_GATE U64 ( .I1(n56), .I2(n2), .O(n57) );
  AND3_GATE U65 ( .I1(A[27]), .I2(n59), .I3(A[28]), .O(n56) );
  NAND_GATE U66 ( .I1(n60), .I2(n61), .O(SUM[28]) );
  OR_GATE U67 ( .I1(n3), .I2(n62), .O(n61) );
  NAND_GATE U68 ( .I1(n62), .I2(n3), .O(n60) );
  AND_GATE U69 ( .I1(A[27]), .I2(n59), .O(n62) );
  NAND_GATE U70 ( .I1(n63), .I2(n64), .O(SUM[27]) );
  OR_GATE U71 ( .I1(n4), .I2(n59), .O(n64) );
  NAND_GATE U72 ( .I1(n59), .I2(n4), .O(n63) );
  AND3_GATE U73 ( .I1(A[25]), .I2(n65), .I3(A[26]), .O(n59) );
  NAND_GATE U74 ( .I1(n66), .I2(n67), .O(SUM[26]) );
  OR_GATE U75 ( .I1(n5), .I2(n68), .O(n67) );
  NAND_GATE U76 ( .I1(n68), .I2(n5), .O(n66) );
  AND_GATE U77 ( .I1(A[25]), .I2(n65), .O(n68) );
  NAND_GATE U78 ( .I1(n69), .I2(n70), .O(SUM[25]) );
  OR_GATE U79 ( .I1(n6), .I2(n65), .O(n70) );
  NAND_GATE U80 ( .I1(n65), .I2(n6), .O(n69) );
  AND3_GATE U81 ( .I1(A[23]), .I2(n71), .I3(A[24]), .O(n65) );
  NAND_GATE U82 ( .I1(n72), .I2(n73), .O(SUM[24]) );
  OR_GATE U83 ( .I1(n7), .I2(n74), .O(n73) );
  NAND_GATE U84 ( .I1(n74), .I2(n7), .O(n72) );
  AND_GATE U85 ( .I1(A[23]), .I2(n71), .O(n74) );
  NAND_GATE U86 ( .I1(n75), .I2(n76), .O(SUM[23]) );
  OR_GATE U87 ( .I1(n8), .I2(n71), .O(n76) );
  NAND_GATE U88 ( .I1(n71), .I2(n8), .O(n75) );
  AND3_GATE U89 ( .I1(A[21]), .I2(n77), .I3(A[22]), .O(n71) );
  NAND_GATE U90 ( .I1(n78), .I2(n79), .O(SUM[22]) );
  OR_GATE U91 ( .I1(n9), .I2(n80), .O(n79) );
  NAND_GATE U92 ( .I1(n80), .I2(n9), .O(n78) );
  AND_GATE U93 ( .I1(A[21]), .I2(n77), .O(n80) );
  NAND_GATE U94 ( .I1(n81), .I2(n82), .O(SUM[21]) );
  OR_GATE U95 ( .I1(n10), .I2(n77), .O(n82) );
  NAND_GATE U96 ( .I1(n77), .I2(n10), .O(n81) );
  AND3_GATE U97 ( .I1(A[19]), .I2(n83), .I3(A[20]), .O(n77) );
  NAND_GATE U98 ( .I1(n84), .I2(n85), .O(SUM[20]) );
  OR_GATE U99 ( .I1(n11), .I2(n86), .O(n85) );
  NAND_GATE U100 ( .I1(n86), .I2(n11), .O(n84) );
  AND_GATE U101 ( .I1(A[19]), .I2(n83), .O(n86) );
  NAND_GATE U102 ( .I1(n87), .I2(n88), .O(SUM[19]) );
  OR_GATE U103 ( .I1(n12), .I2(n83), .O(n88) );
  NAND_GATE U104 ( .I1(n83), .I2(n12), .O(n87) );
  AND3_GATE U105 ( .I1(A[17]), .I2(n89), .I3(A[18]), .O(n83) );
  NAND_GATE U106 ( .I1(n90), .I2(n91), .O(SUM[18]) );
  OR_GATE U107 ( .I1(n13), .I2(n92), .O(n91) );
  NAND_GATE U108 ( .I1(n92), .I2(n13), .O(n90) );
  AND_GATE U109 ( .I1(A[17]), .I2(n89), .O(n92) );
  NAND_GATE U110 ( .I1(n93), .I2(n94), .O(SUM[17]) );
  OR_GATE U111 ( .I1(n14), .I2(n89), .O(n94) );
  NAND_GATE U112 ( .I1(n89), .I2(n14), .O(n93) );
  AND3_GATE U113 ( .I1(A[15]), .I2(n95), .I3(A[16]), .O(n89) );
  NAND_GATE U114 ( .I1(n96), .I2(n97), .O(SUM[16]) );
  OR_GATE U115 ( .I1(n15), .I2(n98), .O(n97) );
  NAND_GATE U116 ( .I1(n98), .I2(n15), .O(n96) );
  AND_GATE U117 ( .I1(A[15]), .I2(n95), .O(n98) );
  NAND_GATE U118 ( .I1(n99), .I2(n100), .O(SUM[15]) );
  OR_GATE U119 ( .I1(n16), .I2(n95), .O(n100) );
  NAND_GATE U120 ( .I1(n95), .I2(n16), .O(n99) );
  AND3_GATE U121 ( .I1(A[13]), .I2(n101), .I3(A[14]), .O(n95) );
  NAND_GATE U122 ( .I1(n102), .I2(n103), .O(SUM[14]) );
  OR_GATE U123 ( .I1(n17), .I2(n104), .O(n103) );
  NAND_GATE U124 ( .I1(n104), .I2(n17), .O(n102) );
  AND_GATE U125 ( .I1(A[13]), .I2(n101), .O(n104) );
  NAND_GATE U126 ( .I1(n105), .I2(n106), .O(SUM[13]) );
  OR_GATE U127 ( .I1(n18), .I2(n101), .O(n106) );
  NAND_GATE U128 ( .I1(n101), .I2(n18), .O(n105) );
  AND3_GATE U129 ( .I1(A[11]), .I2(n21), .I3(A[12]), .O(n101) );
  NAND_GATE U130 ( .I1(n107), .I2(n108), .O(SUM[12]) );
  OR_GATE U131 ( .I1(n19), .I2(n109), .O(n108) );
  NAND_GATE U132 ( .I1(n109), .I2(n19), .O(n107) );
  AND_GATE U133 ( .I1(A[11]), .I2(n21), .O(n109) );
  NAND_GATE U134 ( .I1(n110), .I2(n111), .O(SUM[11]) );
  NAND_GATE U135 ( .I1(A[11]), .I2(n112), .O(n111) );
  NAND_GATE U136 ( .I1(n21), .I2(n20), .O(n110) );
  NAND3_GATE U137 ( .I1(n32), .I2(A[9]), .I3(A[10]), .O(n112) );
  NAND_GATE U138 ( .I1(n113), .I2(n114), .O(SUM[10]) );
  NAND_GATE U139 ( .I1(A[10]), .I2(n115), .O(n114) );
  OR_GATE U140 ( .I1(n115), .I2(A[10]), .O(n113) );
  NAND_GATE U141 ( .I1(n32), .I2(A[9]), .O(n115) );
  AND3_GATE U142 ( .I1(A[7]), .I2(n36), .I3(A[8]), .O(n32) );
  AND3_GATE U143 ( .I1(A[5]), .I2(n42), .I3(A[6]), .O(n36) );
  AND3_GATE U144 ( .I1(A[3]), .I2(A[2]), .I3(A[4]), .O(n42) );
endmodule


module pps_ex_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310;

  INV_GATE U1 ( .I1(B[0]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[1]), .O(n32) );
  AND_GATE U33 ( .I1(n33), .I2(n34), .O(SUM[9]) );
  NAND_GATE U34 ( .I1(n35), .I2(n36), .O(n34) );
  OR_GATE U35 ( .I1(n35), .I2(n36), .O(n33) );
  AND_GATE U36 ( .I1(n37), .I2(n38), .O(n35) );
  NAND_GATE U37 ( .I1(B[9]), .I2(n24), .O(n38) );
  OR_GATE U38 ( .I1(n24), .I2(B[9]), .O(n37) );
  AND_GATE U39 ( .I1(n39), .I2(n40), .O(SUM[8]) );
  NAND_GATE U40 ( .I1(n41), .I2(n42), .O(n40) );
  OR_GATE U41 ( .I1(n41), .I2(n42), .O(n39) );
  AND_GATE U42 ( .I1(n43), .I2(n44), .O(n41) );
  NAND_GATE U43 ( .I1(B[8]), .I2(n25), .O(n44) );
  OR_GATE U44 ( .I1(n25), .I2(B[8]), .O(n43) );
  AND_GATE U45 ( .I1(n45), .I2(n46), .O(SUM[7]) );
  NAND_GATE U46 ( .I1(n47), .I2(n48), .O(n46) );
  OR_GATE U47 ( .I1(n47), .I2(n48), .O(n45) );
  AND_GATE U48 ( .I1(n49), .I2(n50), .O(n47) );
  NAND_GATE U49 ( .I1(B[7]), .I2(n26), .O(n50) );
  OR_GATE U50 ( .I1(n26), .I2(B[7]), .O(n49) );
  AND_GATE U51 ( .I1(n51), .I2(n52), .O(SUM[6]) );
  NAND_GATE U52 ( .I1(n53), .I2(n54), .O(n52) );
  OR_GATE U53 ( .I1(n53), .I2(n54), .O(n51) );
  AND_GATE U54 ( .I1(n55), .I2(n56), .O(n53) );
  NAND_GATE U55 ( .I1(B[6]), .I2(n27), .O(n56) );
  OR_GATE U56 ( .I1(n27), .I2(B[6]), .O(n55) );
  AND_GATE U57 ( .I1(n57), .I2(n58), .O(SUM[5]) );
  NAND_GATE U58 ( .I1(n59), .I2(n60), .O(n58) );
  OR_GATE U59 ( .I1(n59), .I2(n60), .O(n57) );
  AND_GATE U60 ( .I1(n61), .I2(n62), .O(n59) );
  NAND_GATE U61 ( .I1(B[5]), .I2(n28), .O(n62) );
  OR_GATE U62 ( .I1(n28), .I2(B[5]), .O(n61) );
  AND_GATE U63 ( .I1(n63), .I2(n64), .O(SUM[4]) );
  NAND_GATE U64 ( .I1(n65), .I2(n66), .O(n64) );
  OR_GATE U65 ( .I1(n65), .I2(n66), .O(n63) );
  AND_GATE U66 ( .I1(n67), .I2(n68), .O(n65) );
  NAND_GATE U67 ( .I1(B[4]), .I2(n29), .O(n68) );
  OR_GATE U68 ( .I1(n29), .I2(B[4]), .O(n67) );
  AND_GATE U69 ( .I1(n69), .I2(n70), .O(SUM[3]) );
  NAND_GATE U70 ( .I1(n71), .I2(n72), .O(n70) );
  OR_GATE U71 ( .I1(n71), .I2(n72), .O(n69) );
  AND_GATE U72 ( .I1(n73), .I2(n74), .O(n71) );
  NAND_GATE U73 ( .I1(B[3]), .I2(n30), .O(n74) );
  OR_GATE U74 ( .I1(n30), .I2(B[3]), .O(n73) );
  AND_GATE U75 ( .I1(n75), .I2(n76), .O(SUM[31]) );
  NAND_GATE U76 ( .I1(n77), .I2(n78), .O(n76) );
  OR_GATE U77 ( .I1(n78), .I2(n77), .O(n75) );
  AND_GATE U78 ( .I1(n79), .I2(n80), .O(n77) );
  NAND_GATE U79 ( .I1(B[30]), .I2(n81), .O(n80) );
  NAND_GATE U80 ( .I1(n82), .I2(n3), .O(n81) );
  OR_GATE U81 ( .I1(n3), .I2(n82), .O(n79) );
  AND_GATE U82 ( .I1(n83), .I2(n84), .O(n78) );
  NAND_GATE U83 ( .I1(B[31]), .I2(n2), .O(n84) );
  OR_GATE U84 ( .I1(n2), .I2(B[31]), .O(n83) );
  AND_GATE U85 ( .I1(n85), .I2(n86), .O(SUM[30]) );
  NAND_GATE U86 ( .I1(n87), .I2(n82), .O(n86) );
  OR_GATE U87 ( .I1(n87), .I2(n82), .O(n85) );
  AND_GATE U88 ( .I1(n88), .I2(n89), .O(n82) );
  NAND_GATE U89 ( .I1(B[29]), .I2(n90), .O(n89) );
  NAND_GATE U90 ( .I1(n91), .I2(n4), .O(n90) );
  OR_GATE U91 ( .I1(n4), .I2(n91), .O(n88) );
  AND_GATE U92 ( .I1(n92), .I2(n93), .O(n87) );
  NAND_GATE U93 ( .I1(B[30]), .I2(n3), .O(n93) );
  OR_GATE U94 ( .I1(n3), .I2(B[30]), .O(n92) );
  AND_GATE U95 ( .I1(n94), .I2(n95), .O(SUM[2]) );
  NAND_GATE U96 ( .I1(n96), .I2(n97), .O(n95) );
  OR_GATE U97 ( .I1(n96), .I2(n97), .O(n94) );
  AND_GATE U98 ( .I1(n98), .I2(n99), .O(n96) );
  NAND_GATE U99 ( .I1(B[2]), .I2(n31), .O(n99) );
  OR_GATE U100 ( .I1(n31), .I2(B[2]), .O(n98) );
  AND_GATE U101 ( .I1(n100), .I2(n101), .O(SUM[29]) );
  NAND_GATE U102 ( .I1(n102), .I2(n91), .O(n101) );
  OR_GATE U103 ( .I1(n102), .I2(n91), .O(n100) );
  AND_GATE U104 ( .I1(n103), .I2(n104), .O(n91) );
  NAND_GATE U105 ( .I1(B[28]), .I2(n105), .O(n104) );
  NAND_GATE U106 ( .I1(n106), .I2(n5), .O(n105) );
  OR_GATE U107 ( .I1(n5), .I2(n106), .O(n103) );
  AND_GATE U108 ( .I1(n107), .I2(n108), .O(n102) );
  NAND_GATE U109 ( .I1(B[29]), .I2(n4), .O(n108) );
  OR_GATE U110 ( .I1(n4), .I2(B[29]), .O(n107) );
  AND_GATE U111 ( .I1(n109), .I2(n110), .O(SUM[28]) );
  NAND_GATE U112 ( .I1(n111), .I2(n106), .O(n110) );
  OR_GATE U113 ( .I1(n111), .I2(n106), .O(n109) );
  AND_GATE U114 ( .I1(n112), .I2(n113), .O(n106) );
  NAND_GATE U115 ( .I1(B[27]), .I2(n114), .O(n113) );
  NAND_GATE U116 ( .I1(n115), .I2(n6), .O(n114) );
  OR_GATE U117 ( .I1(n6), .I2(n115), .O(n112) );
  AND_GATE U118 ( .I1(n116), .I2(n117), .O(n111) );
  NAND_GATE U119 ( .I1(B[28]), .I2(n5), .O(n117) );
  OR_GATE U120 ( .I1(n5), .I2(B[28]), .O(n116) );
  AND_GATE U121 ( .I1(n118), .I2(n119), .O(SUM[27]) );
  NAND_GATE U122 ( .I1(n120), .I2(n115), .O(n119) );
  OR_GATE U123 ( .I1(n120), .I2(n115), .O(n118) );
  AND_GATE U124 ( .I1(n121), .I2(n122), .O(n115) );
  NAND_GATE U125 ( .I1(B[26]), .I2(n123), .O(n122) );
  NAND_GATE U126 ( .I1(n124), .I2(n7), .O(n123) );
  OR_GATE U127 ( .I1(n7), .I2(n124), .O(n121) );
  AND_GATE U128 ( .I1(n125), .I2(n126), .O(n120) );
  NAND_GATE U129 ( .I1(B[27]), .I2(n6), .O(n126) );
  OR_GATE U130 ( .I1(n6), .I2(B[27]), .O(n125) );
  AND_GATE U131 ( .I1(n127), .I2(n128), .O(SUM[26]) );
  NAND_GATE U132 ( .I1(n129), .I2(n124), .O(n128) );
  OR_GATE U133 ( .I1(n129), .I2(n124), .O(n127) );
  AND_GATE U134 ( .I1(n130), .I2(n131), .O(n124) );
  NAND_GATE U135 ( .I1(B[25]), .I2(n132), .O(n131) );
  NAND_GATE U136 ( .I1(n133), .I2(n8), .O(n132) );
  OR_GATE U137 ( .I1(n8), .I2(n133), .O(n130) );
  AND_GATE U138 ( .I1(n134), .I2(n135), .O(n129) );
  NAND_GATE U139 ( .I1(B[26]), .I2(n7), .O(n135) );
  OR_GATE U140 ( .I1(n7), .I2(B[26]), .O(n134) );
  AND_GATE U141 ( .I1(n136), .I2(n137), .O(SUM[25]) );
  NAND_GATE U142 ( .I1(n138), .I2(n133), .O(n137) );
  OR_GATE U143 ( .I1(n138), .I2(n133), .O(n136) );
  AND_GATE U144 ( .I1(n139), .I2(n140), .O(n133) );
  NAND_GATE U145 ( .I1(B[24]), .I2(n141), .O(n140) );
  NAND_GATE U146 ( .I1(n142), .I2(n9), .O(n141) );
  OR_GATE U147 ( .I1(n9), .I2(n142), .O(n139) );
  AND_GATE U148 ( .I1(n143), .I2(n144), .O(n138) );
  NAND_GATE U149 ( .I1(B[25]), .I2(n8), .O(n144) );
  OR_GATE U150 ( .I1(n8), .I2(B[25]), .O(n143) );
  AND_GATE U151 ( .I1(n145), .I2(n146), .O(SUM[24]) );
  NAND_GATE U152 ( .I1(n147), .I2(n142), .O(n146) );
  OR_GATE U153 ( .I1(n147), .I2(n142), .O(n145) );
  AND_GATE U154 ( .I1(n148), .I2(n149), .O(n142) );
  NAND_GATE U155 ( .I1(B[23]), .I2(n150), .O(n149) );
  NAND_GATE U156 ( .I1(n151), .I2(n10), .O(n150) );
  OR_GATE U157 ( .I1(n10), .I2(n151), .O(n148) );
  AND_GATE U158 ( .I1(n152), .I2(n153), .O(n147) );
  NAND_GATE U159 ( .I1(B[24]), .I2(n9), .O(n153) );
  OR_GATE U160 ( .I1(n9), .I2(B[24]), .O(n152) );
  AND_GATE U161 ( .I1(n154), .I2(n155), .O(SUM[23]) );
  NAND_GATE U162 ( .I1(n156), .I2(n151), .O(n155) );
  OR_GATE U163 ( .I1(n156), .I2(n151), .O(n154) );
  AND_GATE U164 ( .I1(n157), .I2(n158), .O(n151) );
  NAND_GATE U165 ( .I1(B[22]), .I2(n159), .O(n158) );
  NAND_GATE U166 ( .I1(n160), .I2(n11), .O(n159) );
  OR_GATE U167 ( .I1(n11), .I2(n160), .O(n157) );
  AND_GATE U168 ( .I1(n161), .I2(n162), .O(n156) );
  NAND_GATE U169 ( .I1(B[23]), .I2(n10), .O(n162) );
  OR_GATE U170 ( .I1(n10), .I2(B[23]), .O(n161) );
  AND_GATE U171 ( .I1(n163), .I2(n164), .O(SUM[22]) );
  NAND_GATE U172 ( .I1(n165), .I2(n160), .O(n164) );
  OR_GATE U173 ( .I1(n165), .I2(n160), .O(n163) );
  AND_GATE U174 ( .I1(n166), .I2(n167), .O(n160) );
  NAND_GATE U175 ( .I1(B[21]), .I2(n168), .O(n167) );
  NAND_GATE U176 ( .I1(n169), .I2(n12), .O(n168) );
  OR_GATE U177 ( .I1(n12), .I2(n169), .O(n166) );
  AND_GATE U178 ( .I1(n170), .I2(n171), .O(n165) );
  NAND_GATE U179 ( .I1(B[22]), .I2(n11), .O(n171) );
  OR_GATE U180 ( .I1(n11), .I2(B[22]), .O(n170) );
  AND_GATE U181 ( .I1(n172), .I2(n173), .O(SUM[21]) );
  NAND_GATE U182 ( .I1(n174), .I2(n169), .O(n173) );
  OR_GATE U183 ( .I1(n174), .I2(n169), .O(n172) );
  AND_GATE U184 ( .I1(n175), .I2(n176), .O(n169) );
  NAND_GATE U185 ( .I1(B[20]), .I2(n177), .O(n176) );
  NAND_GATE U186 ( .I1(n178), .I2(n13), .O(n177) );
  OR_GATE U187 ( .I1(n13), .I2(n178), .O(n175) );
  AND_GATE U188 ( .I1(n179), .I2(n180), .O(n174) );
  NAND_GATE U189 ( .I1(B[21]), .I2(n12), .O(n180) );
  OR_GATE U190 ( .I1(n12), .I2(B[21]), .O(n179) );
  AND_GATE U191 ( .I1(n181), .I2(n182), .O(SUM[20]) );
  NAND_GATE U192 ( .I1(n183), .I2(n178), .O(n182) );
  OR_GATE U193 ( .I1(n183), .I2(n178), .O(n181) );
  AND_GATE U194 ( .I1(n184), .I2(n185), .O(n178) );
  NAND_GATE U195 ( .I1(B[19]), .I2(n186), .O(n185) );
  NAND_GATE U196 ( .I1(n187), .I2(n14), .O(n186) );
  OR_GATE U197 ( .I1(n14), .I2(n187), .O(n184) );
  AND_GATE U198 ( .I1(n188), .I2(n189), .O(n183) );
  NAND_GATE U199 ( .I1(B[20]), .I2(n13), .O(n189) );
  OR_GATE U200 ( .I1(n13), .I2(B[20]), .O(n188) );
  NAND_GATE U201 ( .I1(n190), .I2(n191), .O(SUM[1]) );
  NAND_GATE U202 ( .I1(n192), .I2(n193), .O(n191) );
  OR_GATE U203 ( .I1(n192), .I2(n193), .O(n190) );
  AND_GATE U204 ( .I1(n194), .I2(n195), .O(n192) );
  NAND_GATE U205 ( .I1(B[1]), .I2(n32), .O(n195) );
  OR_GATE U206 ( .I1(n32), .I2(B[1]), .O(n194) );
  AND_GATE U207 ( .I1(n196), .I2(n197), .O(SUM[19]) );
  NAND_GATE U208 ( .I1(n198), .I2(n187), .O(n197) );
  OR_GATE U209 ( .I1(n198), .I2(n187), .O(n196) );
  AND_GATE U210 ( .I1(n199), .I2(n200), .O(n187) );
  NAND_GATE U211 ( .I1(B[18]), .I2(n201), .O(n200) );
  NAND_GATE U212 ( .I1(n202), .I2(n15), .O(n201) );
  OR_GATE U213 ( .I1(n15), .I2(n202), .O(n199) );
  AND_GATE U214 ( .I1(n203), .I2(n204), .O(n198) );
  NAND_GATE U215 ( .I1(B[19]), .I2(n14), .O(n204) );
  OR_GATE U216 ( .I1(n14), .I2(B[19]), .O(n203) );
  AND_GATE U217 ( .I1(n205), .I2(n206), .O(SUM[18]) );
  NAND_GATE U218 ( .I1(n207), .I2(n202), .O(n206) );
  OR_GATE U219 ( .I1(n207), .I2(n202), .O(n205) );
  AND_GATE U220 ( .I1(n208), .I2(n209), .O(n202) );
  NAND_GATE U221 ( .I1(B[17]), .I2(n210), .O(n209) );
  NAND_GATE U222 ( .I1(n211), .I2(n16), .O(n210) );
  OR_GATE U223 ( .I1(n16), .I2(n211), .O(n208) );
  AND_GATE U224 ( .I1(n212), .I2(n213), .O(n207) );
  NAND_GATE U225 ( .I1(B[18]), .I2(n15), .O(n213) );
  OR_GATE U226 ( .I1(n15), .I2(B[18]), .O(n212) );
  AND_GATE U227 ( .I1(n214), .I2(n215), .O(SUM[17]) );
  NAND_GATE U228 ( .I1(n216), .I2(n211), .O(n215) );
  OR_GATE U229 ( .I1(n216), .I2(n211), .O(n214) );
  AND_GATE U230 ( .I1(n217), .I2(n218), .O(n211) );
  NAND_GATE U231 ( .I1(B[16]), .I2(n219), .O(n218) );
  NAND_GATE U232 ( .I1(n220), .I2(n17), .O(n219) );
  OR_GATE U233 ( .I1(n17), .I2(n220), .O(n217) );
  AND_GATE U234 ( .I1(n221), .I2(n222), .O(n216) );
  NAND_GATE U235 ( .I1(B[17]), .I2(n16), .O(n222) );
  OR_GATE U236 ( .I1(n16), .I2(B[17]), .O(n221) );
  AND_GATE U237 ( .I1(n223), .I2(n224), .O(SUM[16]) );
  NAND_GATE U238 ( .I1(n225), .I2(n220), .O(n224) );
  OR_GATE U239 ( .I1(n225), .I2(n220), .O(n223) );
  AND_GATE U240 ( .I1(n226), .I2(n227), .O(n220) );
  NAND_GATE U241 ( .I1(B[15]), .I2(n228), .O(n227) );
  NAND_GATE U242 ( .I1(n229), .I2(n18), .O(n228) );
  OR_GATE U243 ( .I1(n18), .I2(n229), .O(n226) );
  AND_GATE U244 ( .I1(n230), .I2(n231), .O(n225) );
  NAND_GATE U245 ( .I1(B[16]), .I2(n17), .O(n231) );
  OR_GATE U246 ( .I1(n17), .I2(B[16]), .O(n230) );
  AND_GATE U247 ( .I1(n232), .I2(n233), .O(SUM[15]) );
  NAND_GATE U248 ( .I1(n234), .I2(n229), .O(n233) );
  OR_GATE U249 ( .I1(n234), .I2(n229), .O(n232) );
  AND_GATE U250 ( .I1(n235), .I2(n236), .O(n229) );
  NAND_GATE U251 ( .I1(B[14]), .I2(n237), .O(n236) );
  NAND_GATE U252 ( .I1(n238), .I2(n19), .O(n237) );
  OR_GATE U253 ( .I1(n19), .I2(n238), .O(n235) );
  AND_GATE U254 ( .I1(n239), .I2(n240), .O(n234) );
  NAND_GATE U255 ( .I1(B[15]), .I2(n18), .O(n240) );
  OR_GATE U256 ( .I1(n18), .I2(B[15]), .O(n239) );
  AND_GATE U257 ( .I1(n241), .I2(n242), .O(SUM[14]) );
  NAND_GATE U258 ( .I1(n243), .I2(n238), .O(n242) );
  OR_GATE U259 ( .I1(n243), .I2(n238), .O(n241) );
  AND_GATE U260 ( .I1(n244), .I2(n245), .O(n238) );
  NAND_GATE U261 ( .I1(B[13]), .I2(n246), .O(n245) );
  NAND_GATE U262 ( .I1(n247), .I2(n20), .O(n246) );
  OR_GATE U263 ( .I1(n20), .I2(n247), .O(n244) );
  AND_GATE U264 ( .I1(n248), .I2(n249), .O(n243) );
  NAND_GATE U265 ( .I1(B[14]), .I2(n19), .O(n249) );
  OR_GATE U266 ( .I1(n19), .I2(B[14]), .O(n248) );
  AND_GATE U267 ( .I1(n250), .I2(n251), .O(SUM[13]) );
  NAND_GATE U268 ( .I1(n252), .I2(n247), .O(n251) );
  OR_GATE U269 ( .I1(n252), .I2(n247), .O(n250) );
  AND_GATE U270 ( .I1(n253), .I2(n254), .O(n247) );
  NAND_GATE U271 ( .I1(B[12]), .I2(n255), .O(n254) );
  NAND_GATE U272 ( .I1(n256), .I2(n21), .O(n255) );
  OR_GATE U273 ( .I1(n21), .I2(n256), .O(n253) );
  AND_GATE U274 ( .I1(n257), .I2(n258), .O(n252) );
  NAND_GATE U275 ( .I1(B[13]), .I2(n20), .O(n258) );
  OR_GATE U276 ( .I1(n20), .I2(B[13]), .O(n257) );
  AND_GATE U277 ( .I1(n259), .I2(n260), .O(SUM[12]) );
  NAND_GATE U278 ( .I1(n261), .I2(n256), .O(n260) );
  OR_GATE U279 ( .I1(n261), .I2(n256), .O(n259) );
  AND_GATE U280 ( .I1(n262), .I2(n263), .O(n256) );
  NAND_GATE U281 ( .I1(B[11]), .I2(n264), .O(n263) );
  NAND_GATE U282 ( .I1(n265), .I2(n22), .O(n264) );
  OR_GATE U283 ( .I1(n22), .I2(n265), .O(n262) );
  AND_GATE U284 ( .I1(n266), .I2(n267), .O(n261) );
  NAND_GATE U285 ( .I1(B[12]), .I2(n21), .O(n267) );
  OR_GATE U286 ( .I1(n21), .I2(B[12]), .O(n266) );
  AND_GATE U287 ( .I1(n268), .I2(n269), .O(SUM[11]) );
  NAND_GATE U288 ( .I1(n270), .I2(n265), .O(n269) );
  OR_GATE U289 ( .I1(n270), .I2(n265), .O(n268) );
  AND_GATE U290 ( .I1(n271), .I2(n272), .O(n265) );
  NAND_GATE U291 ( .I1(B[10]), .I2(n273), .O(n272) );
  NAND_GATE U292 ( .I1(n274), .I2(n23), .O(n273) );
  OR_GATE U293 ( .I1(n23), .I2(n274), .O(n271) );
  AND_GATE U294 ( .I1(n275), .I2(n276), .O(n270) );
  NAND_GATE U295 ( .I1(B[11]), .I2(n22), .O(n276) );
  OR_GATE U296 ( .I1(n22), .I2(B[11]), .O(n275) );
  AND_GATE U297 ( .I1(n277), .I2(n278), .O(SUM[10]) );
  NAND_GATE U298 ( .I1(n279), .I2(n274), .O(n278) );
  OR_GATE U299 ( .I1(n279), .I2(n274), .O(n277) );
  AND_GATE U300 ( .I1(n280), .I2(n281), .O(n274) );
  NAND_GATE U301 ( .I1(B[9]), .I2(n282), .O(n281) );
  NAND_GATE U302 ( .I1(n36), .I2(n24), .O(n282) );
  OR_GATE U303 ( .I1(n24), .I2(n36), .O(n280) );
  AND_GATE U304 ( .I1(n283), .I2(n284), .O(n36) );
  NAND_GATE U305 ( .I1(B[8]), .I2(n285), .O(n284) );
  NAND_GATE U306 ( .I1(n42), .I2(n25), .O(n285) );
  OR_GATE U307 ( .I1(n25), .I2(n42), .O(n283) );
  AND_GATE U308 ( .I1(n286), .I2(n287), .O(n42) );
  NAND_GATE U309 ( .I1(B[7]), .I2(n288), .O(n287) );
  NAND_GATE U310 ( .I1(n48), .I2(n26), .O(n288) );
  OR_GATE U311 ( .I1(n26), .I2(n48), .O(n286) );
  AND_GATE U312 ( .I1(n289), .I2(n290), .O(n48) );
  NAND_GATE U313 ( .I1(B[6]), .I2(n291), .O(n290) );
  NAND_GATE U314 ( .I1(n54), .I2(n27), .O(n291) );
  OR_GATE U315 ( .I1(n27), .I2(n54), .O(n289) );
  AND_GATE U316 ( .I1(n292), .I2(n293), .O(n54) );
  NAND_GATE U317 ( .I1(B[5]), .I2(n294), .O(n293) );
  NAND_GATE U318 ( .I1(n60), .I2(n28), .O(n294) );
  OR_GATE U319 ( .I1(n28), .I2(n60), .O(n292) );
  AND_GATE U320 ( .I1(n295), .I2(n296), .O(n60) );
  NAND_GATE U321 ( .I1(B[4]), .I2(n297), .O(n296) );
  NAND_GATE U322 ( .I1(n66), .I2(n29), .O(n297) );
  OR_GATE U323 ( .I1(n29), .I2(n66), .O(n295) );
  AND_GATE U324 ( .I1(n298), .I2(n299), .O(n66) );
  NAND_GATE U325 ( .I1(B[3]), .I2(n300), .O(n299) );
  NAND_GATE U326 ( .I1(n72), .I2(n30), .O(n300) );
  OR_GATE U327 ( .I1(n30), .I2(n72), .O(n298) );
  AND_GATE U328 ( .I1(n301), .I2(n302), .O(n72) );
  NAND_GATE U329 ( .I1(B[2]), .I2(n303), .O(n302) );
  NAND_GATE U330 ( .I1(n97), .I2(n31), .O(n303) );
  OR_GATE U331 ( .I1(n31), .I2(n97), .O(n301) );
  AND_GATE U332 ( .I1(n304), .I2(n305), .O(n97) );
  NAND_GATE U333 ( .I1(B[1]), .I2(n306), .O(n305) );
  OR_GATE U334 ( .I1(A[1]), .I2(n193), .O(n306) );
  NAND_GATE U335 ( .I1(A[1]), .I2(n193), .O(n304) );
  AND_GATE U336 ( .I1(B[0]), .I2(A[0]), .O(n193) );
  AND_GATE U337 ( .I1(n307), .I2(n308), .O(n279) );
  NAND_GATE U338 ( .I1(B[10]), .I2(n23), .O(n308) );
  OR_GATE U339 ( .I1(n23), .I2(B[10]), .O(n307) );
  NAND_GATE U340 ( .I1(n309), .I2(n310), .O(SUM[0]) );
  OR_GATE U341 ( .I1(n1), .I2(A[0]), .O(n310) );
  NAND_GATE U342 ( .I1(A[0]), .I2(n1), .O(n309) );
endmodule


module predict_nb_record3_1_DW01_cmp6_9 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[0]), .O(n2) );
  INV_GATE U3 ( .I1(A[2]), .O(n3) );
  INV_GATE U4 ( .I1(A[3]), .O(n4) );
  INV_GATE U5 ( .I1(A[4]), .O(n5) );
  INV_GATE U6 ( .I1(A[5]), .O(n6) );
  INV_GATE U7 ( .I1(A[6]), .O(n7) );
  INV_GATE U8 ( .I1(A[7]), .O(n8) );
  INV_GATE U9 ( .I1(A[8]), .O(n9) );
  INV_GATE U10 ( .I1(A[9]), .O(n10) );
  INV_GATE U11 ( .I1(A[10]), .O(n11) );
  INV_GATE U12 ( .I1(A[11]), .O(n12) );
  INV_GATE U13 ( .I1(A[12]), .O(n13) );
  INV_GATE U14 ( .I1(A[13]), .O(n14) );
  INV_GATE U15 ( .I1(A[14]), .O(n15) );
  INV_GATE U16 ( .I1(A[15]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[17]), .O(n18) );
  INV_GATE U19 ( .I1(A[18]), .O(n19) );
  INV_GATE U20 ( .I1(A[19]), .O(n20) );
  INV_GATE U21 ( .I1(A[20]), .O(n21) );
  INV_GATE U22 ( .I1(A[21]), .O(n22) );
  INV_GATE U23 ( .I1(A[22]), .O(n23) );
  INV_GATE U24 ( .I1(A[23]), .O(n24) );
  INV_GATE U25 ( .I1(A[24]), .O(n25) );
  INV_GATE U26 ( .I1(A[25]), .O(n26) );
  INV_GATE U27 ( .I1(A[26]), .O(n27) );
  INV_GATE U28 ( .I1(A[27]), .O(n28) );
  INV_GATE U29 ( .I1(A[28]), .O(n29) );
  INV_GATE U30 ( .I1(A[29]), .O(n30) );
  INV_GATE U31 ( .I1(A[30]), .O(n31) );
  INV_GATE U32 ( .I1(A[31]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n16), .O(n49) );
  OR_GATE U38 ( .I1(n16), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n18), .O(n44) );
  OR_GATE U42 ( .I1(n18), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n19), .O(n42) );
  OR_GATE U44 ( .I1(n19), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n20), .O(n58) );
  OR_GATE U48 ( .I1(n20), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n21), .O(n56) );
  OR_GATE U50 ( .I1(n21), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n22), .O(n53) );
  OR_GATE U52 ( .I1(n22), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n23), .O(n51) );
  OR_GATE U54 ( .I1(n23), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n24), .O(n67) );
  OR_GATE U58 ( .I1(n24), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n25), .O(n65) );
  OR_GATE U60 ( .I1(n25), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n26), .O(n62) );
  OR_GATE U62 ( .I1(n26), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n27), .O(n60) );
  OR_GATE U64 ( .I1(n27), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n28), .O(n76) );
  OR_GATE U68 ( .I1(n28), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n29), .O(n74) );
  OR_GATE U70 ( .I1(n29), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n30), .O(n71) );
  OR_GATE U72 ( .I1(n30), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n31), .O(n69) );
  OR_GATE U74 ( .I1(n31), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n4), .O(n85) );
  OR_GATE U78 ( .I1(n4), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n5), .O(n83) );
  OR_GATE U80 ( .I1(n5), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n6), .O(n89) );
  OR_GATE U83 ( .I1(n6), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n7), .O(n87) );
  OR_GATE U85 ( .I1(n7), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n32), .O(n93) );
  OR_GATE U88 ( .I1(n32), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n3), .O(n91) );
  OR_GATE U90 ( .I1(n3), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n2), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n2), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n8), .O(n108) );
  OR_GATE U102 ( .I1(n8), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n9), .O(n106) );
  OR_GATE U104 ( .I1(n9), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n10), .O(n103) );
  OR_GATE U106 ( .I1(n10), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n11), .O(n101) );
  OR_GATE U108 ( .I1(n11), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n12), .O(n117) );
  OR_GATE U112 ( .I1(n12), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n13), .O(n115) );
  OR_GATE U114 ( .I1(n13), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n14), .O(n112) );
  OR_GATE U116 ( .I1(n14), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n15), .O(n110) );
  OR_GATE U118 ( .I1(n15), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_8 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[0]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n18), .O(n49) );
  OR_GATE U38 ( .I1(n18), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n16), .O(n44) );
  OR_GATE U42 ( .I1(n16), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n15), .O(n42) );
  OR_GATE U44 ( .I1(n15), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n14), .O(n58) );
  OR_GATE U48 ( .I1(n14), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n13), .O(n56) );
  OR_GATE U50 ( .I1(n13), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n12), .O(n53) );
  OR_GATE U52 ( .I1(n12), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n11), .O(n51) );
  OR_GATE U54 ( .I1(n11), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n10), .O(n67) );
  OR_GATE U58 ( .I1(n10), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n9), .O(n65) );
  OR_GATE U60 ( .I1(n9), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n8), .O(n62) );
  OR_GATE U62 ( .I1(n8), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n7), .O(n60) );
  OR_GATE U64 ( .I1(n7), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n6), .O(n76) );
  OR_GATE U68 ( .I1(n6), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n5), .O(n74) );
  OR_GATE U70 ( .I1(n5), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n4), .O(n71) );
  OR_GATE U72 ( .I1(n4), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n3), .O(n69) );
  OR_GATE U74 ( .I1(n3), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n30), .O(n85) );
  OR_GATE U78 ( .I1(n30), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n29), .O(n83) );
  OR_GATE U80 ( .I1(n29), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n28), .O(n89) );
  OR_GATE U83 ( .I1(n28), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n27), .O(n87) );
  OR_GATE U85 ( .I1(n27), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n31), .O(n91) );
  OR_GATE U90 ( .I1(n31), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n26), .O(n108) );
  OR_GATE U102 ( .I1(n26), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n25), .O(n106) );
  OR_GATE U104 ( .I1(n25), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n24), .O(n103) );
  OR_GATE U106 ( .I1(n24), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n23), .O(n101) );
  OR_GATE U108 ( .I1(n23), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n22), .O(n117) );
  OR_GATE U112 ( .I1(n22), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n21), .O(n115) );
  OR_GATE U114 ( .I1(n21), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n20), .O(n112) );
  OR_GATE U116 ( .I1(n20), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n19), .O(n110) );
  OR_GATE U118 ( .I1(n19), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_7 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[0]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n18), .O(n49) );
  OR_GATE U38 ( .I1(n18), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n16), .O(n44) );
  OR_GATE U42 ( .I1(n16), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n15), .O(n42) );
  OR_GATE U44 ( .I1(n15), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n14), .O(n58) );
  OR_GATE U48 ( .I1(n14), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n13), .O(n56) );
  OR_GATE U50 ( .I1(n13), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n12), .O(n53) );
  OR_GATE U52 ( .I1(n12), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n11), .O(n51) );
  OR_GATE U54 ( .I1(n11), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n10), .O(n67) );
  OR_GATE U58 ( .I1(n10), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n9), .O(n65) );
  OR_GATE U60 ( .I1(n9), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n8), .O(n62) );
  OR_GATE U62 ( .I1(n8), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n7), .O(n60) );
  OR_GATE U64 ( .I1(n7), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n6), .O(n76) );
  OR_GATE U68 ( .I1(n6), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n5), .O(n74) );
  OR_GATE U70 ( .I1(n5), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n4), .O(n71) );
  OR_GATE U72 ( .I1(n4), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n3), .O(n69) );
  OR_GATE U74 ( .I1(n3), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n30), .O(n85) );
  OR_GATE U78 ( .I1(n30), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n29), .O(n83) );
  OR_GATE U80 ( .I1(n29), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n28), .O(n89) );
  OR_GATE U83 ( .I1(n28), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n27), .O(n87) );
  OR_GATE U85 ( .I1(n27), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n31), .O(n91) );
  OR_GATE U90 ( .I1(n31), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n26), .O(n108) );
  OR_GATE U102 ( .I1(n26), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n25), .O(n106) );
  OR_GATE U104 ( .I1(n25), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n24), .O(n103) );
  OR_GATE U106 ( .I1(n24), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n23), .O(n101) );
  OR_GATE U108 ( .I1(n23), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n22), .O(n117) );
  OR_GATE U112 ( .I1(n22), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n21), .O(n115) );
  OR_GATE U114 ( .I1(n21), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n20), .O(n112) );
  OR_GATE U116 ( .I1(n20), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n19), .O(n110) );
  OR_GATE U118 ( .I1(n19), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_6 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[0]), .O(n2) );
  INV_GATE U3 ( .I1(A[2]), .O(n3) );
  INV_GATE U4 ( .I1(A[3]), .O(n4) );
  INV_GATE U5 ( .I1(A[4]), .O(n5) );
  INV_GATE U6 ( .I1(A[5]), .O(n6) );
  INV_GATE U7 ( .I1(A[6]), .O(n7) );
  INV_GATE U8 ( .I1(A[7]), .O(n8) );
  INV_GATE U9 ( .I1(A[8]), .O(n9) );
  INV_GATE U10 ( .I1(A[9]), .O(n10) );
  INV_GATE U11 ( .I1(A[10]), .O(n11) );
  INV_GATE U12 ( .I1(A[11]), .O(n12) );
  INV_GATE U13 ( .I1(A[12]), .O(n13) );
  INV_GATE U14 ( .I1(A[13]), .O(n14) );
  INV_GATE U15 ( .I1(A[14]), .O(n15) );
  INV_GATE U16 ( .I1(A[15]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[17]), .O(n18) );
  INV_GATE U19 ( .I1(A[18]), .O(n19) );
  INV_GATE U20 ( .I1(A[19]), .O(n20) );
  INV_GATE U21 ( .I1(A[20]), .O(n21) );
  INV_GATE U22 ( .I1(A[21]), .O(n22) );
  INV_GATE U23 ( .I1(A[22]), .O(n23) );
  INV_GATE U24 ( .I1(A[23]), .O(n24) );
  INV_GATE U25 ( .I1(A[24]), .O(n25) );
  INV_GATE U26 ( .I1(A[25]), .O(n26) );
  INV_GATE U27 ( .I1(A[26]), .O(n27) );
  INV_GATE U28 ( .I1(A[27]), .O(n28) );
  INV_GATE U29 ( .I1(A[28]), .O(n29) );
  INV_GATE U30 ( .I1(A[29]), .O(n30) );
  INV_GATE U31 ( .I1(A[30]), .O(n31) );
  INV_GATE U32 ( .I1(A[31]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n16), .O(n49) );
  OR_GATE U38 ( .I1(n16), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n18), .O(n44) );
  OR_GATE U42 ( .I1(n18), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n19), .O(n42) );
  OR_GATE U44 ( .I1(n19), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n20), .O(n58) );
  OR_GATE U48 ( .I1(n20), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n21), .O(n56) );
  OR_GATE U50 ( .I1(n21), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n22), .O(n53) );
  OR_GATE U52 ( .I1(n22), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n23), .O(n51) );
  OR_GATE U54 ( .I1(n23), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n24), .O(n67) );
  OR_GATE U58 ( .I1(n24), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n25), .O(n65) );
  OR_GATE U60 ( .I1(n25), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n26), .O(n62) );
  OR_GATE U62 ( .I1(n26), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n27), .O(n60) );
  OR_GATE U64 ( .I1(n27), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n28), .O(n76) );
  OR_GATE U68 ( .I1(n28), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n29), .O(n74) );
  OR_GATE U70 ( .I1(n29), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n30), .O(n71) );
  OR_GATE U72 ( .I1(n30), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n31), .O(n69) );
  OR_GATE U74 ( .I1(n31), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n4), .O(n85) );
  OR_GATE U78 ( .I1(n4), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n5), .O(n83) );
  OR_GATE U80 ( .I1(n5), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n6), .O(n89) );
  OR_GATE U83 ( .I1(n6), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n7), .O(n87) );
  OR_GATE U85 ( .I1(n7), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n32), .O(n93) );
  OR_GATE U88 ( .I1(n32), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n3), .O(n91) );
  OR_GATE U90 ( .I1(n3), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n2), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n2), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n8), .O(n108) );
  OR_GATE U102 ( .I1(n8), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n9), .O(n106) );
  OR_GATE U104 ( .I1(n9), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n10), .O(n103) );
  OR_GATE U106 ( .I1(n10), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n11), .O(n101) );
  OR_GATE U108 ( .I1(n11), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n12), .O(n117) );
  OR_GATE U112 ( .I1(n12), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n13), .O(n115) );
  OR_GATE U114 ( .I1(n13), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n14), .O(n112) );
  OR_GATE U116 ( .I1(n14), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n15), .O(n110) );
  OR_GATE U118 ( .I1(n15), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_5 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[0]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n18), .O(n49) );
  OR_GATE U38 ( .I1(n18), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n16), .O(n44) );
  OR_GATE U42 ( .I1(n16), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n15), .O(n42) );
  OR_GATE U44 ( .I1(n15), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n14), .O(n58) );
  OR_GATE U48 ( .I1(n14), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n13), .O(n56) );
  OR_GATE U50 ( .I1(n13), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n12), .O(n53) );
  OR_GATE U52 ( .I1(n12), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n11), .O(n51) );
  OR_GATE U54 ( .I1(n11), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n10), .O(n67) );
  OR_GATE U58 ( .I1(n10), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n9), .O(n65) );
  OR_GATE U60 ( .I1(n9), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n8), .O(n62) );
  OR_GATE U62 ( .I1(n8), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n7), .O(n60) );
  OR_GATE U64 ( .I1(n7), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n6), .O(n76) );
  OR_GATE U68 ( .I1(n6), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n5), .O(n74) );
  OR_GATE U70 ( .I1(n5), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n4), .O(n71) );
  OR_GATE U72 ( .I1(n4), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n3), .O(n69) );
  OR_GATE U74 ( .I1(n3), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n30), .O(n85) );
  OR_GATE U78 ( .I1(n30), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n29), .O(n83) );
  OR_GATE U80 ( .I1(n29), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n28), .O(n89) );
  OR_GATE U83 ( .I1(n28), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n27), .O(n87) );
  OR_GATE U85 ( .I1(n27), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n31), .O(n91) );
  OR_GATE U90 ( .I1(n31), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n26), .O(n108) );
  OR_GATE U102 ( .I1(n26), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n25), .O(n106) );
  OR_GATE U104 ( .I1(n25), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n24), .O(n103) );
  OR_GATE U106 ( .I1(n24), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n23), .O(n101) );
  OR_GATE U108 ( .I1(n23), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n22), .O(n117) );
  OR_GATE U112 ( .I1(n22), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n21), .O(n115) );
  OR_GATE U114 ( .I1(n21), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n20), .O(n112) );
  OR_GATE U116 ( .I1(n20), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n19), .O(n110) );
  OR_GATE U118 ( .I1(n19), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_4 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[0]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n18), .O(n49) );
  OR_GATE U38 ( .I1(n18), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n16), .O(n44) );
  OR_GATE U42 ( .I1(n16), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n15), .O(n42) );
  OR_GATE U44 ( .I1(n15), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n14), .O(n58) );
  OR_GATE U48 ( .I1(n14), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n13), .O(n56) );
  OR_GATE U50 ( .I1(n13), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n12), .O(n53) );
  OR_GATE U52 ( .I1(n12), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n11), .O(n51) );
  OR_GATE U54 ( .I1(n11), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n10), .O(n67) );
  OR_GATE U58 ( .I1(n10), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n9), .O(n65) );
  OR_GATE U60 ( .I1(n9), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n8), .O(n62) );
  OR_GATE U62 ( .I1(n8), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n7), .O(n60) );
  OR_GATE U64 ( .I1(n7), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n6), .O(n76) );
  OR_GATE U68 ( .I1(n6), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n5), .O(n74) );
  OR_GATE U70 ( .I1(n5), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n4), .O(n71) );
  OR_GATE U72 ( .I1(n4), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n3), .O(n69) );
  OR_GATE U74 ( .I1(n3), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n30), .O(n85) );
  OR_GATE U78 ( .I1(n30), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n29), .O(n83) );
  OR_GATE U80 ( .I1(n29), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n28), .O(n89) );
  OR_GATE U83 ( .I1(n28), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n27), .O(n87) );
  OR_GATE U85 ( .I1(n27), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n31), .O(n91) );
  OR_GATE U90 ( .I1(n31), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n26), .O(n108) );
  OR_GATE U102 ( .I1(n26), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n25), .O(n106) );
  OR_GATE U104 ( .I1(n25), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n24), .O(n103) );
  OR_GATE U106 ( .I1(n24), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n23), .O(n101) );
  OR_GATE U108 ( .I1(n23), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n22), .O(n117) );
  OR_GATE U112 ( .I1(n22), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n21), .O(n115) );
  OR_GATE U114 ( .I1(n21), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n20), .O(n112) );
  OR_GATE U116 ( .I1(n20), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n19), .O(n110) );
  OR_GATE U118 ( .I1(n19), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_3 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[0]), .O(n2) );
  INV_GATE U3 ( .I1(A[2]), .O(n3) );
  INV_GATE U4 ( .I1(A[3]), .O(n4) );
  INV_GATE U5 ( .I1(A[4]), .O(n5) );
  INV_GATE U6 ( .I1(A[5]), .O(n6) );
  INV_GATE U7 ( .I1(A[6]), .O(n7) );
  INV_GATE U8 ( .I1(A[7]), .O(n8) );
  INV_GATE U9 ( .I1(A[8]), .O(n9) );
  INV_GATE U10 ( .I1(A[9]), .O(n10) );
  INV_GATE U11 ( .I1(A[10]), .O(n11) );
  INV_GATE U12 ( .I1(A[11]), .O(n12) );
  INV_GATE U13 ( .I1(A[12]), .O(n13) );
  INV_GATE U14 ( .I1(A[13]), .O(n14) );
  INV_GATE U15 ( .I1(A[14]), .O(n15) );
  INV_GATE U16 ( .I1(A[15]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[17]), .O(n18) );
  INV_GATE U19 ( .I1(A[18]), .O(n19) );
  INV_GATE U20 ( .I1(A[19]), .O(n20) );
  INV_GATE U21 ( .I1(A[20]), .O(n21) );
  INV_GATE U22 ( .I1(A[21]), .O(n22) );
  INV_GATE U23 ( .I1(A[22]), .O(n23) );
  INV_GATE U24 ( .I1(A[23]), .O(n24) );
  INV_GATE U25 ( .I1(A[24]), .O(n25) );
  INV_GATE U26 ( .I1(A[25]), .O(n26) );
  INV_GATE U27 ( .I1(A[26]), .O(n27) );
  INV_GATE U28 ( .I1(A[27]), .O(n28) );
  INV_GATE U29 ( .I1(A[28]), .O(n29) );
  INV_GATE U30 ( .I1(A[29]), .O(n30) );
  INV_GATE U31 ( .I1(A[30]), .O(n31) );
  INV_GATE U32 ( .I1(A[31]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n16), .O(n49) );
  OR_GATE U38 ( .I1(n16), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n18), .O(n44) );
  OR_GATE U42 ( .I1(n18), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n19), .O(n42) );
  OR_GATE U44 ( .I1(n19), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n20), .O(n58) );
  OR_GATE U48 ( .I1(n20), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n21), .O(n56) );
  OR_GATE U50 ( .I1(n21), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n22), .O(n53) );
  OR_GATE U52 ( .I1(n22), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n23), .O(n51) );
  OR_GATE U54 ( .I1(n23), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n24), .O(n67) );
  OR_GATE U58 ( .I1(n24), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n25), .O(n65) );
  OR_GATE U60 ( .I1(n25), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n26), .O(n62) );
  OR_GATE U62 ( .I1(n26), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n27), .O(n60) );
  OR_GATE U64 ( .I1(n27), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n28), .O(n76) );
  OR_GATE U68 ( .I1(n28), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n29), .O(n74) );
  OR_GATE U70 ( .I1(n29), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n30), .O(n71) );
  OR_GATE U72 ( .I1(n30), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n31), .O(n69) );
  OR_GATE U74 ( .I1(n31), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n4), .O(n85) );
  OR_GATE U78 ( .I1(n4), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n5), .O(n83) );
  OR_GATE U80 ( .I1(n5), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n6), .O(n89) );
  OR_GATE U83 ( .I1(n6), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n7), .O(n87) );
  OR_GATE U85 ( .I1(n7), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n32), .O(n93) );
  OR_GATE U88 ( .I1(n32), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n3), .O(n91) );
  OR_GATE U90 ( .I1(n3), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n2), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n2), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n8), .O(n108) );
  OR_GATE U102 ( .I1(n8), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n9), .O(n106) );
  OR_GATE U104 ( .I1(n9), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n10), .O(n103) );
  OR_GATE U106 ( .I1(n10), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n11), .O(n101) );
  OR_GATE U108 ( .I1(n11), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n12), .O(n117) );
  OR_GATE U112 ( .I1(n12), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n13), .O(n115) );
  OR_GATE U114 ( .I1(n13), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n14), .O(n112) );
  OR_GATE U116 ( .I1(n14), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n15), .O(n110) );
  OR_GATE U118 ( .I1(n15), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_2 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[0]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n18), .O(n49) );
  OR_GATE U38 ( .I1(n18), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n16), .O(n44) );
  OR_GATE U42 ( .I1(n16), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n15), .O(n42) );
  OR_GATE U44 ( .I1(n15), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n14), .O(n58) );
  OR_GATE U48 ( .I1(n14), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n13), .O(n56) );
  OR_GATE U50 ( .I1(n13), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n12), .O(n53) );
  OR_GATE U52 ( .I1(n12), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n11), .O(n51) );
  OR_GATE U54 ( .I1(n11), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n10), .O(n67) );
  OR_GATE U58 ( .I1(n10), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n9), .O(n65) );
  OR_GATE U60 ( .I1(n9), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n8), .O(n62) );
  OR_GATE U62 ( .I1(n8), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n7), .O(n60) );
  OR_GATE U64 ( .I1(n7), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n6), .O(n76) );
  OR_GATE U68 ( .I1(n6), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n5), .O(n74) );
  OR_GATE U70 ( .I1(n5), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n4), .O(n71) );
  OR_GATE U72 ( .I1(n4), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n3), .O(n69) );
  OR_GATE U74 ( .I1(n3), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n30), .O(n85) );
  OR_GATE U78 ( .I1(n30), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n29), .O(n83) );
  OR_GATE U80 ( .I1(n29), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n28), .O(n89) );
  OR_GATE U83 ( .I1(n28), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n27), .O(n87) );
  OR_GATE U85 ( .I1(n27), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n31), .O(n91) );
  OR_GATE U90 ( .I1(n31), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n26), .O(n108) );
  OR_GATE U102 ( .I1(n26), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n25), .O(n106) );
  OR_GATE U104 ( .I1(n25), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n24), .O(n103) );
  OR_GATE U106 ( .I1(n24), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n23), .O(n101) );
  OR_GATE U108 ( .I1(n23), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n22), .O(n117) );
  OR_GATE U112 ( .I1(n22), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n21), .O(n115) );
  OR_GATE U114 ( .I1(n21), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n20), .O(n112) );
  OR_GATE U116 ( .I1(n20), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n19), .O(n110) );
  OR_GATE U118 ( .I1(n19), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(B[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[31]), .O(n2) );
  INV_GATE U3 ( .I1(A[30]), .O(n3) );
  INV_GATE U4 ( .I1(A[29]), .O(n4) );
  INV_GATE U5 ( .I1(A[28]), .O(n5) );
  INV_GATE U6 ( .I1(A[27]), .O(n6) );
  INV_GATE U7 ( .I1(A[26]), .O(n7) );
  INV_GATE U8 ( .I1(A[25]), .O(n8) );
  INV_GATE U9 ( .I1(A[24]), .O(n9) );
  INV_GATE U10 ( .I1(A[23]), .O(n10) );
  INV_GATE U11 ( .I1(A[22]), .O(n11) );
  INV_GATE U12 ( .I1(A[21]), .O(n12) );
  INV_GATE U13 ( .I1(A[20]), .O(n13) );
  INV_GATE U14 ( .I1(A[19]), .O(n14) );
  INV_GATE U15 ( .I1(A[18]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[16]), .O(n17) );
  INV_GATE U18 ( .I1(A[15]), .O(n18) );
  INV_GATE U19 ( .I1(A[14]), .O(n19) );
  INV_GATE U20 ( .I1(A[13]), .O(n20) );
  INV_GATE U21 ( .I1(A[12]), .O(n21) );
  INV_GATE U22 ( .I1(A[11]), .O(n22) );
  INV_GATE U23 ( .I1(A[10]), .O(n23) );
  INV_GATE U24 ( .I1(A[9]), .O(n24) );
  INV_GATE U25 ( .I1(A[8]), .O(n25) );
  INV_GATE U26 ( .I1(A[7]), .O(n26) );
  INV_GATE U27 ( .I1(A[6]), .O(n27) );
  INV_GATE U28 ( .I1(A[5]), .O(n28) );
  INV_GATE U29 ( .I1(A[4]), .O(n29) );
  INV_GATE U30 ( .I1(A[3]), .O(n30) );
  INV_GATE U31 ( .I1(A[2]), .O(n31) );
  INV_GATE U32 ( .I1(A[0]), .O(n32) );
  AND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(EQ) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[15]), .I2(n18), .O(n49) );
  OR_GATE U38 ( .I1(n18), .I2(B[15]), .O(n48) );
  NAND_GATE U39 ( .I1(B[16]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[16]), .O(n46) );
  NAND_GATE U41 ( .I1(B[17]), .I2(n16), .O(n44) );
  OR_GATE U42 ( .I1(n16), .I2(B[17]), .O(n43) );
  NAND_GATE U43 ( .I1(B[18]), .I2(n15), .O(n42) );
  OR_GATE U44 ( .I1(n15), .I2(B[18]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[19]), .I2(n14), .O(n58) );
  OR_GATE U48 ( .I1(n14), .I2(B[19]), .O(n57) );
  NAND_GATE U49 ( .I1(B[20]), .I2(n13), .O(n56) );
  OR_GATE U50 ( .I1(n13), .I2(B[20]), .O(n55) );
  NAND_GATE U51 ( .I1(B[21]), .I2(n12), .O(n53) );
  OR_GATE U52 ( .I1(n12), .I2(B[21]), .O(n52) );
  NAND_GATE U53 ( .I1(B[22]), .I2(n11), .O(n51) );
  OR_GATE U54 ( .I1(n11), .I2(B[22]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[23]), .I2(n10), .O(n67) );
  OR_GATE U58 ( .I1(n10), .I2(B[23]), .O(n66) );
  NAND_GATE U59 ( .I1(B[24]), .I2(n9), .O(n65) );
  OR_GATE U60 ( .I1(n9), .I2(B[24]), .O(n64) );
  NAND_GATE U61 ( .I1(B[25]), .I2(n8), .O(n62) );
  OR_GATE U62 ( .I1(n8), .I2(B[25]), .O(n61) );
  NAND_GATE U63 ( .I1(B[26]), .I2(n7), .O(n60) );
  OR_GATE U64 ( .I1(n7), .I2(B[26]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[27]), .I2(n6), .O(n76) );
  OR_GATE U68 ( .I1(n6), .I2(B[27]), .O(n75) );
  NAND_GATE U69 ( .I1(B[28]), .I2(n5), .O(n74) );
  OR_GATE U70 ( .I1(n5), .I2(B[28]), .O(n73) );
  NAND_GATE U71 ( .I1(B[29]), .I2(n4), .O(n71) );
  OR_GATE U72 ( .I1(n4), .I2(B[29]), .O(n70) );
  NAND_GATE U73 ( .I1(B[30]), .I2(n3), .O(n69) );
  OR_GATE U74 ( .I1(n3), .I2(B[30]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[3]), .I2(n30), .O(n85) );
  OR_GATE U78 ( .I1(n30), .I2(B[3]), .O(n84) );
  NAND_GATE U79 ( .I1(B[4]), .I2(n29), .O(n83) );
  OR_GATE U80 ( .I1(n29), .I2(B[4]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[5]), .I2(n28), .O(n89) );
  OR_GATE U83 ( .I1(n28), .I2(B[5]), .O(n88) );
  NAND_GATE U84 ( .I1(B[6]), .I2(n27), .O(n87) );
  OR_GATE U85 ( .I1(n27), .I2(B[6]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[31]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[31]), .O(n92) );
  NAND_GATE U89 ( .I1(B[2]), .I2(n31), .O(n91) );
  OR_GATE U90 ( .I1(n31), .I2(B[2]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(n96), .I2(n1), .O(n95) );
  NAND_GATE U93 ( .I1(A[1]), .I2(n96), .O(n94) );
  NAND_GATE U94 ( .I1(B[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n1), .I2(n99), .O(n98) );
  OR_GATE U97 ( .I1(n99), .I2(A[1]), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(B[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[7]), .I2(n26), .O(n108) );
  OR_GATE U102 ( .I1(n26), .I2(B[7]), .O(n107) );
  NAND_GATE U103 ( .I1(B[8]), .I2(n25), .O(n106) );
  OR_GATE U104 ( .I1(n25), .I2(B[8]), .O(n105) );
  NAND_GATE U105 ( .I1(B[9]), .I2(n24), .O(n103) );
  OR_GATE U106 ( .I1(n24), .I2(B[9]), .O(n102) );
  NAND_GATE U107 ( .I1(B[10]), .I2(n23), .O(n101) );
  OR_GATE U108 ( .I1(n23), .I2(B[10]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[11]), .I2(n22), .O(n117) );
  OR_GATE U112 ( .I1(n22), .I2(B[11]), .O(n116) );
  NAND_GATE U113 ( .I1(B[12]), .I2(n21), .O(n115) );
  OR_GATE U114 ( .I1(n21), .I2(B[12]), .O(n114) );
  NAND_GATE U115 ( .I1(B[13]), .I2(n20), .O(n112) );
  OR_GATE U116 ( .I1(n20), .I2(B[13]), .O(n111) );
  NAND_GATE U117 ( .I1(B[14]), .I2(n19), .O(n110) );
  OR_GATE U118 ( .I1(n19), .I2(B[14]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_GATE U1 ( .I1(A[2]), .O(SUM[2]) );
  INV_GATE U2 ( .I1(n112), .O(n2) );
  INV_GATE U3 ( .I1(n32), .O(n3) );
  INV_GATE U4 ( .I1(A[3]), .O(n4) );
  INV_GATE U5 ( .I1(A[4]), .O(n5) );
  INV_GATE U6 ( .I1(A[5]), .O(n6) );
  INV_GATE U7 ( .I1(A[6]), .O(n7) );
  INV_GATE U8 ( .I1(A[7]), .O(n8) );
  INV_GATE U9 ( .I1(A[8]), .O(n9) );
  INV_GATE U10 ( .I1(A[11]), .O(n10) );
  INV_GATE U11 ( .I1(A[12]), .O(n11) );
  INV_GATE U12 ( .I1(A[13]), .O(n12) );
  INV_GATE U13 ( .I1(A[14]), .O(n13) );
  INV_GATE U14 ( .I1(A[15]), .O(n14) );
  INV_GATE U15 ( .I1(A[16]), .O(n15) );
  INV_GATE U16 ( .I1(A[17]), .O(n16) );
  INV_GATE U17 ( .I1(A[18]), .O(n17) );
  INV_GATE U18 ( .I1(A[19]), .O(n18) );
  INV_GATE U19 ( .I1(A[20]), .O(n19) );
  INV_GATE U20 ( .I1(A[21]), .O(n20) );
  INV_GATE U21 ( .I1(A[22]), .O(n21) );
  INV_GATE U22 ( .I1(A[23]), .O(n22) );
  INV_GATE U23 ( .I1(A[24]), .O(n23) );
  INV_GATE U24 ( .I1(A[25]), .O(n24) );
  INV_GATE U25 ( .I1(A[26]), .O(n25) );
  INV_GATE U26 ( .I1(A[27]), .O(n26) );
  INV_GATE U27 ( .I1(A[28]), .O(n27) );
  INV_GATE U28 ( .I1(A[29]), .O(n28) );
  INV_GATE U29 ( .I1(A[30]), .O(n29) );
  NAND_GATE U30 ( .I1(n30), .I2(n31), .O(SUM[9]) );
  NAND_GATE U31 ( .I1(A[9]), .I2(n3), .O(n31) );
  OR_GATE U32 ( .I1(n3), .I2(A[9]), .O(n30) );
  NAND_GATE U33 ( .I1(n33), .I2(n34), .O(SUM[8]) );
  OR_GATE U34 ( .I1(n9), .I2(n35), .O(n34) );
  NAND_GATE U35 ( .I1(n35), .I2(n9), .O(n33) );
  AND_GATE U36 ( .I1(A[7]), .I2(n36), .O(n35) );
  NAND_GATE U37 ( .I1(n37), .I2(n38), .O(SUM[7]) );
  OR_GATE U38 ( .I1(n8), .I2(n36), .O(n38) );
  NAND_GATE U39 ( .I1(n36), .I2(n8), .O(n37) );
  NAND_GATE U40 ( .I1(n39), .I2(n40), .O(SUM[6]) );
  OR_GATE U41 ( .I1(n7), .I2(n41), .O(n40) );
  NAND_GATE U42 ( .I1(n41), .I2(n7), .O(n39) );
  AND_GATE U43 ( .I1(A[5]), .I2(n42), .O(n41) );
  NAND_GATE U44 ( .I1(n43), .I2(n44), .O(SUM[5]) );
  OR_GATE U45 ( .I1(n6), .I2(n42), .O(n44) );
  NAND_GATE U46 ( .I1(n42), .I2(n6), .O(n43) );
  NAND_GATE U47 ( .I1(n45), .I2(n46), .O(SUM[4]) );
  OR_GATE U48 ( .I1(n5), .I2(n47), .O(n46) );
  NAND_GATE U49 ( .I1(n47), .I2(n5), .O(n45) );
  AND_GATE U50 ( .I1(A[3]), .I2(A[2]), .O(n47) );
  NAND_GATE U51 ( .I1(n48), .I2(n49), .O(SUM[3]) );
  NAND_GATE U52 ( .I1(A[3]), .I2(SUM[2]), .O(n49) );
  NAND_GATE U53 ( .I1(A[2]), .I2(n4), .O(n48) );
  NAND_GATE U54 ( .I1(n50), .I2(n51), .O(SUM[31]) );
  NAND_GATE U55 ( .I1(A[31]), .I2(n52), .O(n51) );
  OR_GATE U56 ( .I1(n52), .I2(A[31]), .O(n50) );
  NAND_GATE U57 ( .I1(A[30]), .I2(n53), .O(n52) );
  NAND_GATE U58 ( .I1(n54), .I2(n55), .O(SUM[30]) );
  OR_GATE U59 ( .I1(n29), .I2(n53), .O(n55) );
  NAND_GATE U60 ( .I1(n53), .I2(n29), .O(n54) );
  AND_GATE U61 ( .I1(A[29]), .I2(n56), .O(n53) );
  NAND_GATE U62 ( .I1(n57), .I2(n58), .O(SUM[29]) );
  OR_GATE U63 ( .I1(n28), .I2(n56), .O(n58) );
  NAND_GATE U64 ( .I1(n56), .I2(n28), .O(n57) );
  AND3_GATE U65 ( .I1(A[27]), .I2(n59), .I3(A[28]), .O(n56) );
  NAND_GATE U66 ( .I1(n60), .I2(n61), .O(SUM[28]) );
  OR_GATE U67 ( .I1(n27), .I2(n62), .O(n61) );
  NAND_GATE U68 ( .I1(n62), .I2(n27), .O(n60) );
  AND_GATE U69 ( .I1(A[27]), .I2(n59), .O(n62) );
  NAND_GATE U70 ( .I1(n63), .I2(n64), .O(SUM[27]) );
  OR_GATE U71 ( .I1(n26), .I2(n59), .O(n64) );
  NAND_GATE U72 ( .I1(n59), .I2(n26), .O(n63) );
  AND3_GATE U73 ( .I1(A[25]), .I2(n65), .I3(A[26]), .O(n59) );
  NAND_GATE U74 ( .I1(n66), .I2(n67), .O(SUM[26]) );
  OR_GATE U75 ( .I1(n25), .I2(n68), .O(n67) );
  NAND_GATE U76 ( .I1(n68), .I2(n25), .O(n66) );
  AND_GATE U77 ( .I1(A[25]), .I2(n65), .O(n68) );
  NAND_GATE U78 ( .I1(n69), .I2(n70), .O(SUM[25]) );
  OR_GATE U79 ( .I1(n24), .I2(n65), .O(n70) );
  NAND_GATE U80 ( .I1(n65), .I2(n24), .O(n69) );
  AND3_GATE U81 ( .I1(A[23]), .I2(n71), .I3(A[24]), .O(n65) );
  NAND_GATE U82 ( .I1(n72), .I2(n73), .O(SUM[24]) );
  OR_GATE U83 ( .I1(n23), .I2(n74), .O(n73) );
  NAND_GATE U84 ( .I1(n74), .I2(n23), .O(n72) );
  AND_GATE U85 ( .I1(A[23]), .I2(n71), .O(n74) );
  NAND_GATE U86 ( .I1(n75), .I2(n76), .O(SUM[23]) );
  OR_GATE U87 ( .I1(n22), .I2(n71), .O(n76) );
  NAND_GATE U88 ( .I1(n71), .I2(n22), .O(n75) );
  AND3_GATE U89 ( .I1(A[21]), .I2(n77), .I3(A[22]), .O(n71) );
  NAND_GATE U90 ( .I1(n78), .I2(n79), .O(SUM[22]) );
  OR_GATE U91 ( .I1(n21), .I2(n80), .O(n79) );
  NAND_GATE U92 ( .I1(n80), .I2(n21), .O(n78) );
  AND_GATE U93 ( .I1(A[21]), .I2(n77), .O(n80) );
  NAND_GATE U94 ( .I1(n81), .I2(n82), .O(SUM[21]) );
  OR_GATE U95 ( .I1(n20), .I2(n77), .O(n82) );
  NAND_GATE U96 ( .I1(n77), .I2(n20), .O(n81) );
  AND3_GATE U97 ( .I1(A[19]), .I2(n83), .I3(A[20]), .O(n77) );
  NAND_GATE U98 ( .I1(n84), .I2(n85), .O(SUM[20]) );
  OR_GATE U99 ( .I1(n19), .I2(n86), .O(n85) );
  NAND_GATE U100 ( .I1(n86), .I2(n19), .O(n84) );
  AND_GATE U101 ( .I1(A[19]), .I2(n83), .O(n86) );
  NAND_GATE U102 ( .I1(n87), .I2(n88), .O(SUM[19]) );
  OR_GATE U103 ( .I1(n18), .I2(n83), .O(n88) );
  NAND_GATE U104 ( .I1(n83), .I2(n18), .O(n87) );
  AND3_GATE U105 ( .I1(A[17]), .I2(n89), .I3(A[18]), .O(n83) );
  NAND_GATE U106 ( .I1(n90), .I2(n91), .O(SUM[18]) );
  OR_GATE U107 ( .I1(n17), .I2(n92), .O(n91) );
  NAND_GATE U108 ( .I1(n92), .I2(n17), .O(n90) );
  AND_GATE U109 ( .I1(A[17]), .I2(n89), .O(n92) );
  NAND_GATE U110 ( .I1(n93), .I2(n94), .O(SUM[17]) );
  OR_GATE U111 ( .I1(n16), .I2(n89), .O(n94) );
  NAND_GATE U112 ( .I1(n89), .I2(n16), .O(n93) );
  AND3_GATE U113 ( .I1(A[15]), .I2(n95), .I3(A[16]), .O(n89) );
  NAND_GATE U114 ( .I1(n96), .I2(n97), .O(SUM[16]) );
  OR_GATE U115 ( .I1(n15), .I2(n98), .O(n97) );
  NAND_GATE U116 ( .I1(n98), .I2(n15), .O(n96) );
  AND_GATE U117 ( .I1(A[15]), .I2(n95), .O(n98) );
  NAND_GATE U118 ( .I1(n99), .I2(n100), .O(SUM[15]) );
  OR_GATE U119 ( .I1(n14), .I2(n95), .O(n100) );
  NAND_GATE U120 ( .I1(n95), .I2(n14), .O(n99) );
  AND3_GATE U121 ( .I1(A[13]), .I2(n101), .I3(A[14]), .O(n95) );
  NAND_GATE U122 ( .I1(n102), .I2(n103), .O(SUM[14]) );
  OR_GATE U123 ( .I1(n13), .I2(n104), .O(n103) );
  NAND_GATE U124 ( .I1(n104), .I2(n13), .O(n102) );
  AND_GATE U125 ( .I1(A[13]), .I2(n101), .O(n104) );
  NAND_GATE U126 ( .I1(n105), .I2(n106), .O(SUM[13]) );
  OR_GATE U127 ( .I1(n12), .I2(n101), .O(n106) );
  NAND_GATE U128 ( .I1(n101), .I2(n12), .O(n105) );
  AND3_GATE U129 ( .I1(A[11]), .I2(n2), .I3(A[12]), .O(n101) );
  NAND_GATE U130 ( .I1(n107), .I2(n108), .O(SUM[12]) );
  OR_GATE U131 ( .I1(n11), .I2(n109), .O(n108) );
  NAND_GATE U132 ( .I1(n109), .I2(n11), .O(n107) );
  AND_GATE U133 ( .I1(A[11]), .I2(n2), .O(n109) );
  NAND_GATE U134 ( .I1(n110), .I2(n111), .O(SUM[11]) );
  NAND_GATE U135 ( .I1(A[11]), .I2(n112), .O(n111) );
  NAND_GATE U136 ( .I1(n2), .I2(n10), .O(n110) );
  NAND3_GATE U137 ( .I1(n32), .I2(A[9]), .I3(A[10]), .O(n112) );
  NAND_GATE U138 ( .I1(n113), .I2(n114), .O(SUM[10]) );
  NAND_GATE U139 ( .I1(A[10]), .I2(n115), .O(n114) );
  OR_GATE U140 ( .I1(n115), .I2(A[10]), .O(n113) );
  NAND_GATE U141 ( .I1(n32), .I2(A[9]), .O(n115) );
  AND3_GATE U142 ( .I1(A[7]), .I2(n36), .I3(A[8]), .O(n32) );
  AND3_GATE U143 ( .I1(A[5]), .I2(n42), .I3(A[6]), .O(n36) );
  AND3_GATE U144 ( .I1(A[3]), .I2(A[2]), .I3(A[4]), .O(n42) );
endmodule


module predict_nb_record3_1_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117;

  INV_GATE U1 ( .I1(A[1]), .O(n1) );
  INV_GATE U2 ( .I1(A[2]), .O(n2) );
  INV_GATE U3 ( .I1(A[3]), .O(n3) );
  INV_GATE U4 ( .I1(A[4]), .O(n4) );
  INV_GATE U5 ( .I1(A[5]), .O(n5) );
  INV_GATE U6 ( .I1(A[6]), .O(n6) );
  INV_GATE U7 ( .I1(A[7]), .O(n7) );
  INV_GATE U8 ( .I1(A[8]), .O(n8) );
  INV_GATE U9 ( .I1(A[9]), .O(n9) );
  INV_GATE U10 ( .I1(A[10]), .O(n10) );
  INV_GATE U11 ( .I1(A[11]), .O(n11) );
  INV_GATE U12 ( .I1(A[12]), .O(n12) );
  INV_GATE U13 ( .I1(A[13]), .O(n13) );
  INV_GATE U14 ( .I1(A[14]), .O(n14) );
  INV_GATE U15 ( .I1(A[15]), .O(n15) );
  INV_GATE U16 ( .I1(A[16]), .O(n16) );
  INV_GATE U17 ( .I1(A[17]), .O(n17) );
  INV_GATE U18 ( .I1(A[18]), .O(n18) );
  INV_GATE U19 ( .I1(A[19]), .O(n19) );
  INV_GATE U20 ( .I1(A[20]), .O(n20) );
  INV_GATE U21 ( .I1(A[21]), .O(n21) );
  INV_GATE U22 ( .I1(A[22]), .O(n22) );
  INV_GATE U23 ( .I1(A[23]), .O(n23) );
  INV_GATE U24 ( .I1(A[24]), .O(n24) );
  INV_GATE U25 ( .I1(A[25]), .O(n25) );
  INV_GATE U26 ( .I1(A[26]), .O(n26) );
  INV_GATE U27 ( .I1(A[27]), .O(n27) );
  INV_GATE U28 ( .I1(A[28]), .O(n28) );
  INV_GATE U29 ( .I1(A[29]), .O(n29) );
  INV_GATE U30 ( .I1(A[30]), .O(n30) );
  INV_GATE U31 ( .I1(A[31]), .O(n31) );
  INV_GATE U32 ( .I1(B[0]), .O(n32) );
  NAND4_GATE U33 ( .I1(n33), .I2(n34), .I3(n35), .I4(n36), .O(NE) );
  AND4_GATE U34 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .O(n36) );
  AND5_GATE U35 ( .I1(n41), .I2(n42), .I3(n43), .I4(n44), .I5(n45), .O(n40) );
  AND4_GATE U36 ( .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n45) );
  NAND_GATE U37 ( .I1(B[16]), .I2(n16), .O(n49) );
  OR_GATE U38 ( .I1(n16), .I2(B[16]), .O(n48) );
  NAND_GATE U39 ( .I1(B[17]), .I2(n17), .O(n47) );
  OR_GATE U40 ( .I1(n17), .I2(B[17]), .O(n46) );
  NAND_GATE U41 ( .I1(B[18]), .I2(n18), .O(n44) );
  OR_GATE U42 ( .I1(n18), .I2(B[18]), .O(n43) );
  NAND_GATE U43 ( .I1(B[19]), .I2(n19), .O(n42) );
  OR_GATE U44 ( .I1(n19), .I2(B[19]), .O(n41) );
  AND5_GATE U45 ( .I1(n50), .I2(n51), .I3(n52), .I4(n53), .I5(n54), .O(n39) );
  AND4_GATE U46 ( .I1(n55), .I2(n56), .I3(n57), .I4(n58), .O(n54) );
  NAND_GATE U47 ( .I1(B[20]), .I2(n20), .O(n58) );
  OR_GATE U48 ( .I1(n20), .I2(B[20]), .O(n57) );
  NAND_GATE U49 ( .I1(B[21]), .I2(n21), .O(n56) );
  OR_GATE U50 ( .I1(n21), .I2(B[21]), .O(n55) );
  NAND_GATE U51 ( .I1(B[22]), .I2(n22), .O(n53) );
  OR_GATE U52 ( .I1(n22), .I2(B[22]), .O(n52) );
  NAND_GATE U53 ( .I1(B[23]), .I2(n23), .O(n51) );
  OR_GATE U54 ( .I1(n23), .I2(B[23]), .O(n50) );
  AND5_GATE U55 ( .I1(n59), .I2(n60), .I3(n61), .I4(n62), .I5(n63), .O(n38) );
  AND4_GATE U56 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n63) );
  NAND_GATE U57 ( .I1(B[24]), .I2(n24), .O(n67) );
  OR_GATE U58 ( .I1(n24), .I2(B[24]), .O(n66) );
  NAND_GATE U59 ( .I1(B[25]), .I2(n25), .O(n65) );
  OR_GATE U60 ( .I1(n25), .I2(B[25]), .O(n64) );
  NAND_GATE U61 ( .I1(B[26]), .I2(n26), .O(n62) );
  OR_GATE U62 ( .I1(n26), .I2(B[26]), .O(n61) );
  NAND_GATE U63 ( .I1(B[27]), .I2(n27), .O(n60) );
  OR_GATE U64 ( .I1(n27), .I2(B[27]), .O(n59) );
  AND5_GATE U65 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .I5(n72), .O(n37) );
  AND4_GATE U66 ( .I1(n73), .I2(n74), .I3(n75), .I4(n76), .O(n72) );
  NAND_GATE U67 ( .I1(B[28]), .I2(n28), .O(n76) );
  OR_GATE U68 ( .I1(n28), .I2(B[28]), .O(n75) );
  NAND_GATE U69 ( .I1(B[29]), .I2(n29), .O(n74) );
  OR_GATE U70 ( .I1(n29), .I2(B[29]), .O(n73) );
  NAND_GATE U71 ( .I1(B[30]), .I2(n30), .O(n71) );
  OR_GATE U72 ( .I1(n30), .I2(B[30]), .O(n70) );
  NAND_GATE U73 ( .I1(B[31]), .I2(n31), .O(n69) );
  OR_GATE U74 ( .I1(n31), .I2(B[31]), .O(n68) );
  AND5_GATE U75 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n35) );
  AND4_GATE U76 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(n81) );
  NAND_GATE U77 ( .I1(B[4]), .I2(n4), .O(n85) );
  OR_GATE U78 ( .I1(n4), .I2(B[4]), .O(n84) );
  NAND_GATE U79 ( .I1(B[5]), .I2(n5), .O(n83) );
  OR_GATE U80 ( .I1(n5), .I2(B[5]), .O(n82) );
  AND4_GATE U81 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(n80) );
  NAND_GATE U82 ( .I1(B[6]), .I2(n6), .O(n89) );
  OR_GATE U83 ( .I1(n6), .I2(B[6]), .O(n88) );
  NAND_GATE U84 ( .I1(B[7]), .I2(n7), .O(n87) );
  OR_GATE U85 ( .I1(n7), .I2(B[7]), .O(n86) );
  AND4_GATE U86 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(n79) );
  NAND_GATE U87 ( .I1(B[2]), .I2(n2), .O(n93) );
  OR_GATE U88 ( .I1(n2), .I2(B[2]), .O(n92) );
  NAND_GATE U89 ( .I1(B[3]), .I2(n3), .O(n91) );
  OR_GATE U90 ( .I1(n3), .I2(B[3]), .O(n90) );
  NAND_GATE U91 ( .I1(n94), .I2(n95), .O(n78) );
  NAND_GATE U92 ( .I1(B[1]), .I2(n96), .O(n95) );
  NAND_GATE U93 ( .I1(n96), .I2(n1), .O(n94) );
  NAND_GATE U94 ( .I1(A[0]), .I2(n32), .O(n96) );
  NAND_GATE U95 ( .I1(n97), .I2(n98), .O(n77) );
  OR_GATE U96 ( .I1(n99), .I2(B[1]), .O(n98) );
  OR_GATE U97 ( .I1(n1), .I2(n99), .O(n97) );
  NOR_GATE U98 ( .I1(n32), .I2(A[0]), .O(n99) );
  AND5_GATE U99 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .I5(n104), .O(
        n34) );
  AND4_GATE U100 ( .I1(n105), .I2(n106), .I3(n107), .I4(n108), .O(n104) );
  NAND_GATE U101 ( .I1(B[8]), .I2(n8), .O(n108) );
  OR_GATE U102 ( .I1(n8), .I2(B[8]), .O(n107) );
  NAND_GATE U103 ( .I1(B[9]), .I2(n9), .O(n106) );
  OR_GATE U104 ( .I1(n9), .I2(B[9]), .O(n105) );
  NAND_GATE U105 ( .I1(B[10]), .I2(n10), .O(n103) );
  OR_GATE U106 ( .I1(n10), .I2(B[10]), .O(n102) );
  NAND_GATE U107 ( .I1(B[11]), .I2(n11), .O(n101) );
  OR_GATE U108 ( .I1(n11), .I2(B[11]), .O(n100) );
  AND5_GATE U109 ( .I1(n109), .I2(n110), .I3(n111), .I4(n112), .I5(n113), .O(
        n33) );
  AND4_GATE U110 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(n113) );
  NAND_GATE U111 ( .I1(B[12]), .I2(n12), .O(n117) );
  OR_GATE U112 ( .I1(n12), .I2(B[12]), .O(n116) );
  NAND_GATE U113 ( .I1(B[13]), .I2(n13), .O(n115) );
  OR_GATE U114 ( .I1(n13), .I2(B[13]), .O(n114) );
  NAND_GATE U115 ( .I1(B[14]), .I2(n14), .O(n112) );
  OR_GATE U116 ( .I1(n14), .I2(B[14]), .O(n111) );
  NAND_GATE U117 ( .I1(B[15]), .I2(n15), .O(n110) );
  OR_GATE U118 ( .I1(n15), .I2(B[15]), .O(n109) );
endmodule


module predict_nb_record3_1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_GATE U1 ( .I1(A[30]), .O(n1) );
  INV_GATE U2 ( .I1(A[29]), .O(n2) );
  INV_GATE U3 ( .I1(A[28]), .O(n3) );
  INV_GATE U4 ( .I1(A[27]), .O(n4) );
  INV_GATE U5 ( .I1(A[26]), .O(n5) );
  INV_GATE U6 ( .I1(A[25]), .O(n6) );
  INV_GATE U7 ( .I1(A[24]), .O(n7) );
  INV_GATE U8 ( .I1(A[23]), .O(n8) );
  INV_GATE U9 ( .I1(A[22]), .O(n9) );
  INV_GATE U10 ( .I1(A[21]), .O(n10) );
  INV_GATE U11 ( .I1(A[20]), .O(n11) );
  INV_GATE U12 ( .I1(A[19]), .O(n12) );
  INV_GATE U13 ( .I1(A[18]), .O(n13) );
  INV_GATE U14 ( .I1(A[17]), .O(n14) );
  INV_GATE U15 ( .I1(A[16]), .O(n15) );
  INV_GATE U16 ( .I1(A[15]), .O(n16) );
  INV_GATE U17 ( .I1(A[14]), .O(n17) );
  INV_GATE U18 ( .I1(A[13]), .O(n18) );
  INV_GATE U19 ( .I1(A[12]), .O(n19) );
  INV_GATE U20 ( .I1(A[11]), .O(n20) );
  INV_GATE U21 ( .I1(n112), .O(n21) );
  INV_GATE U22 ( .I1(A[8]), .O(n22) );
  INV_GATE U23 ( .I1(n32), .O(n23) );
  INV_GATE U24 ( .I1(A[7]), .O(n24) );
  INV_GATE U25 ( .I1(A[6]), .O(n25) );
  INV_GATE U26 ( .I1(A[5]), .O(n26) );
  INV_GATE U27 ( .I1(A[4]), .O(n27) );
  INV_GATE U28 ( .I1(A[3]), .O(n28) );
  INV_GATE U29 ( .I1(A[2]), .O(SUM[2]) );
  NAND_GATE U30 ( .I1(n30), .I2(n31), .O(SUM[9]) );
  NAND_GATE U31 ( .I1(A[9]), .I2(n23), .O(n31) );
  OR_GATE U32 ( .I1(n23), .I2(A[9]), .O(n30) );
  NAND_GATE U33 ( .I1(n33), .I2(n34), .O(SUM[8]) );
  OR_GATE U34 ( .I1(n22), .I2(n35), .O(n34) );
  NAND_GATE U35 ( .I1(n35), .I2(n22), .O(n33) );
  AND_GATE U36 ( .I1(A[7]), .I2(n36), .O(n35) );
  NAND_GATE U37 ( .I1(n37), .I2(n38), .O(SUM[7]) );
  OR_GATE U38 ( .I1(n24), .I2(n36), .O(n38) );
  NAND_GATE U39 ( .I1(n36), .I2(n24), .O(n37) );
  NAND_GATE U40 ( .I1(n39), .I2(n40), .O(SUM[6]) );
  OR_GATE U41 ( .I1(n25), .I2(n41), .O(n40) );
  NAND_GATE U42 ( .I1(n41), .I2(n25), .O(n39) );
  AND_GATE U43 ( .I1(A[5]), .I2(n42), .O(n41) );
  NAND_GATE U44 ( .I1(n43), .I2(n44), .O(SUM[5]) );
  OR_GATE U45 ( .I1(n26), .I2(n42), .O(n44) );
  NAND_GATE U46 ( .I1(n42), .I2(n26), .O(n43) );
  NAND_GATE U47 ( .I1(n45), .I2(n46), .O(SUM[4]) );
  OR_GATE U48 ( .I1(n27), .I2(n47), .O(n46) );
  NAND_GATE U49 ( .I1(n47), .I2(n27), .O(n45) );
  AND_GATE U50 ( .I1(A[3]), .I2(A[2]), .O(n47) );
  NAND_GATE U51 ( .I1(n48), .I2(n49), .O(SUM[3]) );
  NAND_GATE U52 ( .I1(A[3]), .I2(SUM[2]), .O(n49) );
  NAND_GATE U53 ( .I1(A[2]), .I2(n28), .O(n48) );
  NAND_GATE U54 ( .I1(n50), .I2(n51), .O(SUM[31]) );
  NAND_GATE U55 ( .I1(A[31]), .I2(n52), .O(n51) );
  OR_GATE U56 ( .I1(n52), .I2(A[31]), .O(n50) );
  NAND_GATE U57 ( .I1(A[30]), .I2(n53), .O(n52) );
  NAND_GATE U58 ( .I1(n54), .I2(n55), .O(SUM[30]) );
  OR_GATE U59 ( .I1(n1), .I2(n53), .O(n55) );
  NAND_GATE U60 ( .I1(n53), .I2(n1), .O(n54) );
  AND_GATE U61 ( .I1(A[29]), .I2(n56), .O(n53) );
  NAND_GATE U62 ( .I1(n57), .I2(n58), .O(SUM[29]) );
  OR_GATE U63 ( .I1(n2), .I2(n56), .O(n58) );
  NAND_GATE U64 ( .I1(n56), .I2(n2), .O(n57) );
  AND3_GATE U65 ( .I1(A[27]), .I2(n59), .I3(A[28]), .O(n56) );
  NAND_GATE U66 ( .I1(n60), .I2(n61), .O(SUM[28]) );
  OR_GATE U67 ( .I1(n3), .I2(n62), .O(n61) );
  NAND_GATE U68 ( .I1(n62), .I2(n3), .O(n60) );
  AND_GATE U69 ( .I1(A[27]), .I2(n59), .O(n62) );
  NAND_GATE U70 ( .I1(n63), .I2(n64), .O(SUM[27]) );
  OR_GATE U71 ( .I1(n4), .I2(n59), .O(n64) );
  NAND_GATE U72 ( .I1(n59), .I2(n4), .O(n63) );
  AND3_GATE U73 ( .I1(A[25]), .I2(n65), .I3(A[26]), .O(n59) );
  NAND_GATE U74 ( .I1(n66), .I2(n67), .O(SUM[26]) );
  OR_GATE U75 ( .I1(n5), .I2(n68), .O(n67) );
  NAND_GATE U76 ( .I1(n68), .I2(n5), .O(n66) );
  AND_GATE U77 ( .I1(A[25]), .I2(n65), .O(n68) );
  NAND_GATE U78 ( .I1(n69), .I2(n70), .O(SUM[25]) );
  OR_GATE U79 ( .I1(n6), .I2(n65), .O(n70) );
  NAND_GATE U80 ( .I1(n65), .I2(n6), .O(n69) );
  AND3_GATE U81 ( .I1(A[23]), .I2(n71), .I3(A[24]), .O(n65) );
  NAND_GATE U82 ( .I1(n72), .I2(n73), .O(SUM[24]) );
  OR_GATE U83 ( .I1(n7), .I2(n74), .O(n73) );
  NAND_GATE U84 ( .I1(n74), .I2(n7), .O(n72) );
  AND_GATE U85 ( .I1(A[23]), .I2(n71), .O(n74) );
  NAND_GATE U86 ( .I1(n75), .I2(n76), .O(SUM[23]) );
  OR_GATE U87 ( .I1(n8), .I2(n71), .O(n76) );
  NAND_GATE U88 ( .I1(n71), .I2(n8), .O(n75) );
  AND3_GATE U89 ( .I1(A[21]), .I2(n77), .I3(A[22]), .O(n71) );
  NAND_GATE U90 ( .I1(n78), .I2(n79), .O(SUM[22]) );
  OR_GATE U91 ( .I1(n9), .I2(n80), .O(n79) );
  NAND_GATE U92 ( .I1(n80), .I2(n9), .O(n78) );
  AND_GATE U93 ( .I1(A[21]), .I2(n77), .O(n80) );
  NAND_GATE U94 ( .I1(n81), .I2(n82), .O(SUM[21]) );
  OR_GATE U95 ( .I1(n10), .I2(n77), .O(n82) );
  NAND_GATE U96 ( .I1(n77), .I2(n10), .O(n81) );
  AND3_GATE U97 ( .I1(A[19]), .I2(n83), .I3(A[20]), .O(n77) );
  NAND_GATE U98 ( .I1(n84), .I2(n85), .O(SUM[20]) );
  OR_GATE U99 ( .I1(n11), .I2(n86), .O(n85) );
  NAND_GATE U100 ( .I1(n86), .I2(n11), .O(n84) );
  AND_GATE U101 ( .I1(A[19]), .I2(n83), .O(n86) );
  NAND_GATE U102 ( .I1(n87), .I2(n88), .O(SUM[19]) );
  OR_GATE U103 ( .I1(n12), .I2(n83), .O(n88) );
  NAND_GATE U104 ( .I1(n83), .I2(n12), .O(n87) );
  AND3_GATE U105 ( .I1(A[17]), .I2(n89), .I3(A[18]), .O(n83) );
  NAND_GATE U106 ( .I1(n90), .I2(n91), .O(SUM[18]) );
  OR_GATE U107 ( .I1(n13), .I2(n92), .O(n91) );
  NAND_GATE U108 ( .I1(n92), .I2(n13), .O(n90) );
  AND_GATE U109 ( .I1(A[17]), .I2(n89), .O(n92) );
  NAND_GATE U110 ( .I1(n93), .I2(n94), .O(SUM[17]) );
  OR_GATE U111 ( .I1(n14), .I2(n89), .O(n94) );
  NAND_GATE U112 ( .I1(n89), .I2(n14), .O(n93) );
  AND3_GATE U113 ( .I1(A[15]), .I2(n95), .I3(A[16]), .O(n89) );
  NAND_GATE U114 ( .I1(n96), .I2(n97), .O(SUM[16]) );
  OR_GATE U115 ( .I1(n15), .I2(n98), .O(n97) );
  NAND_GATE U116 ( .I1(n98), .I2(n15), .O(n96) );
  AND_GATE U117 ( .I1(A[15]), .I2(n95), .O(n98) );
  NAND_GATE U118 ( .I1(n99), .I2(n100), .O(SUM[15]) );
  OR_GATE U119 ( .I1(n16), .I2(n95), .O(n100) );
  NAND_GATE U120 ( .I1(n95), .I2(n16), .O(n99) );
  AND3_GATE U121 ( .I1(A[13]), .I2(n101), .I3(A[14]), .O(n95) );
  NAND_GATE U122 ( .I1(n102), .I2(n103), .O(SUM[14]) );
  OR_GATE U123 ( .I1(n17), .I2(n104), .O(n103) );
  NAND_GATE U124 ( .I1(n104), .I2(n17), .O(n102) );
  AND_GATE U125 ( .I1(A[13]), .I2(n101), .O(n104) );
  NAND_GATE U126 ( .I1(n105), .I2(n106), .O(SUM[13]) );
  OR_GATE U127 ( .I1(n18), .I2(n101), .O(n106) );
  NAND_GATE U128 ( .I1(n101), .I2(n18), .O(n105) );
  AND3_GATE U129 ( .I1(A[11]), .I2(n21), .I3(A[12]), .O(n101) );
  NAND_GATE U130 ( .I1(n107), .I2(n108), .O(SUM[12]) );
  OR_GATE U131 ( .I1(n19), .I2(n109), .O(n108) );
  NAND_GATE U132 ( .I1(n109), .I2(n19), .O(n107) );
  AND_GATE U133 ( .I1(A[11]), .I2(n21), .O(n109) );
  NAND_GATE U134 ( .I1(n110), .I2(n111), .O(SUM[11]) );
  NAND_GATE U135 ( .I1(A[11]), .I2(n112), .O(n111) );
  NAND_GATE U136 ( .I1(n21), .I2(n20), .O(n110) );
  NAND3_GATE U137 ( .I1(n32), .I2(A[9]), .I3(A[10]), .O(n112) );
  NAND_GATE U138 ( .I1(n113), .I2(n114), .O(SUM[10]) );
  NAND_GATE U139 ( .I1(A[10]), .I2(n115), .O(n114) );
  OR_GATE U140 ( .I1(n115), .I2(A[10]), .O(n113) );
  NAND_GATE U141 ( .I1(n32), .I2(A[9]), .O(n115) );
  AND3_GATE U142 ( .I1(A[7]), .I2(n36), .I3(A[8]), .O(n32) );
  AND3_GATE U143 ( .I1(A[5]), .I2(n42), .I3(A[6]), .O(n36) );
  AND3_GATE U144 ( .I1(A[3]), .I2(A[2]), .I3(A[4]), .O(n42) );
endmodule


module alu ( clock, reset, op1, op2, ctrl, res, overflow );
  input [31:0] op1;
  input [31:0] op2;
  input [27:0] ctrl;
  output [31:0] res;
  input clock, reset;
  output overflow;
  wire   \efct_op1[32] , N710, N711, N712, N713, N714, N715, N716, N717, N718,
         N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729,
         N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740,
         N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751,
         N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762,
         N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838, N1035, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n169, n170, n171,
         n172, n174, n175, n177, n178, n205, n206, n207, n208, n209, n210,
         n211, n212, n214, n215, n216, n222, n223, n224, n225, n226, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n251, n253, n254, n255, n256, n257, n258, n269, n270, n271, n272,
         n273, n274, n275, n276, n278, n279, n280, n281, n284, n286, n287,
         n288, n289, n290, n291, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n314, n316, n317, n318, n319, n320, n321, n327,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n344, n346, n348, n349, n350, n351, n352, n361, n362, n363, n364,
         n365, n374, n375, n376, n377, n379, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n396, n397, n398, n399, n400,
         n401, n403, n417, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n479, n481, n482, n483, n484,
         n485, n493, n494, n495, n496, n497, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n522, n523, n525, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n562, n563,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n612, n613, n614, n615, n619, n631, n632, n652, n653, n654, n655,
         n657, n667, n672, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n709, n710, n715, n716, n717,
         n731, n732, n733, n734, n735, n737, n738, n740, n741, n751, n752,
         n757, n758, n759, n760, n774, n775, n776, n777, n778, n779, n780,
         n781, n791, n792, n793, n794, n799, n800, n801, n802, n816, n817,
         n818, n819, n820, n821, n822, n823, n833, n834, n835, n840, n841,
         n842, n843, n844, n858, n859, n860, n861, n862, n863, n873, n874,
         n875, n880, n881, n882, n896, n897, n898, n899, n909, n910, n911,
         n916, n917, n918, n919, n920, n921, n922, n923, n931, n932, n933,
         n934, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n964, n965, n967, n982, n983, n984, n985, n995, n996, n997,
         n1002, n1003, n1004, n1005, n1020, n1021, n1022, n1023, n1033, n1034,
         n1035, n1036, n1037, n1042, n1043, n1044, n1045, n1059, n1060, n1061,
         n1062, n1072, n1073, n1074, n1075, n1080, n1081, n1082, n1083, n1096,
         n1097, n1098, n1099, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1145, n1146, n1147, n1148, n1149, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1216, n1217, n1218, n1219, n1221, n1222, n1223,
         n1224, n1225, n1230, n1231, n1232, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1290, n1291, n1292, n1293, n1294, n1295, n1318, n1319, n1320, n1321,
         n1322, n1323, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1338,
         n1343, n1344, n1345, n1346, n1347, n1348, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1411, n1412, n1413,
         n1414, n1415, n1416, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1446, n1457, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1505, n1506, n1697, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1909, n1910, n1911, n1922, n1923, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n168, n173, n176, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n213, n217, n218, n219, n220, n221, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n249, n250, n252, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n277, n282, n283,
         n285, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n312, n313, n315, n322, n323, n324, n325, n326, n328, n329, n330,
         n342, n343, n345, n347, n353, n354, n355, n356, n357, n358, n359,
         n360, n366, n367, n368, n369, n370, n371, n372, n373, n378, n380,
         n392, n393, n394, n395, n402, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n418, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n470, n471, n472, n473, n474, n475, n476, n477, n478, n480,
         n486, n487, n488, n489, n490, n491, n492, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n518, n519, n520, n521, n524, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n558, n559,
         n560, n561, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n616, n617, n618, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n656, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n668, n669, n670, n671, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n711, n712,
         n713, n714, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n736, n739, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n753, n754, n755, n756, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n795, n796, n797,
         n798, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n836, n837, n838, n839, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n876, n877, n878, n879, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n912, n913,
         n914, n915, n924, n925, n926, n927, n928, n929, n930, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n956, n957, n958,
         n959, n960, n961, n962, n963, n966, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n998, n999, n1000, n1001,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1038, n1039, n1040, n1041, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1076,
         n1077, n1078, n1079, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1212, n1213, n1214,
         n1215, n1220, n1226, n1227, n1228, n1229, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1287, n1288, n1289, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1324, n1325, n1326, n1327, n1335, n1336, n1337, n1339, n1340, n1341,
         n1342, n1349, n1350, n1351, n1352, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1407, n1408,
         n1409, n1410, n1417, n1418, n1419, n1420, n1421, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1458, n1459, n1460,
         n1461, n1462, n1463, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1499, n1500, n1501, n1502, n1503,
         n1504, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1924, n1925, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058;
  wire   [32:0] efct_op2;
  wire   [32:0] res_add;
  wire   [63:0] hilo;
  assign overflow = N1035;

  FLIP_FLOP_D \hilo_reg[63]  ( .D(n1926), .CK(clock), .Q(hilo[63]) );
  FLIP_FLOP_D \hilo_reg[62]  ( .D(n1927), .CK(clock), .Q(hilo[62]) );
  FLIP_FLOP_D \hilo_reg[61]  ( .D(n1928), .CK(clock), .Q(hilo[61]) );
  FLIP_FLOP_D \hilo_reg[60]  ( .D(n1929), .CK(clock), .Q(hilo[60]) );
  FLIP_FLOP_D \hilo_reg[59]  ( .D(n1930), .CK(clock), .Q(hilo[59]) );
  FLIP_FLOP_D \hilo_reg[58]  ( .D(n1931), .CK(clock), .Q(hilo[58]) );
  FLIP_FLOP_D \hilo_reg[57]  ( .D(n1932), .CK(clock), .Q(hilo[57]) );
  FLIP_FLOP_D \hilo_reg[56]  ( .D(n1933), .CK(clock), .Q(hilo[56]) );
  FLIP_FLOP_D \hilo_reg[55]  ( .D(n1934), .CK(clock), .Q(hilo[55]) );
  FLIP_FLOP_D \hilo_reg[54]  ( .D(n1935), .CK(clock), .Q(hilo[54]) );
  FLIP_FLOP_D \hilo_reg[53]  ( .D(n1936), .CK(clock), .Q(hilo[53]) );
  FLIP_FLOP_D \hilo_reg[52]  ( .D(n1937), .CK(clock), .Q(hilo[52]) );
  FLIP_FLOP_D \hilo_reg[51]  ( .D(n1938), .CK(clock), .Q(hilo[51]) );
  FLIP_FLOP_D \hilo_reg[50]  ( .D(n1939), .CK(clock), .Q(hilo[50]) );
  FLIP_FLOP_D \hilo_reg[49]  ( .D(n1940), .CK(clock), .Q(hilo[49]) );
  FLIP_FLOP_D \hilo_reg[48]  ( .D(n1941), .CK(clock), .Q(hilo[48]) );
  FLIP_FLOP_D \hilo_reg[47]  ( .D(n1942), .CK(clock), .Q(hilo[47]) );
  FLIP_FLOP_D \hilo_reg[46]  ( .D(n1943), .CK(clock), .Q(hilo[46]) );
  FLIP_FLOP_D \hilo_reg[45]  ( .D(n1944), .CK(clock), .Q(hilo[45]) );
  FLIP_FLOP_D \hilo_reg[44]  ( .D(n1945), .CK(clock), .Q(hilo[44]) );
  FLIP_FLOP_D \hilo_reg[43]  ( .D(n1946), .CK(clock), .Q(hilo[43]) );
  FLIP_FLOP_D \hilo_reg[42]  ( .D(n1947), .CK(clock), .Q(hilo[42]) );
  FLIP_FLOP_D \hilo_reg[41]  ( .D(n1948), .CK(clock), .Q(hilo[41]) );
  FLIP_FLOP_D \hilo_reg[40]  ( .D(n1949), .CK(clock), .Q(hilo[40]) );
  FLIP_FLOP_D \hilo_reg[39]  ( .D(n1950), .CK(clock), .Q(hilo[39]) );
  FLIP_FLOP_D \hilo_reg[38]  ( .D(n1951), .CK(clock), .Q(hilo[38]) );
  FLIP_FLOP_D \hilo_reg[37]  ( .D(n1952), .CK(clock), .Q(hilo[37]) );
  FLIP_FLOP_D \hilo_reg[36]  ( .D(n1953), .CK(clock), .Q(hilo[36]) );
  FLIP_FLOP_D \hilo_reg[35]  ( .D(n1954), .CK(clock), .Q(hilo[35]) );
  FLIP_FLOP_D \hilo_reg[34]  ( .D(n1955), .CK(clock), .Q(hilo[34]) );
  FLIP_FLOP_D \hilo_reg[33]  ( .D(n1956), .CK(clock), .Q(hilo[33]) );
  FLIP_FLOP_D \hilo_reg[32]  ( .D(n1957), .CK(clock), .Q(hilo[32]) );
  FLIP_FLOP_D \hilo_reg[31]  ( .D(n1958), .CK(clock), .Q(hilo[31]) );
  FLIP_FLOP_D \hilo_reg[30]  ( .D(n1959), .CK(clock), .Q(hilo[30]) );
  FLIP_FLOP_D \hilo_reg[29]  ( .D(n1960), .CK(clock), .Q(hilo[29]) );
  FLIP_FLOP_D \hilo_reg[28]  ( .D(n1961), .CK(clock), .Q(hilo[28]) );
  FLIP_FLOP_D \hilo_reg[27]  ( .D(n1962), .CK(clock), .Q(hilo[27]) );
  FLIP_FLOP_D \hilo_reg[26]  ( .D(n1963), .CK(clock), .Q(hilo[26]) );
  FLIP_FLOP_D \hilo_reg[25]  ( .D(n1964), .CK(clock), .Q(hilo[25]) );
  FLIP_FLOP_D \hilo_reg[24]  ( .D(n1965), .CK(clock), .Q(hilo[24]) );
  FLIP_FLOP_D \hilo_reg[23]  ( .D(n1966), .CK(clock), .Q(hilo[23]) );
  FLIP_FLOP_D \hilo_reg[22]  ( .D(n1967), .CK(clock), .Q(hilo[22]) );
  FLIP_FLOP_D \hilo_reg[21]  ( .D(n1968), .CK(clock), .Q(hilo[21]) );
  FLIP_FLOP_D \hilo_reg[20]  ( .D(n1969), .CK(clock), .Q(hilo[20]) );
  FLIP_FLOP_D \hilo_reg[19]  ( .D(n1970), .CK(clock), .Q(hilo[19]) );
  FLIP_FLOP_D \hilo_reg[18]  ( .D(n1971), .CK(clock), .Q(hilo[18]) );
  FLIP_FLOP_D \hilo_reg[17]  ( .D(n1972), .CK(clock), .Q(hilo[17]) );
  FLIP_FLOP_D \hilo_reg[16]  ( .D(n1973), .CK(clock), .Q(hilo[16]) );
  FLIP_FLOP_D \hilo_reg[15]  ( .D(n1974), .CK(clock), .Q(hilo[15]) );
  FLIP_FLOP_D \hilo_reg[14]  ( .D(n1975), .CK(clock), .Q(hilo[14]) );
  FLIP_FLOP_D \hilo_reg[13]  ( .D(n1976), .CK(clock), .Q(hilo[13]) );
  FLIP_FLOP_D \hilo_reg[12]  ( .D(n1977), .CK(clock), .Q(hilo[12]) );
  FLIP_FLOP_D \hilo_reg[11]  ( .D(n1978), .CK(clock), .Q(hilo[11]) );
  FLIP_FLOP_D \hilo_reg[10]  ( .D(n1979), .CK(clock), .Q(hilo[10]) );
  FLIP_FLOP_D \hilo_reg[9]  ( .D(n1980), .CK(clock), .Q(hilo[9]) );
  FLIP_FLOP_D \hilo_reg[8]  ( .D(n1981), .CK(clock), .Q(hilo[8]) );
  FLIP_FLOP_D \hilo_reg[7]  ( .D(n1982), .CK(clock), .Q(hilo[7]) );
  FLIP_FLOP_D \hilo_reg[6]  ( .D(n1983), .CK(clock), .Q(hilo[6]) );
  FLIP_FLOP_D \hilo_reg[5]  ( .D(n1984), .CK(clock), .Q(hilo[5]) );
  FLIP_FLOP_D \hilo_reg[4]  ( .D(n1985), .CK(clock), .Q(hilo[4]) );
  FLIP_FLOP_D \hilo_reg[3]  ( .D(n1986), .CK(clock), .Q(hilo[3]) );
  FLIP_FLOP_D \hilo_reg[2]  ( .D(n1987), .CK(clock), .Q(hilo[2]) );
  FLIP_FLOP_D \hilo_reg[1]  ( .D(n1988), .CK(clock), .Q(hilo[1]) );
  FLIP_FLOP_D \hilo_reg[0]  ( .D(n1989), .CK(clock), .Q(hilo[0]) );
  NAND4_GATE U142 ( .I1(n160), .I2(n161), .I3(n162), .I4(n163), .O(n159) );
  AND3_GATE U143 ( .I1(n164), .I2(n165), .I3(n166), .O(n163) );
  NAND_GATE U144 ( .I1(n167), .I2(n2030), .O(n166) );
  OR_GATE U145 ( .I1(n169), .I2(n170), .O(n165) );
  OR_GATE U146 ( .I1(n171), .I2(n172), .O(n164) );
  NAND_GATE U147 ( .I1(n2041), .I2(n174), .O(n162) );
  NAND_GATE U148 ( .I1(n175), .I2(n2026), .O(n161) );
  NAND_GATE U149 ( .I1(n2042), .I2(n177), .O(n160) );
  NAND4_GATE U170 ( .I1(n206), .I2(n207), .I3(n208), .I4(n209), .O(n205) );
  AND3_GATE U171 ( .I1(n210), .I2(n211), .I3(n212), .O(n209) );
  NAND_GATE U172 ( .I1(n2043), .I2(n167), .O(n212) );
  NAND_GATE U173 ( .I1(n2035), .I2(n2046), .O(n211) );
  OR_GATE U174 ( .I1(n214), .I2(n171), .O(n210) );
  NAND_GATE U175 ( .I1(n2041), .I2(n215), .O(n208) );
  NAND_GATE U176 ( .I1(n2045), .I2(n175), .O(n207) );
  NAND_GATE U177 ( .I1(n216), .I2(n2042), .O(n206) );
  NAND5_GATE U188 ( .I1(n222), .I2(n223), .I3(n224), .I4(n225), .I5(n226), .O(
        res[7]) );
  NAND4_GATE U198 ( .I1(n238), .I2(n239), .I3(n240), .I4(n241), .O(n237) );
  AND3_GATE U199 ( .I1(n242), .I2(n243), .I3(n244), .O(n241) );
  NAND_GATE U200 ( .I1(n2031), .I2(n167), .O(n244) );
  OR_GATE U201 ( .I1(n245), .I2(n169), .O(n243) );
  OR_GATE U202 ( .I1(n246), .I2(n171), .O(n242) );
  NAND_GATE U203 ( .I1(n2041), .I2(n247), .O(n240) );
  NAND_GATE U204 ( .I1(n2024), .I2(n175), .O(n239) );
  NAND_GATE U205 ( .I1(n248), .I2(n2042), .O(n238) );
  NAND_GATE U211 ( .I1(op2[7]), .I2(n251), .O(n224) );
  NAND_GATE U215 ( .I1(n52), .I2(n253), .O(n222) );
  NAND5_GATE U216 ( .I1(n254), .I2(n255), .I3(n256), .I4(n257), .I5(n258), .O(
        res[6]) );
  NAND4_GATE U226 ( .I1(n270), .I2(n271), .I3(n272), .I4(n273), .O(n269) );
  AND3_GATE U227 ( .I1(n274), .I2(n275), .I3(n276), .O(n273) );
  NAND_GATE U228 ( .I1(n2034), .I2(n167), .O(n276) );
  OR_GATE U229 ( .I1(n278), .I2(n169), .O(n275) );
  OR_GATE U230 ( .I1(n279), .I2(n171), .O(n274) );
  NAND_GATE U231 ( .I1(n2041), .I2(n280), .O(n272) );
  NAND_GATE U232 ( .I1(n2025), .I2(n175), .O(n271) );
  NAND_GATE U233 ( .I1(n281), .I2(n2042), .O(n270) );
  NAND_GATE U239 ( .I1(op2[6]), .I2(n284), .O(n256) );
  NAND_GATE U243 ( .I1(n52), .I2(n286), .O(n254) );
  NAND5_GATE U244 ( .I1(n287), .I2(n288), .I3(n289), .I4(n290), .I5(n291), .O(
        res[5]) );
  NAND4_GATE U254 ( .I1(n303), .I2(n304), .I3(n305), .I4(n306), .O(n302) );
  AND3_GATE U255 ( .I1(n307), .I2(n308), .I3(n309), .O(n306) );
  NAND_GATE U256 ( .I1(n2026), .I2(n167), .O(n309) );
  NAND_GATE U257 ( .I1(n2030), .I2(n2046), .O(n308) );
  OR_GATE U258 ( .I1(n171), .I2(n170), .O(n307) );
  NAND_GATE U259 ( .I1(n2041), .I2(n310), .O(n305) );
  NAND_GATE U260 ( .I1(n2027), .I2(n175), .O(n304) );
  NAND_GATE U261 ( .I1(n311), .I2(n2042), .O(n303) );
  NAND_GATE U267 ( .I1(op2[5]), .I2(n314), .O(n289) );
  NAND_GATE U271 ( .I1(n52), .I2(n316), .O(n287) );
  NAND5_GATE U272 ( .I1(n317), .I2(n318), .I3(n319), .I4(n320), .I5(n321), .O(
        res[4]) );
  NAND4_GATE U280 ( .I1(n332), .I2(n333), .I3(n334), .I4(n335), .O(n331) );
  AND3_GATE U281 ( .I1(n336), .I2(n337), .I3(n338), .O(n335) );
  NAND_GATE U282 ( .I1(n2045), .I2(n167), .O(n338) );
  OR_GATE U283 ( .I1(n339), .I2(n169), .O(n337) );
  NAND_GATE U284 ( .I1(n2035), .I2(n2047), .O(n336) );
  NAND_GATE U285 ( .I1(n2041), .I2(n340), .O(n334) );
  NAND_GATE U286 ( .I1(n2044), .I2(n175), .O(n333) );
  NAND_GATE U287 ( .I1(n341), .I2(n2042), .O(n332) );
  NAND_GATE U293 ( .I1(op2[4]), .I2(n344), .O(n319) );
  NAND_GATE U296 ( .I1(op2[4]), .I2(n346), .O(n318) );
  NAND5_GATE U300 ( .I1(n348), .I2(n349), .I3(n350), .I4(n351), .I5(n352), .O(
        res[3]) );
  AND3_GATE U309 ( .I1(n362), .I2(n363), .I3(n364), .O(n351) );
  OR_GATE U319 ( .I1(n379), .I2(n114), .O(n365) );
  NAND_GATE U320 ( .I1(n6), .I2(n381), .O(n363) );
  NAND5_GATE U321 ( .I1(n382), .I2(n383), .I3(n384), .I4(n385), .I5(n386), .O(
        n381) );
  AND4_GATE U322 ( .I1(n387), .I2(n388), .I3(n389), .I4(n390), .O(n386) );
  NAND_GATE U323 ( .I1(n376), .I2(op2[6]), .O(n390) );
  NAND_GATE U324 ( .I1(n377), .I2(op2[5]), .O(n389) );
  NAND_GATE U325 ( .I1(n375), .I2(op2[4]), .O(n388) );
  NAND_GATE U326 ( .I1(n374), .I2(op2[3]), .O(n387) );
  OR_GATE U327 ( .I1(n391), .I2(n169), .O(n385) );
  OR_GATE U328 ( .I1(n245), .I2(n171), .O(n384) );
  NAND_GATE U329 ( .I1(n2024), .I2(n167), .O(n383) );
  NAND_GATE U335 ( .I1(n400), .I2(op1[4]), .O(n382) );
  NAND_GATE U336 ( .I1(hilo[3]), .I2(n178), .O(n362) );
  NAND_GATE U337 ( .I1(op2[3]), .I2(n401), .O(n350) );
  NAND_GATE U341 ( .I1(op1[3]), .I2(n403), .O(n348) );
  NAND5_GATE U350 ( .I1(n420), .I2(n421), .I3(n422), .I4(n423), .I5(n424), .O(
        n419) );
  AND4_GATE U351 ( .I1(n425), .I2(n426), .I3(n427), .I4(n428), .O(n424) );
  NAND_GATE U352 ( .I1(op2[28]), .I2(n376), .O(n428) );
  NAND_GATE U353 ( .I1(n377), .I2(op2[29]), .O(n427) );
  NAND_GATE U354 ( .I1(n375), .I2(op2[30]), .O(n426) );
  NAND_GATE U355 ( .I1(n374), .I2(op2[31]), .O(n425) );
  NAND_GATE U356 ( .I1(n2046), .I2(n429), .O(n423) );
  NAND_GATE U357 ( .I1(n2047), .I2(n430), .O(n422) );
  NAND_GATE U358 ( .I1(n167), .I2(n431), .O(n421) );
  NAND_GATE U359 ( .I1(n432), .I2(op1[4]), .O(n420) );
  AND4_GATE U384 ( .I1(n463), .I2(n464), .I3(n465), .I4(n466), .O(n462) );
  NAND_GATE U385 ( .I1(op2[27]), .I2(n376), .O(n466) );
  NAND_GATE U386 ( .I1(op2[28]), .I2(n377), .O(n465) );
  NAND_GATE U387 ( .I1(n375), .I2(op2[29]), .O(n464) );
  NAND_GATE U388 ( .I1(n374), .I2(op2[30]), .O(n463) );
  NAND_GATE U389 ( .I1(n2046), .I2(n467), .O(n461) );
  NAND_GATE U390 ( .I1(n2047), .I2(n468), .O(n460) );
  NAND_GATE U391 ( .I1(n167), .I2(n469), .O(n459) );
  NAND5_GATE U405 ( .I1(n481), .I2(n482), .I3(n483), .I4(n484), .I5(n485), .O(
        res[2]) );
  AND3_GATE U414 ( .I1(n494), .I2(n495), .I3(n496), .O(n484) );
  OR_GATE U424 ( .I1(n507), .I2(n114), .O(n497) );
  NAND_GATE U425 ( .I1(n6), .I2(n508), .O(n495) );
  NAND5_GATE U426 ( .I1(n509), .I2(n510), .I3(n511), .I4(n512), .I5(n513), .O(
        n508) );
  AND4_GATE U427 ( .I1(n514), .I2(n515), .I3(n516), .I4(n517), .O(n513) );
  NAND_GATE U428 ( .I1(n376), .I2(op2[5]), .O(n517) );
  NAND_GATE U429 ( .I1(n377), .I2(op2[4]), .O(n516) );
  NAND_GATE U430 ( .I1(n375), .I2(op2[3]), .O(n515) );
  NAND_GATE U431 ( .I1(n374), .I2(op2[2]), .O(n514) );
  NAND_GATE U432 ( .I1(n2034), .I2(n2046), .O(n512) );
  OR_GATE U433 ( .I1(n278), .I2(n171), .O(n511) );
  NAND_GATE U434 ( .I1(n2025), .I2(n167), .O(n510) );
  NAND_GATE U440 ( .I1(n522), .I2(op1[4]), .O(n509) );
  NAND_GATE U441 ( .I1(hilo[2]), .I2(n178), .O(n494) );
  NAND_GATE U442 ( .I1(op2[2]), .I2(n523), .O(n483) );
  NAND_GATE U446 ( .I1(op1[2]), .I2(n525), .O(n481) );
  AND4_GATE U465 ( .I1(n551), .I2(n552), .I3(n553), .I4(n554), .O(n550) );
  NAND_GATE U466 ( .I1(op2[26]), .I2(n376), .O(n554) );
  NAND_GATE U467 ( .I1(op2[27]), .I2(n377), .O(n553) );
  NAND_GATE U468 ( .I1(op2[28]), .I2(n375), .O(n552) );
  NAND_GATE U469 ( .I1(n374), .I2(op2[29]), .O(n551) );
  NAND_GATE U470 ( .I1(n2046), .I2(n555), .O(n549) );
  NAND_GATE U471 ( .I1(n2047), .I2(n556), .O(n548) );
  NAND_GATE U472 ( .I1(n167), .I2(n557), .O(n547) );
  AND4_GATE U491 ( .I1(n584), .I2(n585), .I3(n586), .I4(n587), .O(n583) );
  NAND_GATE U492 ( .I1(op2[25]), .I2(n376), .O(n587) );
  NAND_GATE U493 ( .I1(op2[26]), .I2(n377), .O(n586) );
  NAND_GATE U494 ( .I1(op2[27]), .I2(n375), .O(n585) );
  NAND_GATE U495 ( .I1(op2[28]), .I2(n374), .O(n584) );
  NAND_GATE U496 ( .I1(n2046), .I2(n588), .O(n582) );
  NAND_GATE U497 ( .I1(n2047), .I2(n589), .O(n581) );
  NAND_GATE U498 ( .I1(n167), .I2(n590), .O(n580) );
  NAND4_GATE U519 ( .I1(n612), .I2(n613), .I3(n614), .I4(n615), .O(n431) );
  NAND_GATE U520 ( .I1(op2[24]), .I2(n396), .O(n615) );
  NAND_GATE U521 ( .I1(op2[25]), .I2(n397), .O(n614) );
  NAND_GATE U522 ( .I1(op2[26]), .I2(n398), .O(n613) );
  NAND_GATE U523 ( .I1(op2[27]), .I2(n399), .O(n612) );
  NAND4_GATE U551 ( .I1(n652), .I2(n653), .I3(n654), .I4(n655), .O(n469) );
  NAND_GATE U552 ( .I1(op2[23]), .I2(n396), .O(n655) );
  NAND_GATE U553 ( .I1(op2[24]), .I2(n397), .O(n654) );
  NAND_GATE U554 ( .I1(op2[25]), .I2(n398), .O(n653) );
  NAND_GATE U555 ( .I1(op2[26]), .I2(n399), .O(n652) );
  NAND4_GATE U583 ( .I1(n686), .I2(n687), .I3(n688), .I4(n689), .O(n557) );
  NAND_GATE U584 ( .I1(op2[22]), .I2(n396), .O(n689) );
  NAND_GATE U585 ( .I1(op2[23]), .I2(n397), .O(n688) );
  NAND_GATE U586 ( .I1(op2[24]), .I2(n398), .O(n687) );
  NAND_GATE U587 ( .I1(op2[25]), .I2(n399), .O(n686) );
  NAND_GATE U591 ( .I1(n693), .I2(n694), .O(n692) );
  NAND_GATE U592 ( .I1(n695), .I2(n696), .O(n691) );
  NAND_GATE U593 ( .I1(n697), .I2(n698), .O(n690) );
  NAND_GATE U609 ( .I1(n709), .I2(n710), .O(n174) );
  NAND_GATE U610 ( .I1(n2057), .I2(n697), .O(n710) );
  NAND_GATE U611 ( .I1(n693), .I2(n562), .O(n709) );
  AND_GATE U615 ( .I1(n715), .I2(n716), .O(n177) );
  NAND_GATE U616 ( .I1(n697), .I2(n717), .O(n716) );
  NAND_GATE U617 ( .I1(n693), .I2(n563), .O(n715) );
  NAND4_GATE U625 ( .I1(n731), .I2(n732), .I3(n733), .I4(n734), .O(n590) );
  NAND_GATE U626 ( .I1(op2[21]), .I2(n396), .O(n734) );
  NAND_GATE U627 ( .I1(op2[22]), .I2(n397), .O(n733) );
  NAND_GATE U628 ( .I1(op2[23]), .I2(n398), .O(n732) );
  NAND_GATE U629 ( .I1(op2[24]), .I2(n399), .O(n731) );
  NAND_GATE U633 ( .I1(n693), .I2(n738), .O(n737) );
  NAND_GATE U635 ( .I1(n697), .I2(n740), .O(n735) );
  NAND_GATE U651 ( .I1(n751), .I2(n752), .O(n215) );
  NAND_GATE U652 ( .I1(n2052), .I2(n697), .O(n752) );
  NAND_GATE U653 ( .I1(n2049), .I2(n693), .O(n751) );
  AND_GATE U657 ( .I1(n757), .I2(n758), .O(n216) );
  NAND_GATE U658 ( .I1(n697), .I2(n759), .O(n758) );
  NAND_GATE U659 ( .I1(n693), .I2(n760), .O(n757) );
  NAND4_GATE U667 ( .I1(n774), .I2(n775), .I3(n776), .I4(n777), .O(n429) );
  NAND_GATE U668 ( .I1(op2[20]), .I2(n396), .O(n777) );
  NAND_GATE U669 ( .I1(op2[21]), .I2(n397), .O(n776) );
  NAND_GATE U670 ( .I1(op2[22]), .I2(n398), .O(n775) );
  NAND_GATE U671 ( .I1(op2[23]), .I2(n399), .O(n774) );
  NAND_GATE U674 ( .I1(n778), .I2(n779), .O(n253) );
  NAND_GATE U675 ( .I1(n697), .I2(n780), .O(n779) );
  NAND_GATE U676 ( .I1(n693), .I2(n361), .O(n778) );
  NAND3_GATE U692 ( .I1(n791), .I2(n792), .I3(n793), .O(n247) );
  NAND_GATE U693 ( .I1(n2055), .I2(n693), .O(n793) );
  NAND_GATE U694 ( .I1(n794), .I2(n695), .O(n792) );
  NAND_GATE U695 ( .I1(n2056), .I2(n697), .O(n791) );
  AND_GATE U699 ( .I1(n799), .I2(n800), .O(n248) );
  NAND_GATE U700 ( .I1(n697), .I2(n801), .O(n800) );
  NAND_GATE U701 ( .I1(n693), .I2(n802), .O(n799) );
  NAND4_GATE U709 ( .I1(n816), .I2(n817), .I3(n818), .I4(n819), .O(n467) );
  NAND_GATE U710 ( .I1(op2[19]), .I2(n396), .O(n819) );
  NAND_GATE U711 ( .I1(op2[20]), .I2(n397), .O(n818) );
  NAND_GATE U712 ( .I1(op2[21]), .I2(n398), .O(n817) );
  NAND_GATE U713 ( .I1(op2[22]), .I2(n399), .O(n816) );
  NAND_GATE U716 ( .I1(n820), .I2(n821), .O(n286) );
  NAND_GATE U717 ( .I1(n697), .I2(n822), .O(n821) );
  NAND_GATE U718 ( .I1(n693), .I2(n493), .O(n820) );
  NAND3_GATE U734 ( .I1(n833), .I2(n834), .I3(n835), .O(n280) );
  NAND_GATE U735 ( .I1(n2053), .I2(n693), .O(n835) );
  NAND_GATE U736 ( .I1(n695), .I2(n479), .O(n834) );
  NAND_GATE U737 ( .I1(n2054), .I2(n697), .O(n833) );
  AND3_GATE U741 ( .I1(n840), .I2(n841), .I3(n842), .O(n281) );
  NAND_GATE U742 ( .I1(n693), .I2(n843), .O(n842) );
  NAND_GATE U743 ( .I1(n695), .I2(n2038), .O(n841) );
  NAND_GATE U744 ( .I1(n697), .I2(n844), .O(n840) );
  NAND4_GATE U752 ( .I1(n858), .I2(n859), .I3(n860), .I4(n861), .O(n555) );
  NAND_GATE U753 ( .I1(op2[18]), .I2(n396), .O(n861) );
  NAND_GATE U754 ( .I1(op2[19]), .I2(n397), .O(n860) );
  NAND_GATE U755 ( .I1(op2[20]), .I2(n398), .O(n859) );
  NAND_GATE U756 ( .I1(op2[21]), .I2(n399), .O(n858) );
  NAND_GATE U759 ( .I1(n862), .I2(n863), .O(n316) );
  NAND_GATE U760 ( .I1(n697), .I2(n694), .O(n863) );
  NAND_GATE U761 ( .I1(n693), .I2(n696), .O(n862) );
  NAND3_GATE U777 ( .I1(n873), .I2(n874), .I3(n875), .O(n310) );
  NAND_GATE U778 ( .I1(n2057), .I2(n693), .O(n875) );
  NAND_GATE U779 ( .I1(n695), .I2(n562), .O(n874) );
  NAND_GATE U780 ( .I1(n697), .I2(n2029), .O(n873) );
  AND3_GATE U784 ( .I1(n880), .I2(n881), .I3(n882), .O(n311) );
  NAND_GATE U785 ( .I1(n693), .I2(n717), .O(n882) );
  NAND_GATE U786 ( .I1(n695), .I2(n563), .O(n881) );
  NAND_GATE U787 ( .I1(n697), .I2(n172), .O(n880) );
  NAND4_GATE U795 ( .I1(n896), .I2(n897), .I3(n898), .I4(n899), .O(n588) );
  NAND_GATE U796 ( .I1(op2[17]), .I2(n396), .O(n899) );
  NAND_GATE U797 ( .I1(op2[18]), .I2(n397), .O(n898) );
  NAND_GATE U798 ( .I1(op2[19]), .I2(n398), .O(n897) );
  NAND_GATE U799 ( .I1(op2[20]), .I2(n399), .O(n896) );
  NAND3_GATE U817 ( .I1(n909), .I2(n910), .I3(n911), .O(n340) );
  NAND_GATE U818 ( .I1(n2052), .I2(n693), .O(n911) );
  NAND_GATE U819 ( .I1(n2049), .I2(n695), .O(n910) );
  NAND_GATE U820 ( .I1(n2036), .I2(n697), .O(n909) );
  AND3_GATE U824 ( .I1(n916), .I2(n917), .I3(n918), .O(n341) );
  NAND_GATE U825 ( .I1(n693), .I2(n759), .O(n918) );
  NAND_GATE U826 ( .I1(n695), .I2(n760), .O(n917) );
  NAND_GATE U827 ( .I1(n697), .I2(n214), .O(n916) );
  NAND5_GATE U831 ( .I1(n919), .I2(n920), .I3(n921), .I4(n922), .I5(n923), .O(
        res[1]) );
  AND3_GATE U840 ( .I1(n931), .I2(n932), .I3(n933), .O(n922) );
  OR_GATE U850 ( .I1(n945), .I2(n114), .O(n934) );
  NAND_GATE U851 ( .I1(n6), .I2(n946), .O(n932) );
  NAND5_GATE U852 ( .I1(n947), .I2(n948), .I3(n949), .I4(n950), .I5(n951), .O(
        n946) );
  AND4_GATE U853 ( .I1(n952), .I2(n953), .I3(n954), .I4(n955), .O(n951) );
  NAND_GATE U854 ( .I1(n376), .I2(op2[4]), .O(n955) );
  NAND_GATE U855 ( .I1(n377), .I2(op2[3]), .O(n954) );
  NAND_GATE U856 ( .I1(n375), .I2(op2[2]), .O(n953) );
  NAND_GATE U857 ( .I1(n374), .I2(op2[1]), .O(n952) );
  NAND_GATE U858 ( .I1(n2026), .I2(n2046), .O(n950) );
  NAND_GATE U864 ( .I1(n2030), .I2(n2047), .O(n949) );
  NAND_GATE U865 ( .I1(n2027), .I2(n167), .O(n948) );
  NAND_GATE U871 ( .I1(n964), .I2(op1[4]), .O(n947) );
  NAND_GATE U872 ( .I1(hilo[1]), .I2(n178), .O(n931) );
  NAND_GATE U873 ( .I1(op2[1]), .I2(n965), .O(n921) );
  NAND_GATE U877 ( .I1(op1[1]), .I2(n967), .O(n919) );
  NAND4_GATE U884 ( .I1(n982), .I2(n983), .I3(n984), .I4(n985), .O(n430) );
  NAND_GATE U885 ( .I1(op2[16]), .I2(n396), .O(n985) );
  NAND_GATE U886 ( .I1(op2[17]), .I2(n397), .O(n984) );
  NAND_GATE U887 ( .I1(op2[18]), .I2(n398), .O(n983) );
  NAND_GATE U888 ( .I1(op2[19]), .I2(n399), .O(n982) );
  NAND3_GATE U906 ( .I1(n995), .I2(n996), .I3(n997), .O(n400) );
  NAND_GATE U907 ( .I1(op1[3]), .I2(n632), .O(n997) );
  NAND_GATE U908 ( .I1(n2040), .I2(n697), .O(n996) );
  NAND_GATE U909 ( .I1(n2056), .I2(n693), .O(n995) );
  AND3_GATE U913 ( .I1(n1002), .I2(n1003), .I3(n1004), .O(n379) );
  NAND_GATE U914 ( .I1(op1[3]), .I2(n1005), .O(n1004) );
  NAND_GATE U915 ( .I1(n697), .I2(n246), .O(n1003) );
  NAND_GATE U916 ( .I1(n693), .I2(n801), .O(n1002) );
  NAND4_GATE U924 ( .I1(n1020), .I2(n1021), .I3(n1022), .I4(n1023), .O(n468)
         );
  NAND_GATE U925 ( .I1(op2[15]), .I2(n396), .O(n1023) );
  NAND_GATE U926 ( .I1(op2[16]), .I2(n397), .O(n1022) );
  NAND_GATE U927 ( .I1(op2[17]), .I2(n398), .O(n1021) );
  NAND_GATE U928 ( .I1(op2[18]), .I2(n399), .O(n1020) );
  NAND4_GATE U946 ( .I1(n1033), .I2(n1034), .I3(n1035), .I4(n1036), .O(n522)
         );
  NAND_GATE U947 ( .I1(n1037), .I2(n479), .O(n1036) );
  NAND_GATE U948 ( .I1(n2053), .I2(n695), .O(n1035) );
  NAND_GATE U949 ( .I1(n2033), .I2(n697), .O(n1034) );
  NAND_GATE U950 ( .I1(n2054), .I2(n693), .O(n1033) );
  AND4_GATE U954 ( .I1(n1042), .I2(n1043), .I3(n1044), .I4(n1045), .O(n507) );
  NAND_GATE U955 ( .I1(n1037), .I2(n2038), .O(n1045) );
  NAND_GATE U956 ( .I1(n695), .I2(n843), .O(n1044) );
  NAND_GATE U957 ( .I1(n697), .I2(n279), .O(n1043) );
  NAND_GATE U958 ( .I1(n693), .I2(n844), .O(n1042) );
  NAND4_GATE U966 ( .I1(n1059), .I2(n1060), .I3(n1061), .I4(n1062), .O(n556)
         );
  NAND_GATE U967 ( .I1(op2[14]), .I2(n396), .O(n1062) );
  NAND_GATE U968 ( .I1(op2[15]), .I2(n397), .O(n1061) );
  NAND_GATE U969 ( .I1(op2[16]), .I2(n398), .O(n1060) );
  NAND_GATE U970 ( .I1(op2[17]), .I2(n399), .O(n1059) );
  NAND4_GATE U988 ( .I1(n1072), .I2(n1073), .I3(n1074), .I4(n1075), .O(n964)
         );
  NAND_GATE U989 ( .I1(n1037), .I2(n562), .O(n1075) );
  NAND_GATE U990 ( .I1(n695), .I2(n2057), .O(n1074) );
  NAND_GATE U991 ( .I1(n697), .I2(n2028), .O(n1073) );
  NAND_GATE U992 ( .I1(n693), .I2(n2029), .O(n1072) );
  AND4_GATE U996 ( .I1(n1080), .I2(n1081), .I3(n1082), .I4(n1083), .O(n945) );
  NAND_GATE U997 ( .I1(n1037), .I2(n563), .O(n1083) );
  NAND_GATE U998 ( .I1(n695), .I2(n717), .O(n1082) );
  NAND_GATE U999 ( .I1(n697), .I2(n170), .O(n1081) );
  NAND_GATE U1000 ( .I1(n693), .I2(n172), .O(n1080) );
  NAND4_GATE U1012 ( .I1(n1096), .I2(n1097), .I3(n1098), .I4(n1099), .O(n589)
         );
  NAND_GATE U1013 ( .I1(op2[13]), .I2(n396), .O(n1099) );
  NAND_GATE U1014 ( .I1(op2[14]), .I2(n397), .O(n1098) );
  NAND_GATE U1015 ( .I1(op2[15]), .I2(n398), .O(n1097) );
  NAND_GATE U1016 ( .I1(op2[16]), .I2(n399), .O(n1096) );
  NAND_GATE U1054 ( .I1(n1037), .I2(n361), .O(n1132) );
  NAND_GATE U1055 ( .I1(n695), .I2(n780), .O(n1131) );
  NAND_GATE U1056 ( .I1(n697), .I2(n619), .O(n1130) );
  NAND4_GATE U1057 ( .I1(n1133), .I2(n1134), .I3(n1135), .I4(n1136), .O(n619)
         );
  NAND_GATE U1058 ( .I1(op2[12]), .I2(n396), .O(n1136) );
  NAND_GATE U1059 ( .I1(op2[13]), .I2(n397), .O(n1135) );
  NAND_GATE U1060 ( .I1(op2[14]), .I2(n398), .O(n1134) );
  NAND_GATE U1061 ( .I1(op2[15]), .I2(n399), .O(n1133) );
  NAND_GATE U1062 ( .I1(n693), .I2(n781), .O(n1129) );
  NAND4_GATE U1071 ( .I1(n1146), .I2(n1147), .I3(n1148), .I4(n1149), .O(n1145)
         );
  NAND_GATE U1072 ( .I1(n2056), .I2(n2046), .O(n1149) );
  NAND_GATE U1073 ( .I1(n2055), .I2(n2047), .O(n1148) );
  NAND_GATE U1074 ( .I1(n2040), .I2(n167), .O(n1147) );
  NAND_GATE U1075 ( .I1(n2039), .I2(n175), .O(n1146) );
  NAND5_GATE U1095 ( .I1(n1167), .I2(n1168), .I3(n1169), .I4(n1170), .I5(n1171), .O(n1166) );
  NAND_GATE U1096 ( .I1(n1172), .I2(n2051), .O(n1171) );
  NAND3_GATE U1097 ( .I1(n1173), .I2(n1174), .I3(n1175), .O(n1172) );
  NAND_GATE U1098 ( .I1(n2033), .I2(n693), .O(n1175) );
  NAND_GATE U1099 ( .I1(n1037), .I2(n2053), .O(n1174) );
  NAND_GATE U1100 ( .I1(n2054), .I2(n695), .O(n1173) );
  OR_GATE U1101 ( .I1(n2050), .I2(n2038), .O(n1170) );
  NAND_GATE U1102 ( .I1(n2032), .I2(n175), .O(n1169) );
  NAND_GATE U1103 ( .I1(n11), .I2(n479), .O(n1167) );
  NAND_GATE U1115 ( .I1(n1037), .I2(n493), .O(n1186) );
  NAND_GATE U1116 ( .I1(n695), .I2(n822), .O(n1185) );
  NAND_GATE U1117 ( .I1(n697), .I2(n657), .O(n1184) );
  NAND4_GATE U1118 ( .I1(n1187), .I2(n1188), .I3(n1189), .I4(n1190), .O(n657)
         );
  NAND_GATE U1119 ( .I1(op2[11]), .I2(n396), .O(n1190) );
  NAND_GATE U1120 ( .I1(op2[12]), .I2(n397), .O(n1189) );
  NAND_GATE U1121 ( .I1(op2[13]), .I2(n398), .O(n1188) );
  NAND_GATE U1122 ( .I1(op2[14]), .I2(n399), .O(n1187) );
  NAND_GATE U1123 ( .I1(n693), .I2(n823), .O(n1183) );
  NAND5_GATE U1134 ( .I1(n1204), .I2(n1168), .I3(n1205), .I4(n1206), .I5(n1207), .O(n1203) );
  NAND_GATE U1135 ( .I1(n1208), .I2(n2051), .O(n1207) );
  NAND3_GATE U1136 ( .I1(n1209), .I2(n1210), .I3(n1211), .O(n1208) );
  NAND_GATE U1137 ( .I1(n693), .I2(n2028), .O(n1211) );
  NAND_GATE U1143 ( .I1(n1037), .I2(n2057), .O(n1210) );
  NAND4_GATE U1144 ( .I1(n1216), .I2(n1217), .I3(n1218), .I4(n1219), .O(n717)
         );
  NAND_GATE U1145 ( .I1(n396), .I2(n106), .O(n1219) );
  NAND_GATE U1146 ( .I1(n397), .I2(n105), .O(n1218) );
  NAND_GATE U1147 ( .I1(n398), .I2(n104), .O(n1217) );
  NAND_GATE U1148 ( .I1(n399), .I2(n103), .O(n1216) );
  NAND_GATE U1149 ( .I1(n695), .I2(n2029), .O(n1209) );
  NAND_GATE U1151 ( .I1(n396), .I2(n102), .O(n1223) );
  NAND_GATE U1152 ( .I1(n397), .I2(n101), .O(n1222) );
  NAND_GATE U1153 ( .I1(n398), .I2(n100), .O(n1221) );
  OR_GATE U1155 ( .I1(n563), .I2(n2050), .O(n1206) );
  NAND_GATE U1157 ( .I1(n398), .I2(n108), .O(n1225) );
  NAND_GATE U1158 ( .I1(n399), .I2(n107), .O(n1224) );
  NAND_GATE U1159 ( .I1(n175), .I2(n2030), .O(n1205) );
  NAND_GATE U1165 ( .I1(n11), .I2(n562), .O(n1204) );
  NAND3_GATE U1166 ( .I1(n1230), .I2(n1231), .I3(n1232), .O(n562) );
  NAND_GATE U1167 ( .I1(op2[29]), .I2(n399), .O(n1232) );
  NAND_GATE U1168 ( .I1(op2[31]), .I2(n397), .O(n1231) );
  NAND_GATE U1169 ( .I1(op2[30]), .I2(n398), .O(n1230) );
  NAND_GATE U1181 ( .I1(n1037), .I2(n696), .O(n1243) );
  NAND_GATE U1182 ( .I1(n1244), .I2(n1245), .O(n696) );
  NAND_GATE U1183 ( .I1(op2[0]), .I2(n398), .O(n1245) );
  NAND_GATE U1184 ( .I1(op2[1]), .I2(n399), .O(n1244) );
  NAND_GATE U1185 ( .I1(n695), .I2(n694), .O(n1242) );
  NAND4_GATE U1186 ( .I1(n1246), .I2(n1247), .I3(n1248), .I4(n1249), .O(n694)
         );
  NAND_GATE U1187 ( .I1(op2[2]), .I2(n396), .O(n1249) );
  NAND_GATE U1188 ( .I1(op2[3]), .I2(n397), .O(n1248) );
  NAND_GATE U1189 ( .I1(op2[4]), .I2(n398), .O(n1247) );
  NAND_GATE U1190 ( .I1(op2[5]), .I2(n399), .O(n1246) );
  NAND_GATE U1191 ( .I1(n697), .I2(n699), .O(n1241) );
  NAND4_GATE U1192 ( .I1(n1250), .I2(n1251), .I3(n1252), .I4(n1253), .O(n699)
         );
  NAND_GATE U1193 ( .I1(op2[10]), .I2(n396), .O(n1253) );
  NAND_GATE U1194 ( .I1(op2[11]), .I2(n397), .O(n1252) );
  NAND_GATE U1195 ( .I1(op2[12]), .I2(n398), .O(n1251) );
  NAND_GATE U1196 ( .I1(op2[13]), .I2(n399), .O(n1250) );
  NAND_GATE U1197 ( .I1(n693), .I2(n698), .O(n1240) );
  NAND4_GATE U1198 ( .I1(n1254), .I2(n1255), .I3(n1256), .I4(n1257), .O(n698)
         );
  NAND_GATE U1199 ( .I1(op2[6]), .I2(n396), .O(n1257) );
  NAND_GATE U1200 ( .I1(op2[7]), .I2(n397), .O(n1256) );
  NAND_GATE U1201 ( .I1(op2[8]), .I2(n398), .O(n1255) );
  NAND_GATE U1202 ( .I1(n399), .I2(op2[9]), .O(n1254) );
  NAND_GATE U1213 ( .I1(op1[3]), .I2(n327), .O(n1272) );
  NAND_GATE U1214 ( .I1(n1273), .I2(n1274), .O(n327) );
  NAND_GATE U1215 ( .I1(n53), .I2(op1[2]), .O(n1274) );
  NAND_GATE U1216 ( .I1(n738), .I2(n112), .O(n1273) );
  NAND4_GATE U1217 ( .I1(n1275), .I2(n1276), .I3(n1277), .I4(n1278), .O(n738)
         );
  NAND_GATE U1218 ( .I1(op2[1]), .I2(n396), .O(n1278) );
  NAND_GATE U1219 ( .I1(op2[2]), .I2(n397), .O(n1277) );
  NAND_GATE U1220 ( .I1(op2[3]), .I2(n398), .O(n1276) );
  NAND_GATE U1221 ( .I1(op2[4]), .I2(n399), .O(n1275) );
  NAND_GATE U1222 ( .I1(n697), .I2(n741), .O(n1271) );
  NAND4_GATE U1223 ( .I1(n1279), .I2(n1280), .I3(n1281), .I4(n1282), .O(n741)
         );
  NAND_GATE U1224 ( .I1(n396), .I2(op2[9]), .O(n1282) );
  NAND_GATE U1225 ( .I1(op2[10]), .I2(n397), .O(n1281) );
  NAND_GATE U1226 ( .I1(op2[11]), .I2(n398), .O(n1280) );
  NAND_GATE U1227 ( .I1(op2[12]), .I2(n399), .O(n1279) );
  NAND_GATE U1228 ( .I1(n693), .I2(n740), .O(n1270) );
  NAND4_GATE U1229 ( .I1(n1283), .I2(n1284), .I3(n1285), .I4(n1286), .O(n740)
         );
  NAND_GATE U1230 ( .I1(op2[5]), .I2(n396), .O(n1286) );
  NAND_GATE U1231 ( .I1(op2[6]), .I2(n397), .O(n1285) );
  NAND_GATE U1232 ( .I1(op2[7]), .I2(n398), .O(n1284) );
  NAND_GATE U1233 ( .I1(op2[8]), .I2(n399), .O(n1283) );
  NAND_GATE U1237 ( .I1(n2049), .I2(n1291), .O(n1290) );
  OR_GATE U1238 ( .I1(n2042), .I2(n11), .O(n1291) );
  NAND3_GATE U1242 ( .I1(n1293), .I2(n1294), .I3(n1295), .O(n1292) );
  NAND_GATE U1243 ( .I1(n2035), .I2(n693), .O(n1295) );
  NAND_GATE U1244 ( .I1(n1037), .I2(n2052), .O(n1294) );
  NAND_GATE U1245 ( .I1(n2036), .I2(n695), .O(n1293) );
  NAND5_GATE U1266 ( .I1(n1319), .I2(n1320), .I3(n1321), .I4(n1322), .I5(n1323), .O(n1318) );
  NAND_GATE U1267 ( .I1(n2031), .I2(n175), .O(n1323) );
  NAND_GATE U1273 ( .I1(n2042), .I2(n631), .O(n1322) );
  NAND_GATE U1274 ( .I1(n113), .I2(n1005), .O(n631) );
  NOR_GATE U1275 ( .I1(n2055), .I2(op1[2]), .O(n1005) );
  NAND_GATE U1276 ( .I1(n1328), .I2(n2051), .O(n1321) );
  NAND_GATE U1277 ( .I1(n1329), .I2(n1330), .O(n1328) );
  NAND_GATE U1278 ( .I1(n1037), .I2(n2056), .O(n1330) );
  NAND4_GATE U1279 ( .I1(n1331), .I2(n1332), .I3(n1333), .I4(n1334), .O(n801)
         );
  NAND_GATE U1280 ( .I1(n396), .I2(n104), .O(n1334) );
  NAND_GATE U1281 ( .I1(n397), .I2(n103), .O(n1333) );
  NAND_GATE U1282 ( .I1(n398), .I2(n102), .O(n1332) );
  NAND_GATE U1283 ( .I1(n399), .I2(n101), .O(n1331) );
  NAND_GATE U1284 ( .I1(n2040), .I2(n695), .O(n1329) );
  NAND_GATE U1286 ( .I1(n396), .I2(n100), .O(n1338) );
  NAND_GATE U1290 ( .I1(n2039), .I2(n167), .O(n1320) );
  NAND3_GATE U1296 ( .I1(n632), .I2(n113), .I3(n2041), .O(n1319) );
  NAND_GATE U1297 ( .I1(n1343), .I2(n1344), .O(n632) );
  NAND_GATE U1298 ( .I1(n794), .I2(op1[2]), .O(n1344) );
  AND_GATE U1299 ( .I1(op2[31]), .I2(n399), .O(n794) );
  NAND_GATE U1300 ( .I1(n2055), .I2(n112), .O(n1343) );
  NAND4_GATE U1301 ( .I1(n1345), .I2(n1346), .I3(n1347), .I4(n1348), .O(n802)
         );
  NAND_GATE U1302 ( .I1(n396), .I2(n108), .O(n1348) );
  NAND_GATE U1303 ( .I1(n397), .I2(n107), .O(n1347) );
  NAND_GATE U1304 ( .I1(n398), .I2(n106), .O(n1346) );
  NAND_GATE U1305 ( .I1(n399), .I2(n105), .O(n1345) );
  NAND_GATE U1317 ( .I1(n693), .I2(n780), .O(n1355) );
  NAND4_GATE U1318 ( .I1(n1356), .I2(n1357), .I3(n1358), .I4(n1359), .O(n780)
         );
  NAND_GATE U1319 ( .I1(op2[4]), .I2(n396), .O(n1359) );
  NAND_GATE U1320 ( .I1(op2[5]), .I2(n397), .O(n1358) );
  NAND_GATE U1321 ( .I1(op2[6]), .I2(n398), .O(n1357) );
  NAND_GATE U1322 ( .I1(op2[7]), .I2(n399), .O(n1356) );
  NAND_GATE U1323 ( .I1(n695), .I2(n361), .O(n1354) );
  NAND4_GATE U1324 ( .I1(n1360), .I2(n1361), .I3(n1362), .I4(n1363), .O(n361)
         );
  NAND_GATE U1325 ( .I1(op2[0]), .I2(n396), .O(n1363) );
  NAND_GATE U1326 ( .I1(op2[1]), .I2(n397), .O(n1362) );
  NAND_GATE U1327 ( .I1(op2[2]), .I2(n398), .O(n1361) );
  NAND_GATE U1328 ( .I1(op2[3]), .I2(n399), .O(n1360) );
  NAND_GATE U1329 ( .I1(n697), .I2(n781), .O(n1353) );
  NAND4_GATE U1330 ( .I1(n1364), .I2(n1365), .I3(n1366), .I4(n1367), .O(n781)
         );
  NAND_GATE U1331 ( .I1(op2[8]), .I2(n396), .O(n1367) );
  NAND_GATE U1332 ( .I1(n397), .I2(op2[9]), .O(n1366) );
  NAND_GATE U1333 ( .I1(op2[10]), .I2(n398), .O(n1365) );
  NAND_GATE U1334 ( .I1(op2[11]), .I2(n399), .O(n1364) );
  NAND4_GATE U1345 ( .I1(n1384), .I2(n1385), .I3(n1386), .I4(n1387), .O(n1383)
         );
  AND3_GATE U1346 ( .I1(n1388), .I2(n1389), .I3(n1390), .O(n1387) );
  NAND_GATE U1347 ( .I1(n2032), .I2(n167), .O(n1390) );
  NAND_GATE U1353 ( .I1(n2033), .I2(n2046), .O(n1389) );
  NAND_GATE U1359 ( .I1(n2054), .I2(n2047), .O(n1388) );
  NAND4_GATE U1360 ( .I1(n1399), .I2(n1400), .I3(n1401), .I4(n1402), .O(n844)
         );
  NAND_GATE U1361 ( .I1(n396), .I2(n103), .O(n1402) );
  NAND_GATE U1362 ( .I1(n397), .I2(n102), .O(n1401) );
  NAND_GATE U1363 ( .I1(n398), .I2(n101), .O(n1400) );
  NAND_GATE U1364 ( .I1(n399), .I2(n100), .O(n1399) );
  NAND_GATE U1365 ( .I1(n2041), .I2(n667), .O(n1386) );
  NAND_GATE U1366 ( .I1(n1403), .I2(n1404), .O(n667) );
  NAND_GATE U1367 ( .I1(n2053), .I2(n697), .O(n1404) );
  NAND_GATE U1368 ( .I1(n693), .I2(n479), .O(n1403) );
  NAND_GATE U1369 ( .I1(n1405), .I2(n1406), .O(n479) );
  NAND_GATE U1370 ( .I1(op2[31]), .I2(n398), .O(n1406) );
  NAND_GATE U1371 ( .I1(op2[30]), .I2(n399), .O(n1405) );
  NAND_GATE U1373 ( .I1(n2034), .I2(n175), .O(n1385) );
  NAND_GATE U1379 ( .I1(n672), .I2(n2042), .O(n1384) );
  AND_GATE U1381 ( .I1(n1411), .I2(n1412), .O(n672) );
  NAND_GATE U1382 ( .I1(n697), .I2(n843), .O(n1412) );
  NAND4_GATE U1383 ( .I1(n1413), .I2(n1414), .I3(n1415), .I4(n1416), .O(n843)
         );
  NAND_GATE U1384 ( .I1(n396), .I2(n107), .O(n1416) );
  NAND_GATE U1385 ( .I1(n397), .I2(n106), .O(n1415) );
  NAND_GATE U1386 ( .I1(n398), .I2(n105), .O(n1414) );
  NAND_GATE U1387 ( .I1(n399), .I2(n104), .O(n1413) );
  NAND_GATE U1388 ( .I1(n693), .I2(n2038), .O(n1411) );
  NAND_GATE U1402 ( .I1(n693), .I2(n822), .O(n1424) );
  NAND4_GATE U1403 ( .I1(n1425), .I2(n1426), .I3(n1427), .I4(n1428), .O(n822)
         );
  NAND_GATE U1404 ( .I1(op2[3]), .I2(n396), .O(n1428) );
  NAND_GATE U1405 ( .I1(op2[4]), .I2(n397), .O(n1427) );
  NAND_GATE U1406 ( .I1(op2[5]), .I2(n398), .O(n1426) );
  NAND_GATE U1407 ( .I1(op2[6]), .I2(n399), .O(n1425) );
  NAND_GATE U1408 ( .I1(n695), .I2(n493), .O(n1423) );
  NAND3_GATE U1409 ( .I1(n1429), .I2(n1430), .I3(n1431), .O(n493) );
  NAND_GATE U1410 ( .I1(op2[2]), .I2(n399), .O(n1431) );
  NAND_GATE U1411 ( .I1(op2[0]), .I2(n397), .O(n1430) );
  NAND_GATE U1412 ( .I1(op2[1]), .I2(n398), .O(n1429) );
  NAND_GATE U1413 ( .I1(n697), .I2(n823), .O(n1422) );
  NAND4_GATE U1414 ( .I1(n1432), .I2(n1433), .I3(n1434), .I4(n1435), .O(n823)
         );
  NAND_GATE U1415 ( .I1(op2[7]), .I2(n396), .O(n1435) );
  NAND_GATE U1416 ( .I1(op2[8]), .I2(n397), .O(n1434) );
  NAND_GATE U1417 ( .I1(n398), .I2(op2[9]), .O(n1433) );
  NAND_GATE U1418 ( .I1(op2[10]), .I2(n399), .O(n1432) );
  NAND_GATE U1433 ( .I1(n1457), .I2(op1[4]), .O(n1446) );
  NAND5_GATE U1439 ( .I1(n1465), .I2(n1466), .I3(n1467), .I4(n1468), .I5(n1469), .O(n1464) );
  AND4_GATE U1440 ( .I1(n1470), .I2(n1471), .I3(n1472), .I4(n1473), .O(n1469)
         );
  NAND_GATE U1441 ( .I1(n376), .I2(op2[3]), .O(n1473) );
  AND_GATE U1442 ( .I1(n175), .I2(n396), .O(n376) );
  NAND_GATE U1443 ( .I1(n377), .I2(op2[2]), .O(n1472) );
  AND_GATE U1444 ( .I1(n175), .I2(n397), .O(n377) );
  NAND_GATE U1445 ( .I1(n375), .I2(op2[1]), .O(n1471) );
  AND_GATE U1446 ( .I1(n175), .I2(n398), .O(n375) );
  NAND_GATE U1447 ( .I1(n374), .I2(op2[0]), .O(n1470) );
  AND_GATE U1448 ( .I1(n175), .I2(n399), .O(n374) );
  NAND_GATE U1449 ( .I1(n2045), .I2(n2046), .O(n1468) );
  NAND_GATE U1450 ( .I1(n1474), .I2(n112), .O(n169) );
  NAND_GATE U1456 ( .I1(n2043), .I2(n2047), .O(n1467) );
  NAND_GATE U1457 ( .I1(op1[2]), .I2(n1474), .O(n171) );
  NOR_GATE U1458 ( .I1(n113), .I2(op1[4]), .O(n1474) );
  NAND_GATE U1464 ( .I1(n2044), .I2(n167), .O(n1466) );
  AND_GATE U1465 ( .I1(n693), .I2(n114), .O(n167) );
  NAND_GATE U1471 ( .I1(n2048), .I2(op1[4]), .O(n1465) );
  NAND4_GATE U1472 ( .I1(n1487), .I2(n1488), .I3(n1489), .I4(n1490), .O(n1457)
         );
  NAND_GATE U1473 ( .I1(n1037), .I2(n760), .O(n1490) );
  NAND4_GATE U1474 ( .I1(n1491), .I2(n1492), .I3(n1493), .I4(n1494), .O(n760)
         );
  NAND_GATE U1475 ( .I1(n396), .I2(n109), .O(n1494) );
  NAND_GATE U1476 ( .I1(n397), .I2(n108), .O(n1493) );
  NAND_GATE U1477 ( .I1(n398), .I2(n107), .O(n1492) );
  NAND_GATE U1478 ( .I1(n399), .I2(n106), .O(n1491) );
  NOR_GATE U1479 ( .I1(n112), .I2(n113), .O(n1037) );
  NAND_GATE U1480 ( .I1(n695), .I2(n759), .O(n1489) );
  NAND4_GATE U1481 ( .I1(n1495), .I2(n1496), .I3(n1497), .I4(n1498), .O(n759)
         );
  NAND_GATE U1482 ( .I1(n396), .I2(n105), .O(n1498) );
  NAND_GATE U1483 ( .I1(n397), .I2(n104), .O(n1497) );
  NAND_GATE U1484 ( .I1(n398), .I2(n103), .O(n1496) );
  NAND_GATE U1485 ( .I1(n399), .I2(n102), .O(n1495) );
  NOR_GATE U1486 ( .I1(n113), .I2(op1[2]), .O(n695) );
  OR_GATE U1487 ( .I1(n76), .I2(n2035), .O(n1488) );
  NAND_GATE U1493 ( .I1(n693), .I2(n214), .O(n1487) );
  NAND_GATE U1495 ( .I1(n396), .I2(n101), .O(n1506) );
  NOR_GATE U1496 ( .I1(n111), .I2(n110), .O(n396) );
  NAND_GATE U1497 ( .I1(n397), .I2(n100), .O(n1505) );
  NOR_GATE U1498 ( .I1(n111), .I2(op1[0]), .O(n397) );
  NOR_GATE U1500 ( .I1(n110), .I2(op1[1]), .O(n398) );
  NOR_GATE U1502 ( .I1(n112), .I2(op1[3]), .O(n693) );
  NOR_GATE U1514 ( .I1(op1[1]), .I2(op1[0]), .O(n399) );
  AND_GATE U1516 ( .I1(n697), .I2(n114), .O(n175) );
  AND_GATE U1517 ( .I1(n113), .I2(n112), .O(n697) );
  NAND4_GATE U1814 ( .I1(n1774), .I2(n1775), .I3(n1776), .I4(n1777), .O(n1978)
         );
  NAND_GATE U1815 ( .I1(N786), .I2(n9), .O(n1777) );
  NAND_GATE U1816 ( .I1(n2037), .I2(op1[11]), .O(n1776) );
  NAND_GATE U1817 ( .I1(N721), .I2(n10), .O(n1775) );
  NAND_GATE U1818 ( .I1(hilo[11]), .I2(n1697), .O(n1774) );
  NAND4_GATE U1819 ( .I1(n1778), .I2(n1779), .I3(n1780), .I4(n1781), .O(n1979)
         );
  NAND_GATE U1820 ( .I1(N785), .I2(n9), .O(n1781) );
  NAND_GATE U1821 ( .I1(n2037), .I2(op1[10]), .O(n1780) );
  NAND_GATE U1822 ( .I1(N720), .I2(n10), .O(n1779) );
  NAND_GATE U1823 ( .I1(hilo[10]), .I2(n1697), .O(n1778) );
  NAND4_GATE U1824 ( .I1(n1782), .I2(n1783), .I3(n1784), .I4(n1785), .O(n1980)
         );
  NAND_GATE U1825 ( .I1(N784), .I2(n9), .O(n1785) );
  NAND_GATE U1826 ( .I1(n2037), .I2(op1[9]), .O(n1784) );
  NAND_GATE U1827 ( .I1(N719), .I2(n10), .O(n1783) );
  NAND_GATE U1828 ( .I1(hilo[9]), .I2(n1697), .O(n1782) );
  NAND4_GATE U1829 ( .I1(n1786), .I2(n1787), .I3(n1788), .I4(n1789), .O(n1981)
         );
  NAND_GATE U1830 ( .I1(N783), .I2(n9), .O(n1789) );
  NAND_GATE U1831 ( .I1(n2037), .I2(op1[8]), .O(n1788) );
  NAND_GATE U1832 ( .I1(N718), .I2(n10), .O(n1787) );
  NAND_GATE U1833 ( .I1(hilo[8]), .I2(n1697), .O(n1786) );
  NAND4_GATE U1834 ( .I1(n1790), .I2(n1791), .I3(n1792), .I4(n1793), .O(n1982)
         );
  NAND_GATE U1835 ( .I1(N782), .I2(n9), .O(n1793) );
  NAND_GATE U1836 ( .I1(n2037), .I2(op1[7]), .O(n1792) );
  NAND_GATE U1837 ( .I1(N717), .I2(n10), .O(n1791) );
  NAND_GATE U1838 ( .I1(hilo[7]), .I2(n1697), .O(n1790) );
  NAND4_GATE U1839 ( .I1(n1794), .I2(n1795), .I3(n1796), .I4(n1797), .O(n1983)
         );
  NAND_GATE U1840 ( .I1(N781), .I2(n9), .O(n1797) );
  NAND_GATE U1841 ( .I1(n2037), .I2(op1[6]), .O(n1796) );
  NAND_GATE U1842 ( .I1(N716), .I2(n10), .O(n1795) );
  NAND_GATE U1843 ( .I1(hilo[6]), .I2(n1697), .O(n1794) );
  NAND4_GATE U1844 ( .I1(n1798), .I2(n1799), .I3(n1800), .I4(n1801), .O(n1984)
         );
  NAND_GATE U1845 ( .I1(N780), .I2(n9), .O(n1801) );
  NAND_GATE U1846 ( .I1(n2037), .I2(op1[5]), .O(n1800) );
  NAND_GATE U1847 ( .I1(N715), .I2(n10), .O(n1799) );
  NAND_GATE U1848 ( .I1(hilo[5]), .I2(n1697), .O(n1798) );
  NAND4_GATE U1849 ( .I1(n1802), .I2(n1803), .I3(n1804), .I4(n1805), .O(n1985)
         );
  NAND_GATE U1850 ( .I1(N779), .I2(n9), .O(n1805) );
  NAND_GATE U1851 ( .I1(n2037), .I2(op1[4]), .O(n1804) );
  NAND_GATE U1852 ( .I1(N714), .I2(n10), .O(n1803) );
  NAND_GATE U1853 ( .I1(hilo[4]), .I2(n1697), .O(n1802) );
  NAND4_GATE U1854 ( .I1(n1806), .I2(n1807), .I3(n1808), .I4(n1809), .O(n1986)
         );
  NAND_GATE U1855 ( .I1(N778), .I2(n9), .O(n1809) );
  NAND_GATE U1856 ( .I1(n2037), .I2(op1[3]), .O(n1808) );
  NAND_GATE U1857 ( .I1(N713), .I2(n10), .O(n1807) );
  NAND_GATE U1858 ( .I1(hilo[3]), .I2(n1697), .O(n1806) );
  NAND4_GATE U1859 ( .I1(n1810), .I2(n1811), .I3(n1812), .I4(n1813), .O(n1987)
         );
  NAND_GATE U1860 ( .I1(N777), .I2(n9), .O(n1813) );
  NAND_GATE U1861 ( .I1(n2037), .I2(op1[2]), .O(n1812) );
  NAND_GATE U1862 ( .I1(N712), .I2(n10), .O(n1811) );
  NAND_GATE U1863 ( .I1(hilo[2]), .I2(n1697), .O(n1810) );
  NAND4_GATE U1864 ( .I1(n1814), .I2(n1815), .I3(n1816), .I4(n1817), .O(n1988)
         );
  NAND_GATE U1865 ( .I1(N776), .I2(n9), .O(n1817) );
  NAND_GATE U1866 ( .I1(n2037), .I2(op1[1]), .O(n1816) );
  NAND_GATE U1867 ( .I1(N711), .I2(n10), .O(n1815) );
  NAND_GATE U1868 ( .I1(hilo[1]), .I2(n1697), .O(n1814) );
  NAND4_GATE U1869 ( .I1(n1818), .I2(n1819), .I3(n1820), .I4(n1821), .O(n1989)
         );
  NAND_GATE U1870 ( .I1(N775), .I2(n9), .O(n1821) );
  NAND_GATE U1872 ( .I1(n2037), .I2(op1[0]), .O(n1820) );
  NAND_GATE U1874 ( .I1(N710), .I2(n10), .O(n1819) );
  NAND_GATE U1876 ( .I1(hilo[0]), .I2(n1697), .O(n1818) );
  NAND_GATE U2001 ( .I1(n1910), .I2(n1911), .O(n1909) );
  NAND_GATE U2002 ( .I1(op1[31]), .I2(efct_op2[31]), .O(n1911) );
  NAND_GATE U2003 ( .I1(n2058), .I2(n141), .O(n1910) );
  NAND_GATE U2042 ( .I1(n1922), .I2(n1923), .O(n417) );
  NAND_GATE U2043 ( .I1(op2[31]), .I2(n141), .O(n1923) );
  NAND_GATE U2044 ( .I1(op1[31]), .I2(n109), .O(n1922) );
  alu_DW01_add_0 add_1_root_add_125_2 ( .A({\efct_op1[32] , op1}), .B(efct_op2), .CI(n77), .SUM(res_add) );
  alu_DW02_mult_1 mult_138_2 ( .A(op1), .B(op2), .TC(1'b0), .PRODUCT({N838, 
        N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, 
        N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, 
        N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, 
        N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, 
        N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, 
        N777, N776, N775}) );
  alu_DW02_mult_0 mult_138 ( .A(op1), .B(op2), .TC(1'b1), .PRODUCT({N773, N772, 
        N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, 
        N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, 
        N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, 
        N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, 
        N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, 
        N711, N710}) );
  NAND_GATE U2 ( .I1(n402), .I2(n4), .O(n1) );
  NAND_GATE U3 ( .I1(n1), .I2(n2), .O(n570) );
  OR_GATE U4 ( .I1(n3), .I2(n404), .O(n2) );
  INV_GATE U5 ( .I1(n439), .O(n3) );
  AND_GATE U6 ( .I1(n395), .I2(n439), .O(n4) );
  AND_GATE U7 ( .I1(n8), .I2(n1839), .O(n5) );
  AND_GATE U8 ( .I1(n1512), .I2(n1701), .O(n6) );
  AND_GATE U9 ( .I1(n327), .I2(n113), .O(n7) );
  NOR_GATE U10 ( .I1(n1521), .I2(reset), .O(n8) );
  AND_GATE U11 ( .I1(n1526), .I2(n5), .O(n9) );
  NOR_GATE U12 ( .I1(n1523), .I2(reset), .O(n10) );
  AND_GATE U13 ( .I1(n697), .I2(n2041), .O(n11) );
  AND_GATE U14 ( .I1(n1688), .I2(n1696), .O(n12) );
  AND_GATE U15 ( .I1(n175), .I2(n1507), .O(n13) );
  AND_GATE U16 ( .I1(n2047), .I2(n1507), .O(n14) );
  AND_GATE U17 ( .I1(n167), .I2(n1507), .O(n15) );
  AND_GATE U18 ( .I1(n697), .I2(n51), .O(n16) );
  AND_GATE U19 ( .I1(n2046), .I2(n1507), .O(n17) );
  NAND_GATE U20 ( .I1(n458), .I2(n21), .O(n18) );
  AND_GATE U21 ( .I1(n18), .I2(n19), .O(n569) );
  OR_GATE U22 ( .I1(n20), .I2(n473), .O(n19) );
  INV_GATE U23 ( .I1(n49), .O(n20) );
  AND_GATE U24 ( .I1(n470), .I2(n49), .O(n21) );
  OR3_GATE U25 ( .I1(n22), .I2(n23), .I3(n27), .O(n1941) );
  AND_GATE U26 ( .I1(N823), .I2(n9), .O(n22) );
  AND_GATE U27 ( .I1(N758), .I2(n10), .O(n23) );
  OR3_GATE U28 ( .I1(n24), .I2(n25), .I3(n26), .O(n1926) );
  AND_GATE U29 ( .I1(N838), .I2(n9), .O(n24) );
  AND_GATE U30 ( .I1(N773), .I2(n10), .O(n25) );
  NAND_GATE U31 ( .I1(n2023), .I2(n2022), .O(n26) );
  NAND_GATE U32 ( .I1(n1902), .I2(n1901), .O(n27) );
  AND_GATE U33 ( .I1(n47), .I2(n29), .O(n28) );
  AND_GATE U34 ( .I1(n46), .I2(n41), .O(n29) );
  AND_GATE U35 ( .I1(n47), .I2(n48), .O(n30) );
  AND_GATE U36 ( .I1(n48), .I2(n29), .O(n31) );
  AND_GATE U37 ( .I1(n50), .I2(n44), .O(n32) );
  OR3_GATE U38 ( .I1(n33), .I2(n34), .I3(n72), .O(n1933) );
  AND_GATE U39 ( .I1(N766), .I2(n10), .O(n33) );
  AND_GATE U40 ( .I1(N831), .I2(n9), .O(n34) );
  OR3_GATE U41 ( .I1(n35), .I2(n36), .I3(n69), .O(n1927) );
  AND_GATE U42 ( .I1(N837), .I2(n9), .O(n35) );
  AND_GATE U43 ( .I1(N772), .I2(n10), .O(n36) );
  OR3_GATE U44 ( .I1(n37), .I2(n38), .I3(n73), .O(n1948) );
  AND_GATE U45 ( .I1(N816), .I2(n9), .O(n37) );
  AND_GATE U46 ( .I1(N751), .I2(n10), .O(n38) );
  AND_GATE U47 ( .I1(n143), .I2(n28), .O(n39) );
  AND_GATE U48 ( .I1(n527), .I2(n55), .O(n40) );
  AND_GATE U49 ( .I1(n153), .I2(n43), .O(n41) );
  AND_GATE U50 ( .I1(n145), .I2(n40), .O(n42) );
  AND3_GATE U51 ( .I1(n57), .I2(n44), .I3(n154), .O(n43) );
  AND_GATE U52 ( .I1(n455), .I2(n56), .O(n44) );
  OR_GATE U53 ( .I1(n45), .I2(n546), .O(n560) );
  INV_GATE U54 ( .I1(n545), .O(n45) );
  AND3_GATE U55 ( .I1(n486), .I2(n58), .I3(n59), .O(n46) );
  AND_GATE U56 ( .I1(n61), .I2(n60), .O(n47) );
  AND3_GATE U57 ( .I1(n143), .I2(n505), .I3(n501), .O(n48) );
  AND3_GATE U58 ( .I1(n50), .I2(n57), .I3(n154), .O(n49) );
  AND3_GATE U59 ( .I1(n46), .I2(n30), .I3(n153), .O(n50) );
  AND_GATE U60 ( .I1(op1[4]), .I2(n1507), .O(n51) );
  AND_GATE U61 ( .I1(n114), .I2(n1507), .O(n52) );
  AND_GATE U62 ( .I1(n399), .I2(op2[0]), .O(n53) );
  AND3_GATE U63 ( .I1(n190), .I2(n189), .I3(n188), .O(n54) );
  AND3_GATE U64 ( .I1(n144), .I2(n39), .I3(n501), .O(n55) );
  NOR_GATE U65 ( .I1(ctrl[14]), .I2(ctrl[13]), .O(n56) );
  NOR_GATE U66 ( .I1(ctrl[2]), .I2(ctrl[11]), .O(n57) );
  NOR4_GATE U67 ( .I1(ctrl[21]), .I2(ctrl[20]), .I3(ctrl[17]), .I4(ctrl[16]), 
        .O(n58) );
  NOR_GATE U68 ( .I1(ctrl[22]), .I2(ctrl[23]), .O(n59) );
  NOR_GATE U69 ( .I1(ctrl[5]), .I2(ctrl[3]), .O(n60) );
  NOR_GATE U70 ( .I1(ctrl[9]), .I2(ctrl[6]), .O(n61) );
  OR3_GATE U71 ( .I1(n62), .I2(n63), .I3(n71), .O(n1944) );
  AND_GATE U72 ( .I1(N820), .I2(n9), .O(n62) );
  AND_GATE U73 ( .I1(N755), .I2(n10), .O(n63) );
  OR3_GATE U74 ( .I1(n64), .I2(n65), .I3(n70), .O(n1928) );
  AND_GATE U75 ( .I1(N836), .I2(n9), .O(n64) );
  AND_GATE U76 ( .I1(N771), .I2(n10), .O(n65) );
  OR3_GATE U77 ( .I1(n66), .I2(n67), .I3(n68), .O(n1929) );
  AND_GATE U78 ( .I1(N770), .I2(n10), .O(n66) );
  AND_GATE U79 ( .I1(N835), .I2(n9), .O(n67) );
  NAND_GATE U80 ( .I1(n2015), .I2(n2014), .O(n68) );
  NAND_GATE U81 ( .I1(n2019), .I2(n2018), .O(n69) );
  NAND_GATE U82 ( .I1(n2017), .I2(n2016), .O(n70) );
  NAND_GATE U83 ( .I1(n1891), .I2(n1892), .O(n71) );
  NAND_GATE U84 ( .I1(n2001), .I2(n2000), .O(n72) );
  NAND_GATE U85 ( .I1(n1878), .I2(n1877), .O(n73) );
  INV_GATE U86 ( .I1(n1452), .O(n74) );
  INV_GATE U87 ( .I1(n1499), .O(n75) );
  INV_GATE U88 ( .I1(n697), .O(n76) );
  INV_GATE U89 ( .I1(n54), .O(n77) );
  INV_GATE U90 ( .I1(op2[0]), .O(n78) );
  INV_GATE U91 ( .I1(op2[1]), .O(n79) );
  INV_GATE U92 ( .I1(op2[2]), .O(n80) );
  INV_GATE U93 ( .I1(op2[3]), .O(n81) );
  INV_GATE U94 ( .I1(op2[4]), .O(n82) );
  INV_GATE U95 ( .I1(op2[5]), .O(n83) );
  INV_GATE U96 ( .I1(op2[6]), .O(n84) );
  INV_GATE U97 ( .I1(op2[7]), .O(n85) );
  INV_GATE U98 ( .I1(op2[8]), .O(n86) );
  INV_GATE U99 ( .I1(op2[9]), .O(n87) );
  INV_GATE U100 ( .I1(op2[10]), .O(n88) );
  INV_GATE U101 ( .I1(op2[11]), .O(n89) );
  INV_GATE U102 ( .I1(op2[12]), .O(n90) );
  INV_GATE U103 ( .I1(op2[13]), .O(n91) );
  INV_GATE U104 ( .I1(op2[14]), .O(n92) );
  INV_GATE U105 ( .I1(op2[15]), .O(n93) );
  INV_GATE U106 ( .I1(op2[16]), .O(n94) );
  INV_GATE U107 ( .I1(op2[17]), .O(n95) );
  INV_GATE U108 ( .I1(op2[18]), .O(n96) );
  INV_GATE U109 ( .I1(op2[19]), .O(n97) );
  INV_GATE U110 ( .I1(op2[20]), .O(n98) );
  INV_GATE U111 ( .I1(op2[21]), .O(n99) );
  INV_GATE U112 ( .I1(op2[22]), .O(n100) );
  INV_GATE U113 ( .I1(op2[23]), .O(n101) );
  INV_GATE U114 ( .I1(op2[24]), .O(n102) );
  INV_GATE U115 ( .I1(op2[25]), .O(n103) );
  INV_GATE U116 ( .I1(op2[26]), .O(n104) );
  INV_GATE U117 ( .I1(op2[27]), .O(n105) );
  INV_GATE U118 ( .I1(op2[28]), .O(n106) );
  INV_GATE U119 ( .I1(op2[29]), .O(n107) );
  INV_GATE U120 ( .I1(op2[30]), .O(n108) );
  INV_GATE U121 ( .I1(op2[31]), .O(n109) );
  INV_GATE U122 ( .I1(op1[0]), .O(n110) );
  INV_GATE U123 ( .I1(op1[1]), .O(n111) );
  INV_GATE U124 ( .I1(op1[2]), .O(n112) );
  INV_GATE U125 ( .I1(op1[3]), .O(n113) );
  INV_GATE U126 ( .I1(op1[4]), .O(n114) );
  INV_GATE U127 ( .I1(op1[5]), .O(n115) );
  INV_GATE U128 ( .I1(op1[6]), .O(n116) );
  INV_GATE U129 ( .I1(op1[7]), .O(n117) );
  INV_GATE U130 ( .I1(op1[8]), .O(n118) );
  INV_GATE U131 ( .I1(op1[9]), .O(n119) );
  INV_GATE U132 ( .I1(op1[10]), .O(n120) );
  INV_GATE U133 ( .I1(op1[11]), .O(n121) );
  INV_GATE U134 ( .I1(op1[12]), .O(n122) );
  INV_GATE U135 ( .I1(op1[13]), .O(n123) );
  INV_GATE U136 ( .I1(op1[14]), .O(n124) );
  INV_GATE U137 ( .I1(op1[15]), .O(n125) );
  INV_GATE U138 ( .I1(op1[16]), .O(n126) );
  INV_GATE U139 ( .I1(op1[17]), .O(n127) );
  INV_GATE U140 ( .I1(op1[18]), .O(n128) );
  INV_GATE U141 ( .I1(op1[19]), .O(n129) );
  INV_GATE U150 ( .I1(op1[20]), .O(n130) );
  INV_GATE U151 ( .I1(op1[21]), .O(n131) );
  INV_GATE U152 ( .I1(op1[22]), .O(n132) );
  INV_GATE U153 ( .I1(op1[23]), .O(n133) );
  INV_GATE U154 ( .I1(op1[24]), .O(n134) );
  INV_GATE U155 ( .I1(op1[25]), .O(n135) );
  INV_GATE U156 ( .I1(op1[26]), .O(n136) );
  INV_GATE U157 ( .I1(op1[27]), .O(n137) );
  INV_GATE U158 ( .I1(op1[28]), .O(n138) );
  INV_GATE U159 ( .I1(op1[29]), .O(n139) );
  INV_GATE U160 ( .I1(op1[30]), .O(n140) );
  INV_GATE U161 ( .I1(op1[31]), .O(n141) );
  NAND_GATE U162 ( .I1(ctrl[15]), .I2(n58), .O(n142) );
  INV_GATE U163 ( .I1(ctrl[8]), .O(n143) );
  OR3_GATE U164 ( .I1(ctrl[19]), .I2(ctrl[18]), .I3(ctrl[1]), .O(n147) );
  INV_GATE U165 ( .I1(ctrl[24]), .O(n145) );
  OR_GATE U166 ( .I1(ctrl[27]), .I2(ctrl[25]), .O(n531) );
  INV_GATE U167 ( .I1(n531), .O(n187) );
  NAND_GATE U168 ( .I1(n145), .I2(n187), .O(n371) );
  NOR4_GATE U169 ( .I1(n147), .I2(n371), .I3(ctrl[4]), .I4(ctrl[26]), .O(n505)
         );
  INV_GATE U178 ( .I1(ctrl[7]), .O(n501) );
  INV_GATE U179 ( .I1(ctrl[0]), .O(n153) );
  INV_GATE U180 ( .I1(ctrl[12]), .O(n455) );
  INV_GATE U181 ( .I1(ctrl[10]), .O(n154) );
  NAND3_GATE U182 ( .I1(n30), .I2(n41), .I3(n59), .O(n488) );
  OR_GATE U183 ( .I1(n142), .I2(n488), .O(n474) );
  INV_GATE U184 ( .I1(ctrl[26]), .O(n527) );
  INV_GATE U185 ( .I1(ctrl[4]), .O(n144) );
  INV_GATE U186 ( .I1(ctrl[15]), .O(n486) );
  NOR_GATE U187 ( .I1(ctrl[18]), .I2(ctrl[1]), .O(n146) );
  NAND3_GATE U189 ( .I1(ctrl[19]), .I2(n187), .I3(n146), .O(n151) );
  INV_GATE U190 ( .I1(n147), .O(n532) );
  INV_GATE U191 ( .I1(ctrl[27]), .O(n148) );
  NAND_GATE U192 ( .I1(ctrl[25]), .I2(n148), .O(n183) );
  INV_GATE U193 ( .I1(ctrl[25]), .O(n354) );
  NAND_GATE U194 ( .I1(n354), .I2(ctrl[27]), .O(n149) );
  NAND_GATE U195 ( .I1(n183), .I2(n149), .O(n524) );
  NAND_GATE U196 ( .I1(n532), .I2(n524), .O(n150) );
  NAND_GATE U197 ( .I1(n151), .I2(n150), .O(n152) );
  NAND_GATE U206 ( .I1(n42), .I2(n152), .O(n173) );
  INV_GATE U207 ( .I1(ctrl[14]), .O(n470) );
  NAND_GATE U208 ( .I1(ctrl[13]), .I2(n470), .O(n156) );
  INV_GATE U209 ( .I1(ctrl[13]), .O(n440) );
  NAND_GATE U210 ( .I1(n440), .I2(ctrl[14]), .O(n155) );
  NAND_GATE U212 ( .I1(n156), .I2(n155), .O(n157) );
  NAND3_GATE U213 ( .I1(n49), .I2(n157), .I3(n455), .O(n192) );
  NAND3_GATE U214 ( .I1(ctrl[12]), .I2(n49), .I3(n56), .O(n158) );
  AND_GATE U217 ( .I1(n192), .I2(n158), .O(n168) );
  NAND3_GATE U218 ( .I1(n474), .I2(n173), .I3(n168), .O(n191) );
  AND_GATE U219 ( .I1(op1[31]), .I2(n191), .O(\efct_op1[32] ) );
  NOR4_GATE U220 ( .I1(ctrl[21]), .I2(n488), .I3(ctrl[20]), .I4(ctrl[15]), .O(
        n180) );
  INV_GATE U221 ( .I1(ctrl[16]), .O(n176) );
  NAND3_GATE U222 ( .I1(ctrl[17]), .I2(n180), .I3(n176), .O(n545) );
  INV_GATE U223 ( .I1(ctrl[17]), .O(n179) );
  NAND3_GATE U224 ( .I1(ctrl[16]), .I2(n180), .I3(n179), .O(n558) );
  AND_GATE U225 ( .I1(n545), .I2(n558), .O(n190) );
  INV_GATE U234 ( .I1(ctrl[19]), .O(n394) );
  NAND_GATE U235 ( .I1(ctrl[18]), .I2(n394), .O(n182) );
  INV_GATE U236 ( .I1(ctrl[18]), .O(n393) );
  NAND_GATE U237 ( .I1(n393), .I2(ctrl[19]), .O(n181) );
  NAND_GATE U238 ( .I1(n182), .I2(n181), .O(n380) );
  INV_GATE U240 ( .I1(ctrl[1]), .O(n392) );
  NAND3_GATE U241 ( .I1(n380), .I2(n392), .I3(n187), .O(n185) );
  INV_GATE U242 ( .I1(n183), .O(n355) );
  NAND_GATE U245 ( .I1(n532), .I2(n355), .O(n184) );
  NAND_GATE U246 ( .I1(n185), .I2(n184), .O(n186) );
  NAND_GATE U247 ( .I1(n42), .I2(n186), .O(n189) );
  NAND4_GATE U248 ( .I1(ctrl[24]), .I2(n532), .I3(n40), .I4(n187), .O(n188) );
  NAND_GATE U249 ( .I1(op2[31]), .I2(n191), .O(n193) );
  NAND_GATE U250 ( .I1(n77), .I2(n193), .O(n195) );
  NAND_GATE U251 ( .I1(n54), .I2(n192), .O(n196) );
  OR_GATE U252 ( .I1(n196), .I2(n193), .O(n194) );
  NAND_GATE U253 ( .I1(n195), .I2(n194), .O(efct_op2[32]) );
  NAND_GATE U262 ( .I1(n109), .I2(n77), .O(n198) );
  INV_GATE U263 ( .I1(n196), .O(n342) );
  NAND_GATE U264 ( .I1(op2[31]), .I2(n342), .O(n197) );
  NAND_GATE U265 ( .I1(n198), .I2(n197), .O(efct_op2[31]) );
  NAND_GATE U266 ( .I1(op2[30]), .I2(n342), .O(n200) );
  NAND_GATE U268 ( .I1(n108), .I2(n77), .O(n199) );
  NAND_GATE U269 ( .I1(n200), .I2(n199), .O(efct_op2[30]) );
  NAND_GATE U270 ( .I1(op2[29]), .I2(n342), .O(n202) );
  NAND_GATE U273 ( .I1(n107), .I2(n77), .O(n201) );
  NAND_GATE U274 ( .I1(n202), .I2(n201), .O(efct_op2[29]) );
  NAND_GATE U275 ( .I1(op2[28]), .I2(n342), .O(n204) );
  NAND_GATE U276 ( .I1(n106), .I2(n77), .O(n203) );
  NAND_GATE U277 ( .I1(n204), .I2(n203), .O(efct_op2[28]) );
  NAND_GATE U278 ( .I1(op2[27]), .I2(n342), .O(n217) );
  NAND_GATE U279 ( .I1(n105), .I2(n77), .O(n213) );
  NAND_GATE U288 ( .I1(n217), .I2(n213), .O(efct_op2[27]) );
  NAND_GATE U289 ( .I1(op2[26]), .I2(n342), .O(n219) );
  NAND_GATE U290 ( .I1(n104), .I2(n77), .O(n218) );
  NAND_GATE U291 ( .I1(n219), .I2(n218), .O(efct_op2[26]) );
  NAND_GATE U292 ( .I1(op2[25]), .I2(n342), .O(n221) );
  NAND_GATE U294 ( .I1(n103), .I2(n77), .O(n220) );
  NAND_GATE U295 ( .I1(n221), .I2(n220), .O(efct_op2[25]) );
  NAND_GATE U297 ( .I1(op2[24]), .I2(n342), .O(n228) );
  NAND_GATE U298 ( .I1(n102), .I2(n77), .O(n227) );
  NAND_GATE U299 ( .I1(n228), .I2(n227), .O(efct_op2[24]) );
  NAND_GATE U301 ( .I1(op2[23]), .I2(n342), .O(n230) );
  NAND_GATE U302 ( .I1(n101), .I2(n77), .O(n229) );
  NAND_GATE U303 ( .I1(n230), .I2(n229), .O(efct_op2[23]) );
  NAND_GATE U304 ( .I1(op2[22]), .I2(n342), .O(n232) );
  NAND_GATE U305 ( .I1(n100), .I2(n77), .O(n231) );
  NAND_GATE U306 ( .I1(n232), .I2(n231), .O(efct_op2[22]) );
  NAND_GATE U307 ( .I1(op2[21]), .I2(n342), .O(n234) );
  NAND_GATE U308 ( .I1(n99), .I2(n77), .O(n233) );
  NAND_GATE U310 ( .I1(n234), .I2(n233), .O(efct_op2[21]) );
  NAND_GATE U311 ( .I1(op2[20]), .I2(n342), .O(n236) );
  NAND_GATE U312 ( .I1(n98), .I2(n77), .O(n235) );
  NAND_GATE U313 ( .I1(n236), .I2(n235), .O(efct_op2[20]) );
  NAND_GATE U314 ( .I1(op2[19]), .I2(n342), .O(n250) );
  NAND_GATE U315 ( .I1(n97), .I2(n77), .O(n249) );
  NAND_GATE U316 ( .I1(n250), .I2(n249), .O(efct_op2[19]) );
  NAND_GATE U317 ( .I1(op2[18]), .I2(n342), .O(n259) );
  NAND_GATE U318 ( .I1(n96), .I2(n77), .O(n252) );
  NAND_GATE U330 ( .I1(n259), .I2(n252), .O(efct_op2[18]) );
  NAND_GATE U331 ( .I1(op2[17]), .I2(n342), .O(n261) );
  NAND_GATE U332 ( .I1(n95), .I2(n77), .O(n260) );
  NAND_GATE U333 ( .I1(n261), .I2(n260), .O(efct_op2[17]) );
  NAND_GATE U334 ( .I1(op2[16]), .I2(n342), .O(n263) );
  NAND_GATE U338 ( .I1(n94), .I2(n77), .O(n262) );
  NAND_GATE U339 ( .I1(n263), .I2(n262), .O(efct_op2[16]) );
  NAND_GATE U340 ( .I1(op2[15]), .I2(n342), .O(n265) );
  NAND_GATE U342 ( .I1(n93), .I2(n77), .O(n264) );
  NAND_GATE U343 ( .I1(n265), .I2(n264), .O(efct_op2[15]) );
  NAND_GATE U344 ( .I1(op2[14]), .I2(n342), .O(n267) );
  NAND_GATE U345 ( .I1(n92), .I2(n77), .O(n266) );
  NAND_GATE U346 ( .I1(n267), .I2(n266), .O(efct_op2[14]) );
  NAND_GATE U347 ( .I1(op2[13]), .I2(n342), .O(n277) );
  NAND_GATE U348 ( .I1(n91), .I2(n77), .O(n268) );
  NAND_GATE U349 ( .I1(n277), .I2(n268), .O(efct_op2[13]) );
  NAND_GATE U360 ( .I1(op2[12]), .I2(n342), .O(n283) );
  NAND_GATE U361 ( .I1(n90), .I2(n77), .O(n282) );
  NAND_GATE U362 ( .I1(n283), .I2(n282), .O(efct_op2[12]) );
  NAND_GATE U363 ( .I1(op2[11]), .I2(n342), .O(n292) );
  NAND_GATE U364 ( .I1(n89), .I2(n77), .O(n285) );
  NAND_GATE U365 ( .I1(n292), .I2(n285), .O(efct_op2[11]) );
  NAND_GATE U366 ( .I1(op2[10]), .I2(n342), .O(n294) );
  NAND_GATE U367 ( .I1(n88), .I2(n77), .O(n293) );
  NAND_GATE U368 ( .I1(n294), .I2(n293), .O(efct_op2[10]) );
  NAND_GATE U369 ( .I1(op2[9]), .I2(n342), .O(n296) );
  NAND_GATE U370 ( .I1(n87), .I2(n77), .O(n295) );
  NAND_GATE U371 ( .I1(n296), .I2(n295), .O(efct_op2[9]) );
  NAND_GATE U372 ( .I1(op2[8]), .I2(n342), .O(n298) );
  NAND_GATE U373 ( .I1(n86), .I2(n77), .O(n297) );
  NAND_GATE U374 ( .I1(n298), .I2(n297), .O(efct_op2[8]) );
  NAND_GATE U375 ( .I1(op2[7]), .I2(n342), .O(n300) );
  NAND_GATE U376 ( .I1(n85), .I2(n77), .O(n299) );
  NAND_GATE U377 ( .I1(n300), .I2(n299), .O(efct_op2[7]) );
  NAND_GATE U378 ( .I1(op2[6]), .I2(n342), .O(n312) );
  NAND_GATE U379 ( .I1(n84), .I2(n77), .O(n301) );
  NAND_GATE U380 ( .I1(n312), .I2(n301), .O(efct_op2[6]) );
  NAND_GATE U381 ( .I1(op2[5]), .I2(n342), .O(n315) );
  NAND_GATE U382 ( .I1(n83), .I2(n77), .O(n313) );
  NAND_GATE U383 ( .I1(n315), .I2(n313), .O(efct_op2[5]) );
  NAND_GATE U392 ( .I1(op2[4]), .I2(n342), .O(n323) );
  NAND_GATE U393 ( .I1(n82), .I2(n77), .O(n322) );
  NAND_GATE U394 ( .I1(n323), .I2(n322), .O(efct_op2[4]) );
  NAND_GATE U395 ( .I1(op2[3]), .I2(n342), .O(n325) );
  NAND_GATE U396 ( .I1(n81), .I2(n77), .O(n324) );
  NAND_GATE U397 ( .I1(n325), .I2(n324), .O(efct_op2[3]) );
  NAND_GATE U398 ( .I1(op2[2]), .I2(n342), .O(n328) );
  NAND_GATE U399 ( .I1(n80), .I2(n77), .O(n326) );
  NAND_GATE U400 ( .I1(n328), .I2(n326), .O(efct_op2[2]) );
  NAND_GATE U401 ( .I1(op2[1]), .I2(n342), .O(n330) );
  NAND_GATE U402 ( .I1(n79), .I2(n77), .O(n329) );
  NAND_GATE U403 ( .I1(n330), .I2(n329), .O(efct_op2[1]) );
  NAND_GATE U404 ( .I1(op2[0]), .I2(n342), .O(n345) );
  NAND_GATE U406 ( .I1(n78), .I2(n77), .O(n343) );
  NAND_GATE U407 ( .I1(n345), .I2(n343), .O(efct_op2[0]) );
  OR_GATE U408 ( .I1(n141), .I2(res_add[31]), .O(n353) );
  NAND_GATE U409 ( .I1(res_add[31]), .I2(n141), .O(n347) );
  NAND_GATE U410 ( .I1(n353), .I2(n347), .O(n360) );
  NAND3_GATE U411 ( .I1(n1909), .I2(ctrl[27]), .I3(n354), .O(n357) );
  NAND_GATE U412 ( .I1(n417), .I2(n355), .O(n356) );
  NAND_GATE U413 ( .I1(n357), .I2(n356), .O(n359) );
  AND_GATE U415 ( .I1(n532), .I2(n42), .O(n358) );
  AND3_GATE U416 ( .I1(n360), .I2(n359), .I3(n358), .O(N1035) );
  NAND_GATE U417 ( .I1(n399), .I2(n90), .O(n369) );
  NAND_GATE U418 ( .I1(n398), .I2(n91), .O(n368) );
  NAND_GATE U419 ( .I1(n397), .I2(n92), .O(n367) );
  NAND_GATE U420 ( .I1(n396), .I2(n93), .O(n366) );
  NAND4_GATE U421 ( .I1(n369), .I2(n368), .I3(n367), .I4(n366), .O(n339) );
  NOR_GATE U422 ( .I1(ctrl[2]), .I2(ctrl[10]), .O(n370) );
  NAND3_GATE U423 ( .I1(ctrl[11]), .I2(n32), .I3(n370), .O(n1523) );
  NAND3_GATE U435 ( .I1(ctrl[10]), .I2(n57), .I3(n32), .O(n1525) );
  AND_GATE U436 ( .I1(ctrl[4]), .I2(n532), .O(n373) );
  INV_GATE U437 ( .I1(n371), .O(n528) );
  AND3_GATE U438 ( .I1(n501), .I2(n528), .I3(n527), .O(n372) );
  NAND3_GATE U439 ( .I1(n39), .I2(n373), .I3(n372), .O(n378) );
  NAND3_GATE U443 ( .I1(n1523), .I2(n1525), .I3(n378), .O(n178) );
  AND_GATE U444 ( .I1(n528), .I2(n40), .O(n404) );
  NAND3_GATE U445 ( .I1(n392), .I2(n380), .I3(res_add[32]), .O(n402) );
  NAND3_GATE U447 ( .I1(n394), .I2(n393), .I3(ctrl[1]), .O(n395) );
  NAND_GATE U448 ( .I1(n376), .I2(n81), .O(n406) );
  NAND_GATE U449 ( .I1(n377), .I2(n80), .O(n405) );
  AND_GATE U450 ( .I1(n406), .I2(n405), .O(n438) );
  NAND_GATE U451 ( .I1(n375), .I2(n79), .O(n408) );
  NAND_GATE U452 ( .I1(n374), .I2(n78), .O(n407) );
  AND_GATE U453 ( .I1(n408), .I2(n407), .O(n437) );
  INV_GATE U454 ( .I1(n171), .O(n2047) );
  NAND_GATE U455 ( .I1(n2047), .I2(n339), .O(n414) );
  NAND_GATE U456 ( .I1(n399), .I2(n82), .O(n412) );
  NAND_GATE U457 ( .I1(n398), .I2(n83), .O(n411) );
  NAND_GATE U458 ( .I1(n397), .I2(n84), .O(n410) );
  NAND_GATE U459 ( .I1(n396), .I2(n85), .O(n409) );
  NAND4_GATE U460 ( .I1(n412), .I2(n411), .I3(n410), .I4(n409), .O(n1533) );
  NAND_GATE U461 ( .I1(n167), .I2(n1533), .O(n413) );
  AND_GATE U462 ( .I1(n414), .I2(n413), .O(n436) );
  INV_GATE U463 ( .I1(n169), .O(n2046) );
  NAND_GATE U464 ( .I1(n399), .I2(n86), .O(n433) );
  NAND_GATE U473 ( .I1(n398), .I2(n87), .O(n418) );
  NAND_GATE U474 ( .I1(n397), .I2(n88), .O(n416) );
  NAND_GATE U475 ( .I1(n396), .I2(n89), .O(n415) );
  NAND4_GATE U476 ( .I1(n433), .I2(n418), .I3(n416), .I4(n415), .O(n1534) );
  NAND_GATE U477 ( .I1(n2046), .I2(n1534), .O(n435) );
  NAND4_GATE U478 ( .I1(op2[31]), .I2(ctrl[7]), .I3(n39), .I4(n505), .O(n1512)
         );
  INV_GATE U479 ( .I1(n1512), .O(n1635) );
  AND_GATE U480 ( .I1(n1446), .I2(n1635), .O(n434) );
  NAND5_GATE U481 ( .I1(n438), .I2(n437), .I3(n436), .I4(n435), .I5(n434), .O(
        n439) );
  NAND3_GATE U482 ( .I1(n440), .I2(n141), .I3(ctrl[12]), .O(n457) );
  NOR_GATE U483 ( .I1(res_add[14]), .I2(res_add[15]), .O(n454) );
  NOR4_GATE U484 ( .I1(res_add[2]), .I2(res_add[3]), .I3(res_add[1]), .I4(
        res_add[0]), .O(n445) );
  NOR_GATE U485 ( .I1(res_add[5]), .I2(res_add[4]), .O(n444) );
  NOR_GATE U486 ( .I1(res_add[6]), .I2(res_add[7]), .O(n443) );
  NOR4_GATE U487 ( .I1(res_add[10]), .I2(res_add[11]), .I3(res_add[9]), .I4(
        res_add[8]), .O(n442) );
  NOR_GATE U488 ( .I1(res_add[13]), .I2(res_add[12]), .O(n441) );
  AND5_GATE U489 ( .I1(n445), .I2(n444), .I3(n443), .I4(n442), .I5(n441), .O(
        n453) );
  NOR_GATE U490 ( .I1(res_add[31]), .I2(res_add[30]), .O(n452) );
  NOR4_GATE U499 ( .I1(res_add[18]), .I2(res_add[19]), .I3(res_add[17]), .I4(
        res_add[16]), .O(n450) );
  NOR_GATE U500 ( .I1(res_add[21]), .I2(res_add[20]), .O(n449) );
  NOR_GATE U501 ( .I1(res_add[22]), .I2(res_add[23]), .O(n448) );
  NOR4_GATE U502 ( .I1(res_add[26]), .I2(res_add[27]), .I3(res_add[25]), .I4(
        res_add[24]), .O(n447) );
  NOR_GATE U503 ( .I1(res_add[29]), .I2(res_add[28]), .O(n446) );
  AND5_GATE U504 ( .I1(n450), .I2(n449), .I3(n448), .I4(n447), .I5(n446), .O(
        n451) );
  NAND4_GATE U505 ( .I1(n454), .I2(n453), .I3(n452), .I4(n451), .O(n546) );
  NAND_GATE U506 ( .I1(n141), .I2(n546), .O(n471) );
  NAND3_GATE U507 ( .I1(n455), .I2(ctrl[13]), .I3(n471), .O(n456) );
  NAND_GATE U508 ( .I1(n457), .I2(n456), .O(n458) );
  NOR3_GATE U509 ( .I1(n471), .I2(ctrl[13]), .I3(ctrl[12]), .O(n472) );
  NAND_GATE U510 ( .I1(n472), .I2(ctrl[14]), .O(n473) );
  INV_GATE U511 ( .I1(n474), .O(n475) );
  NAND_GATE U512 ( .I1(op1[31]), .I2(n475), .O(n519) );
  INV_GATE U513 ( .I1(ctrl[5]), .O(n477) );
  AND_GATE U514 ( .I1(ctrl[3]), .I2(n61), .O(n476) );
  NAND3_GATE U515 ( .I1(n477), .I2(n31), .I3(n476), .O(n1524) );
  NOR_GATE U516 ( .I1(ctrl[11]), .I2(ctrl[10]), .O(n478) );
  NAND3_GATE U517 ( .I1(ctrl[2]), .I2(n32), .I3(n478), .O(n480) );
  NAND_GATE U518 ( .I1(n1524), .I2(n480), .O(n1689) );
  INV_GATE U524 ( .I1(n1689), .O(n1619) );
  AND4_GATE U525 ( .I1(n58), .I2(n41), .I3(n30), .I4(n486), .O(n491) );
  INV_GATE U526 ( .I1(ctrl[23]), .O(n487) );
  NAND3_GATE U527 ( .I1(ctrl[22]), .I2(n491), .I3(n487), .O(n1688) );
  NAND_GATE U528 ( .I1(n1619), .I2(n1688), .O(n1509) );
  INV_GATE U529 ( .I1(n1509), .O(n1456) );
  NOR4_GATE U530 ( .I1(ctrl[17]), .I2(n488), .I3(ctrl[16]), .I4(ctrl[15]), .O(
        n539) );
  INV_GATE U531 ( .I1(ctrl[20]), .O(n489) );
  NAND3_GATE U532 ( .I1(ctrl[21]), .I2(n539), .I3(n489), .O(n1452) );
  NAND_GATE U533 ( .I1(n78), .I2(n1452), .O(n498) );
  INV_GATE U534 ( .I1(ctrl[22]), .O(n490) );
  NAND3_GATE U535 ( .I1(ctrl[23]), .I2(n491), .I3(n490), .O(n1499) );
  NAND_GATE U536 ( .I1(op2[0]), .I2(n1499), .O(n492) );
  NAND_GATE U537 ( .I1(n498), .I2(n492), .O(n499) );
  NAND_GATE U538 ( .I1(n1456), .I2(n499), .O(n500) );
  NAND_GATE U539 ( .I1(op1[0]), .I2(n500), .O(n518) );
  NAND3_GATE U540 ( .I1(n501), .I2(ctrl[8]), .I3(n28), .O(n503) );
  NAND_GATE U541 ( .I1(ctrl[7]), .I2(n39), .O(n502) );
  NAND_GATE U542 ( .I1(n503), .I2(n502), .O(n504) );
  AND_GATE U543 ( .I1(n505), .I2(n504), .O(n1701) );
  NAND_GATE U544 ( .I1(n1464), .I2(n6), .O(n506) );
  AND3_GATE U545 ( .I1(n519), .I2(n518), .I3(n506), .O(n568) );
  NAND3_GATE U546 ( .I1(ctrl[5]), .I2(n61), .I3(n31), .O(n520) );
  NOR_GATE U547 ( .I1(ctrl[3]), .I2(n520), .O(n1700) );
  NAND_GATE U548 ( .I1(hilo[32]), .I2(n1700), .O(n537) );
  NAND3_GATE U549 ( .I1(ctrl[9]), .I2(n60), .I3(n31), .O(n521) );
  NOR_GATE U550 ( .I1(ctrl[6]), .I2(n521), .O(n1507) );
  NAND_GATE U556 ( .I1(n13), .I2(n53), .O(n536) );
  OR_GATE U557 ( .I1(n524), .I2(ctrl[24]), .O(n526) );
  NAND_GATE U558 ( .I1(n527), .I2(n526), .O(n530) );
  NAND_GATE U559 ( .I1(ctrl[26]), .I2(n528), .O(n529) );
  NAND_GATE U560 ( .I1(n530), .I2(n529), .O(n534) );
  NAND_GATE U561 ( .I1(ctrl[24]), .I2(n531), .O(n533) );
  AND4_GATE U562 ( .I1(n534), .I2(n533), .I3(n55), .I4(n532), .O(n1691) );
  NAND_GATE U563 ( .I1(res_add[0]), .I2(n1691), .O(n535) );
  AND3_GATE U564 ( .I1(n537), .I2(n536), .I3(n535), .O(n566) );
  INV_GATE U565 ( .I1(ctrl[21]), .O(n538) );
  NAND3_GATE U566 ( .I1(ctrl[20]), .I2(n539), .I3(n538), .O(n1637) );
  INV_GATE U567 ( .I1(n1637), .O(n1694) );
  NAND_GATE U568 ( .I1(n110), .I2(n1694), .O(n540) );
  NAND_GATE U569 ( .I1(n78), .I2(n540), .O(n544) );
  NAND4_GATE U570 ( .I1(ctrl[0]), .I2(n46), .I3(n43), .I4(n30), .O(n1696) );
  AND_GATE U571 ( .I1(op2[0]), .I2(n12), .O(n542) );
  NAND_GATE U572 ( .I1(n110), .I2(n74), .O(n541) );
  NAND_GATE U573 ( .I1(n542), .I2(n541), .O(n543) );
  NAND_GATE U574 ( .I1(n544), .I2(n543), .O(n565) );
  NAND_GATE U575 ( .I1(n558), .I2(n546), .O(n559) );
  NAND_GATE U576 ( .I1(n560), .I2(n559), .O(n564) );
  NAND_GATE U577 ( .I1(hilo[0]), .I2(n178), .O(n561) );
  AND4_GATE U578 ( .I1(n566), .I2(n565), .I3(n564), .I4(n561), .O(n567) );
  NAND4_GATE U579 ( .I1(n570), .I2(n569), .I3(n568), .I4(n567), .O(res[0]) );
  NAND_GATE U580 ( .I1(res_add[8]), .I2(n1691), .O(n600) );
  NAND_GATE U581 ( .I1(hilo[8]), .I2(n178), .O(n599) );
  NAND_GATE U582 ( .I1(n118), .I2(n1694), .O(n571) );
  NAND_GATE U588 ( .I1(n86), .I2(n571), .O(n575) );
  AND_GATE U589 ( .I1(op2[8]), .I2(n12), .O(n573) );
  NAND_GATE U590 ( .I1(n118), .I2(n74), .O(n572) );
  NAND_GATE U594 ( .I1(n573), .I2(n572), .O(n574) );
  NAND_GATE U595 ( .I1(n575), .I2(n574), .O(n598) );
  NAND_GATE U596 ( .I1(n205), .I2(n1701), .O(n596) );
  NAND_GATE U597 ( .I1(hilo[40]), .I2(n1700), .O(n595) );
  NAND_GATE U598 ( .I1(n86), .I2(n1452), .O(n577) );
  NAND_GATE U599 ( .I1(op2[8]), .I2(n1499), .O(n576) );
  NAND_GATE U600 ( .I1(n577), .I2(n576), .O(n578) );
  NAND_GATE U601 ( .I1(n1456), .I2(n578), .O(n579) );
  NAND_GATE U602 ( .I1(op1[8]), .I2(n579), .O(n593) );
  NAND_GATE U603 ( .I1(n695), .I2(n53), .O(n591) );
  NAND3_GATE U604 ( .I1(n737), .I2(n735), .I3(n591), .O(n1128) );
  NAND_GATE U605 ( .I1(n52), .I2(n1128), .O(n592) );
  AND_GATE U606 ( .I1(n593), .I2(n592), .O(n594) );
  AND3_GATE U607 ( .I1(n596), .I2(n595), .I3(n594), .O(n597) );
  NAND4_GATE U608 ( .I1(n600), .I2(n599), .I3(n598), .I4(n597), .O(res[8]) );
  NAND_GATE U612 ( .I1(res_add[9]), .I2(n1691), .O(n623) );
  NAND_GATE U613 ( .I1(hilo[9]), .I2(n178), .O(n622) );
  NAND_GATE U614 ( .I1(n119), .I2(n1694), .O(n601) );
  NAND_GATE U618 ( .I1(n87), .I2(n601), .O(n605) );
  AND_GATE U619 ( .I1(op2[9]), .I2(n12), .O(n603) );
  NAND_GATE U620 ( .I1(n119), .I2(n74), .O(n602) );
  NAND_GATE U621 ( .I1(n603), .I2(n602), .O(n604) );
  NAND_GATE U622 ( .I1(n605), .I2(n604), .O(n621) );
  NAND_GATE U623 ( .I1(n159), .I2(n1701), .O(n618) );
  NAND_GATE U624 ( .I1(hilo[41]), .I2(n1700), .O(n617) );
  NAND3_GATE U630 ( .I1(n692), .I2(n691), .I3(n690), .O(n1182) );
  NAND_GATE U631 ( .I1(n52), .I2(n1182), .O(n611) );
  NAND_GATE U632 ( .I1(n87), .I2(n1452), .O(n607) );
  NAND_GATE U634 ( .I1(op2[9]), .I2(n1499), .O(n606) );
  NAND_GATE U636 ( .I1(n607), .I2(n606), .O(n608) );
  NAND_GATE U637 ( .I1(n1456), .I2(n608), .O(n609) );
  NAND_GATE U638 ( .I1(op1[9]), .I2(n609), .O(n610) );
  AND_GATE U639 ( .I1(n611), .I2(n610), .O(n616) );
  AND3_GATE U640 ( .I1(n618), .I2(n617), .I3(n616), .O(n620) );
  NAND4_GATE U641 ( .I1(n623), .I2(n622), .I3(n621), .I4(n620), .O(res[9]) );
  NAND_GATE U642 ( .I1(res_add[10]), .I2(n1691), .O(n643) );
  NAND_GATE U643 ( .I1(hilo[10]), .I2(n178), .O(n642) );
  NAND_GATE U644 ( .I1(n120), .I2(n1694), .O(n624) );
  NAND_GATE U645 ( .I1(n88), .I2(n624), .O(n628) );
  AND_GATE U646 ( .I1(op2[10]), .I2(n12), .O(n626) );
  NAND_GATE U647 ( .I1(n120), .I2(n74), .O(n625) );
  NAND_GATE U648 ( .I1(n626), .I2(n625), .O(n627) );
  NAND_GATE U649 ( .I1(n628), .I2(n627), .O(n641) );
  NAND_GATE U650 ( .I1(n1383), .I2(n1701), .O(n639) );
  NAND_GATE U654 ( .I1(hilo[42]), .I2(n1700), .O(n638) );
  NAND3_GATE U655 ( .I1(n1424), .I2(n1423), .I3(n1422), .O(n1238) );
  NAND_GATE U656 ( .I1(n52), .I2(n1238), .O(n636) );
  NAND_GATE U660 ( .I1(n88), .I2(n1452), .O(n630) );
  NAND_GATE U661 ( .I1(op2[10]), .I2(n1499), .O(n629) );
  NAND_GATE U662 ( .I1(n630), .I2(n629), .O(n633) );
  NAND_GATE U663 ( .I1(n1456), .I2(n633), .O(n634) );
  NAND_GATE U664 ( .I1(op1[10]), .I2(n634), .O(n635) );
  AND_GATE U665 ( .I1(n636), .I2(n635), .O(n637) );
  AND3_GATE U666 ( .I1(n639), .I2(n638), .I3(n637), .O(n640) );
  NAND4_GATE U672 ( .I1(n643), .I2(n642), .I3(n641), .I4(n640), .O(res[10]) );
  NAND_GATE U673 ( .I1(res_add[11]), .I2(n1691), .O(n666) );
  NAND_GATE U677 ( .I1(hilo[11]), .I2(n178), .O(n665) );
  NAND_GATE U678 ( .I1(n121), .I2(n1694), .O(n644) );
  NAND_GATE U679 ( .I1(n89), .I2(n644), .O(n648) );
  AND_GATE U680 ( .I1(op2[11]), .I2(n12), .O(n646) );
  NAND_GATE U681 ( .I1(n121), .I2(n74), .O(n645) );
  NAND_GATE U682 ( .I1(n646), .I2(n645), .O(n647) );
  NAND_GATE U683 ( .I1(n648), .I2(n647), .O(n664) );
  NAND_GATE U684 ( .I1(n1318), .I2(n1701), .O(n662) );
  NAND_GATE U685 ( .I1(hilo[43]), .I2(n1700), .O(n661) );
  NAND3_GATE U686 ( .I1(n1355), .I2(n1354), .I3(n1353), .O(n1304) );
  NAND_GATE U687 ( .I1(n52), .I2(n1304), .O(n659) );
  NAND_GATE U688 ( .I1(n89), .I2(n1452), .O(n650) );
  NAND_GATE U689 ( .I1(op2[11]), .I2(n1499), .O(n649) );
  NAND_GATE U690 ( .I1(n650), .I2(n649), .O(n651) );
  NAND_GATE U691 ( .I1(n1456), .I2(n651), .O(n656) );
  NAND_GATE U696 ( .I1(op1[11]), .I2(n656), .O(n658) );
  AND_GATE U697 ( .I1(n659), .I2(n658), .O(n660) );
  AND3_GATE U698 ( .I1(n662), .I2(n661), .I3(n660), .O(n663) );
  NAND4_GATE U702 ( .I1(n666), .I2(n665), .I3(n664), .I4(n663), .O(res[11]) );
  NAND_GATE U703 ( .I1(op1[4]), .I2(n1635), .O(n2050) );
  INV_GATE U704 ( .I1(n2050), .O(n2042) );
  NAND_GATE U705 ( .I1(n76), .I2(n2042), .O(n1168) );
  NAND_GATE U706 ( .I1(op1[4]), .I2(n1512), .O(n2051) );
  NAND_GATE U707 ( .I1(hilo[44]), .I2(n1700), .O(n703) );
  NAND_GATE U708 ( .I1(n90), .I2(n1452), .O(n669) );
  NAND_GATE U714 ( .I1(op2[12]), .I2(n1499), .O(n668) );
  NAND_GATE U715 ( .I1(n669), .I2(n668), .O(n670) );
  NAND_GATE U719 ( .I1(n1456), .I2(n670), .O(n671) );
  NAND_GATE U720 ( .I1(op1[12]), .I2(n671), .O(n702) );
  NAND3_GATE U721 ( .I1(n1272), .I2(n1271), .I3(n1270), .O(n1350) );
  NAND_GATE U722 ( .I1(n52), .I2(n1350), .O(n677) );
  INV_GATE U723 ( .I1(n339), .O(n2043) );
  NAND_GATE U724 ( .I1(n175), .I2(n2043), .O(n674) );
  NAND_GATE U725 ( .I1(n1292), .I2(n2051), .O(n673) );
  NAND4_GATE U726 ( .I1(n674), .I2(n673), .I3(n1168), .I4(n1290), .O(n675) );
  NAND_GATE U727 ( .I1(n1701), .I2(n675), .O(n676) );
  AND_GATE U728 ( .I1(n677), .I2(n676), .O(n701) );
  NAND_GATE U729 ( .I1(n122), .I2(n1694), .O(n678) );
  NAND_GATE U730 ( .I1(n90), .I2(n678), .O(n682) );
  AND_GATE U731 ( .I1(op2[12]), .I2(n12), .O(n680) );
  NAND_GATE U732 ( .I1(n122), .I2(n74), .O(n679) );
  NAND_GATE U733 ( .I1(n680), .I2(n679), .O(n681) );
  NAND_GATE U738 ( .I1(n682), .I2(n681), .O(n700) );
  NAND_GATE U739 ( .I1(hilo[12]), .I2(n178), .O(n684) );
  NAND_GATE U740 ( .I1(res_add[12]), .I2(n1691), .O(n683) );
  AND_GATE U745 ( .I1(n684), .I2(n683), .O(n685) );
  NAND5_GATE U746 ( .I1(n703), .I2(n702), .I3(n701), .I4(n700), .I5(n685), .O(
        res[12]) );
  NAND_GATE U747 ( .I1(res_add[13]), .I2(n1691), .O(n726) );
  NAND_GATE U748 ( .I1(hilo[13]), .I2(n178), .O(n725) );
  NAND_GATE U749 ( .I1(n123), .I2(n1694), .O(n704) );
  NAND_GATE U750 ( .I1(n91), .I2(n704), .O(n708) );
  AND_GATE U751 ( .I1(op2[13]), .I2(n12), .O(n706) );
  NAND_GATE U757 ( .I1(n123), .I2(n74), .O(n705) );
  NAND_GATE U758 ( .I1(n706), .I2(n705), .O(n707) );
  NAND_GATE U762 ( .I1(n708), .I2(n707), .O(n724) );
  NAND_GATE U763 ( .I1(n1203), .I2(n1701), .O(n722) );
  NAND_GATE U764 ( .I1(hilo[45]), .I2(n1700), .O(n721) );
  NAND4_GATE U765 ( .I1(n1243), .I2(n1242), .I3(n1241), .I4(n1240), .O(n1410)
         );
  NAND_GATE U766 ( .I1(n52), .I2(n1410), .O(n719) );
  NAND_GATE U767 ( .I1(n91), .I2(n1452), .O(n712) );
  NAND_GATE U768 ( .I1(op2[13]), .I2(n1499), .O(n711) );
  NAND_GATE U769 ( .I1(n712), .I2(n711), .O(n713) );
  NAND_GATE U770 ( .I1(n1456), .I2(n713), .O(n714) );
  NAND_GATE U771 ( .I1(op1[13]), .I2(n714), .O(n718) );
  AND_GATE U772 ( .I1(n719), .I2(n718), .O(n720) );
  AND3_GATE U773 ( .I1(n722), .I2(n721), .I3(n720), .O(n723) );
  NAND4_GATE U774 ( .I1(n726), .I2(n725), .I3(n724), .I4(n723), .O(res[13]) );
  NAND_GATE U775 ( .I1(res_add[14]), .I2(n1691), .O(n755) );
  NAND_GATE U776 ( .I1(hilo[14]), .I2(n178), .O(n754) );
  NAND_GATE U781 ( .I1(n124), .I2(n1694), .O(n727) );
  NAND_GATE U782 ( .I1(n92), .I2(n727), .O(n736) );
  AND_GATE U783 ( .I1(op2[14]), .I2(n12), .O(n729) );
  NAND_GATE U788 ( .I1(n124), .I2(n74), .O(n728) );
  NAND_GATE U789 ( .I1(n729), .I2(n728), .O(n730) );
  NAND_GATE U790 ( .I1(n736), .I2(n730), .O(n753) );
  NAND_GATE U791 ( .I1(n1166), .I2(n1701), .O(n749) );
  NAND_GATE U792 ( .I1(hilo[46]), .I2(n1700), .O(n748) );
  NAND4_GATE U793 ( .I1(n1186), .I2(n1185), .I3(n1184), .I4(n1183), .O(n1460)
         );
  NAND_GATE U794 ( .I1(n52), .I2(n1460), .O(n746) );
  NAND_GATE U800 ( .I1(n92), .I2(n1452), .O(n742) );
  NAND_GATE U801 ( .I1(op2[14]), .I2(n1499), .O(n739) );
  NAND_GATE U802 ( .I1(n742), .I2(n739), .O(n743) );
  NAND_GATE U803 ( .I1(n1456), .I2(n743), .O(n744) );
  NAND_GATE U804 ( .I1(op1[14]), .I2(n744), .O(n745) );
  AND_GATE U805 ( .I1(n746), .I2(n745), .O(n747) );
  AND3_GATE U806 ( .I1(n749), .I2(n748), .I3(n747), .O(n750) );
  NAND4_GATE U807 ( .I1(n755), .I2(n754), .I3(n753), .I4(n750), .O(res[14]) );
  NAND_GATE U808 ( .I1(n399), .I2(n97), .O(n762) );
  NAND_GATE U809 ( .I1(n398), .I2(n98), .O(n761) );
  NAND_GATE U810 ( .I1(n397), .I2(n99), .O(n756) );
  NAND4_GATE U811 ( .I1(n1338), .I2(n762), .I3(n761), .I4(n756), .O(n246) );
  NAND_GATE U812 ( .I1(n399), .I2(n93), .O(n766) );
  NAND_GATE U813 ( .I1(n398), .I2(n94), .O(n765) );
  NAND_GATE U814 ( .I1(n397), .I2(n95), .O(n764) );
  NAND_GATE U815 ( .I1(n396), .I2(n96), .O(n763) );
  NAND4_GATE U816 ( .I1(n766), .I2(n765), .I3(n764), .I4(n763), .O(n245) );
  NAND4_GATE U821 ( .I1(n1132), .I2(n1131), .I3(n1130), .I4(n1129), .O(n432)
         );
  NAND_GATE U822 ( .I1(n432), .I2(n52), .O(n807) );
  NAND_GATE U823 ( .I1(n93), .I2(n1452), .O(n768) );
  NAND_GATE U828 ( .I1(op2[15]), .I2(n1499), .O(n767) );
  NAND_GATE U829 ( .I1(n768), .I2(n767), .O(n769) );
  NAND_GATE U830 ( .I1(n1456), .I2(n769), .O(n770) );
  NAND_GATE U832 ( .I1(op1[15]), .I2(n770), .O(n806) );
  INV_GATE U833 ( .I1(n2051), .O(n2041) );
  NAND3_GATE U834 ( .I1(n11), .I2(n1701), .I3(n794), .O(n785) );
  NAND_GATE U835 ( .I1(n801), .I2(n2046), .O(n782) );
  NAND_GATE U836 ( .I1(n802), .I2(n2047), .O(n773) );
  NAND_GATE U837 ( .I1(n175), .I2(n245), .O(n772) );
  NAND_GATE U838 ( .I1(n167), .I2(n246), .O(n771) );
  NAND5_GATE U839 ( .I1(n782), .I2(n773), .I3(n772), .I4(n1635), .I5(n771), 
        .O(n784) );
  NAND_GATE U841 ( .I1(n1145), .I2(n6), .O(n783) );
  AND3_GATE U842 ( .I1(n785), .I2(n784), .I3(n783), .O(n805) );
  NAND_GATE U843 ( .I1(n125), .I2(n1694), .O(n786) );
  NAND_GATE U844 ( .I1(n93), .I2(n786), .O(n790) );
  AND_GATE U845 ( .I1(op2[15]), .I2(n12), .O(n788) );
  NAND_GATE U846 ( .I1(n125), .I2(n74), .O(n787) );
  NAND_GATE U847 ( .I1(n788), .I2(n787), .O(n789) );
  NAND_GATE U848 ( .I1(n790), .I2(n789), .O(n796) );
  NAND_GATE U849 ( .I1(hilo[15]), .I2(n178), .O(n795) );
  AND_GATE U859 ( .I1(n796), .I2(n795), .O(n804) );
  NAND_GATE U860 ( .I1(res_add[15]), .I2(n1691), .O(n798) );
  NAND_GATE U861 ( .I1(hilo[47]), .I2(n1700), .O(n797) );
  AND_GATE U862 ( .I1(n798), .I2(n797), .O(n803) );
  NAND5_GATE U863 ( .I1(n807), .I2(n806), .I3(n805), .I4(n804), .I5(n803), .O(
        res[15]) );
  NAND_GATE U866 ( .I1(res_add[16]), .I2(n1691), .O(n850) );
  NAND_GATE U867 ( .I1(hilo[16]), .I2(n178), .O(n849) );
  NAND_GATE U868 ( .I1(n126), .I2(n1694), .O(n808) );
  NAND_GATE U869 ( .I1(n94), .I2(n808), .O(n812) );
  AND_GATE U870 ( .I1(op2[16]), .I2(n12), .O(n810) );
  NAND_GATE U874 ( .I1(n126), .I2(n74), .O(n809) );
  NAND_GATE U875 ( .I1(n810), .I2(n809), .O(n811) );
  NAND_GATE U876 ( .I1(n812), .I2(n811), .O(n848) );
  NAND_GATE U878 ( .I1(n740), .I2(n17), .O(n815) );
  NAND_GATE U879 ( .I1(n589), .I2(n13), .O(n814) );
  NAND_GATE U880 ( .I1(hilo[48]), .I2(n1700), .O(n813) );
  AND3_GATE U881 ( .I1(n815), .I2(n814), .I3(n813), .O(n847) );
  INV_GATE U882 ( .I1(n1457), .O(n2048) );
  NAND_GATE U883 ( .I1(n114), .I2(n6), .O(n876) );
  NAND_GATE U889 ( .I1(n1512), .I2(n876), .O(n824) );
  NAND_GATE U890 ( .I1(n2048), .I2(n824), .O(n845) );
  NAND_GATE U891 ( .I1(n53), .I2(n16), .O(n830) );
  NAND_GATE U892 ( .I1(n94), .I2(n1452), .O(n826) );
  NAND_GATE U893 ( .I1(op2[16]), .I2(n1499), .O(n825) );
  NAND_GATE U894 ( .I1(n826), .I2(n825), .O(n827) );
  NAND_GATE U895 ( .I1(n1456), .I2(n827), .O(n828) );
  NAND_GATE U896 ( .I1(op1[16]), .I2(n828), .O(n829) );
  AND_GATE U897 ( .I1(n830), .I2(n829), .O(n839) );
  NAND_GATE U898 ( .I1(n738), .I2(n14), .O(n837) );
  NAND_GATE U899 ( .I1(n741), .I2(n15), .O(n836) );
  NAND3_GATE U900 ( .I1(ctrl[6]), .I2(n60), .I3(n31), .O(n831) );
  NOR_GATE U901 ( .I1(ctrl[9]), .I2(n831), .O(n1508) );
  NAND_GATE U902 ( .I1(op2[0]), .I2(n1508), .O(n832) );
  AND3_GATE U903 ( .I1(n837), .I2(n836), .I3(n832), .O(n838) );
  AND4_GATE U904 ( .I1(n2050), .I2(n845), .I3(n839), .I4(n838), .O(n846) );
  NAND5_GATE U905 ( .I1(n850), .I2(n849), .I3(n848), .I4(n847), .I5(n846), .O(
        res[16]) );
  NAND_GATE U910 ( .I1(res_add[17]), .I2(n1691), .O(n889) );
  NAND_GATE U911 ( .I1(hilo[17]), .I2(n178), .O(n888) );
  NAND_GATE U912 ( .I1(n127), .I2(n1694), .O(n851) );
  NAND_GATE U917 ( .I1(n95), .I2(n851), .O(n855) );
  AND_GATE U918 ( .I1(op2[17]), .I2(n12), .O(n853) );
  NAND_GATE U919 ( .I1(n127), .I2(n74), .O(n852) );
  NAND_GATE U920 ( .I1(n853), .I2(n852), .O(n854) );
  NAND_GATE U921 ( .I1(n855), .I2(n854), .O(n887) );
  NAND_GATE U922 ( .I1(n698), .I2(n17), .O(n865) );
  NAND_GATE U923 ( .I1(n945), .I2(n1635), .O(n864) );
  NAND_GATE U929 ( .I1(n556), .I2(n13), .O(n857) );
  NAND_GATE U930 ( .I1(hilo[49]), .I2(n1700), .O(n856) );
  AND4_GATE U931 ( .I1(n865), .I2(n864), .I3(n857), .I4(n856), .O(n886) );
  NAND_GATE U932 ( .I1(n95), .I2(n1452), .O(n867) );
  NAND_GATE U933 ( .I1(op2[17]), .I2(n1499), .O(n866) );
  NAND_GATE U934 ( .I1(n867), .I2(n866), .O(n868) );
  NAND_GATE U935 ( .I1(n1456), .I2(n868), .O(n869) );
  NAND_GATE U936 ( .I1(op1[17]), .I2(n869), .O(n884) );
  NAND_GATE U937 ( .I1(n694), .I2(n14), .O(n883) );
  NAND_GATE U938 ( .I1(n696), .I2(n16), .O(n870) );
  AND_GATE U939 ( .I1(n2050), .I2(n870), .O(n879) );
  NAND_GATE U940 ( .I1(n699), .I2(n15), .O(n872) );
  NAND_GATE U941 ( .I1(op2[1]), .I2(n1508), .O(n871) );
  AND_GATE U942 ( .I1(n872), .I2(n871), .O(n878) );
  INV_GATE U943 ( .I1(n876), .O(n1303) );
  NAND_GATE U944 ( .I1(n964), .I2(n1303), .O(n877) );
  AND5_GATE U945 ( .I1(n884), .I2(n883), .I3(n879), .I4(n878), .I5(n877), .O(
        n885) );
  NAND5_GATE U951 ( .I1(n889), .I2(n888), .I3(n887), .I4(n886), .I5(n885), .O(
        res[17]) );
  NAND_GATE U952 ( .I1(res_add[18]), .I2(n1691), .O(n930) );
  NAND_GATE U953 ( .I1(hilo[18]), .I2(n178), .O(n929) );
  NAND_GATE U959 ( .I1(n128), .I2(n1694), .O(n890) );
  NAND_GATE U960 ( .I1(n96), .I2(n890), .O(n894) );
  AND_GATE U961 ( .I1(op2[18]), .I2(n12), .O(n892) );
  NAND_GATE U962 ( .I1(n128), .I2(n74), .O(n891) );
  NAND_GATE U963 ( .I1(n892), .I2(n891), .O(n893) );
  NAND_GATE U964 ( .I1(n894), .I2(n893), .O(n928) );
  NAND_GATE U965 ( .I1(n823), .I2(n17), .O(n902) );
  NAND_GATE U971 ( .I1(n507), .I2(n1635), .O(n901) );
  NAND_GATE U972 ( .I1(n468), .I2(n13), .O(n900) );
  NAND_GATE U973 ( .I1(hilo[50]), .I2(n1700), .O(n895) );
  AND4_GATE U974 ( .I1(n902), .I2(n901), .I3(n900), .I4(n895), .O(n927) );
  NAND_GATE U975 ( .I1(n96), .I2(n1452), .O(n904) );
  NAND_GATE U976 ( .I1(op2[18]), .I2(n1499), .O(n903) );
  NAND_GATE U977 ( .I1(n904), .I2(n903), .O(n905) );
  NAND_GATE U978 ( .I1(n1456), .I2(n905), .O(n906) );
  NAND_GATE U979 ( .I1(op1[18]), .I2(n906), .O(n925) );
  NAND_GATE U980 ( .I1(n822), .I2(n14), .O(n924) );
  NAND_GATE U981 ( .I1(n493), .I2(n16), .O(n907) );
  AND_GATE U982 ( .I1(n2050), .I2(n907), .O(n915) );
  NAND_GATE U983 ( .I1(n657), .I2(n15), .O(n912) );
  NAND_GATE U984 ( .I1(op2[2]), .I2(n1508), .O(n908) );
  AND_GATE U985 ( .I1(n912), .I2(n908), .O(n914) );
  NAND_GATE U986 ( .I1(n522), .I2(n1303), .O(n913) );
  AND5_GATE U987 ( .I1(n925), .I2(n924), .I3(n915), .I4(n914), .I5(n913), .O(
        n926) );
  NAND5_GATE U993 ( .I1(n930), .I2(n929), .I3(n928), .I4(n927), .I5(n926), .O(
        res[18]) );
  NAND_GATE U994 ( .I1(res_add[19]), .I2(n1691), .O(n974) );
  NAND_GATE U995 ( .I1(hilo[19]), .I2(n178), .O(n973) );
  NAND_GATE U1001 ( .I1(n129), .I2(n1694), .O(n935) );
  NAND_GATE U1002 ( .I1(n97), .I2(n935), .O(n939) );
  AND_GATE U1003 ( .I1(op2[19]), .I2(n12), .O(n937) );
  NAND_GATE U1004 ( .I1(n129), .I2(n74), .O(n936) );
  NAND_GATE U1005 ( .I1(n937), .I2(n936), .O(n938) );
  NAND_GATE U1006 ( .I1(n939), .I2(n938), .O(n972) );
  NAND_GATE U1007 ( .I1(n781), .I2(n17), .O(n943) );
  NAND_GATE U1008 ( .I1(n379), .I2(n1635), .O(n942) );
  NAND_GATE U1009 ( .I1(n430), .I2(n13), .O(n941) );
  NAND_GATE U1010 ( .I1(hilo[51]), .I2(n1700), .O(n940) );
  AND4_GATE U1011 ( .I1(n943), .I2(n942), .I3(n941), .I4(n940), .O(n971) );
  NAND_GATE U1017 ( .I1(n97), .I2(n1452), .O(n956) );
  NAND_GATE U1018 ( .I1(op2[19]), .I2(n1499), .O(n944) );
  NAND_GATE U1019 ( .I1(n956), .I2(n944), .O(n957) );
  NAND_GATE U1020 ( .I1(n1456), .I2(n957), .O(n958) );
  NAND_GATE U1021 ( .I1(op1[19]), .I2(n958), .O(n969) );
  NAND_GATE U1022 ( .I1(n780), .I2(n14), .O(n968) );
  NAND_GATE U1023 ( .I1(n361), .I2(n16), .O(n959) );
  AND_GATE U1024 ( .I1(n2050), .I2(n959), .O(n966) );
  NAND_GATE U1025 ( .I1(n619), .I2(n15), .O(n961) );
  NAND_GATE U1026 ( .I1(op2[3]), .I2(n1508), .O(n960) );
  AND_GATE U1027 ( .I1(n961), .I2(n960), .O(n963) );
  NAND_GATE U1028 ( .I1(n400), .I2(n1303), .O(n962) );
  AND5_GATE U1029 ( .I1(n969), .I2(n968), .I3(n966), .I4(n963), .I5(n962), .O(
        n970) );
  NAND5_GATE U1030 ( .I1(n974), .I2(n973), .I3(n972), .I4(n971), .I5(n970), 
        .O(res[19]) );
  NAND_GATE U1031 ( .I1(res_add[20]), .I2(n1691), .O(n1011) );
  NAND_GATE U1032 ( .I1(hilo[20]), .I2(n178), .O(n1010) );
  NAND_GATE U1033 ( .I1(n130), .I2(n1694), .O(n975) );
  NAND_GATE U1034 ( .I1(n98), .I2(n975), .O(n979) );
  AND_GATE U1035 ( .I1(op2[20]), .I2(n12), .O(n977) );
  NAND_GATE U1036 ( .I1(n130), .I2(n74), .O(n976) );
  NAND_GATE U1037 ( .I1(n977), .I2(n976), .O(n978) );
  NAND_GATE U1038 ( .I1(n979), .I2(n978), .O(n1009) );
  NAND_GATE U1039 ( .I1(n741), .I2(n17), .O(n987) );
  NAND_GATE U1040 ( .I1(n341), .I2(n1635), .O(n986) );
  NAND_GATE U1041 ( .I1(n588), .I2(n13), .O(n981) );
  NAND_GATE U1042 ( .I1(hilo[52]), .I2(n1700), .O(n980) );
  AND4_GATE U1043 ( .I1(n987), .I2(n986), .I3(n981), .I4(n980), .O(n1008) );
  NAND_GATE U1044 ( .I1(n98), .I2(n1452), .O(n989) );
  NAND_GATE U1045 ( .I1(op2[20]), .I2(n1499), .O(n988) );
  NAND_GATE U1046 ( .I1(n989), .I2(n988), .O(n990) );
  NAND_GATE U1047 ( .I1(n1456), .I2(n990), .O(n991) );
  NAND_GATE U1048 ( .I1(op1[20]), .I2(n991), .O(n1006) );
  NAND_GATE U1049 ( .I1(n740), .I2(n14), .O(n1001) );
  NAND_GATE U1050 ( .I1(n51), .I2(n7), .O(n992) );
  AND_GATE U1051 ( .I1(n2050), .I2(n992), .O(n1000) );
  NAND_GATE U1052 ( .I1(n589), .I2(n15), .O(n994) );
  NAND_GATE U1053 ( .I1(op2[4]), .I2(n1508), .O(n993) );
  AND_GATE U1063 ( .I1(n994), .I2(n993), .O(n999) );
  NAND_GATE U1064 ( .I1(n340), .I2(n1303), .O(n998) );
  AND5_GATE U1065 ( .I1(n1006), .I2(n1001), .I3(n1000), .I4(n999), .I5(n998), 
        .O(n1007) );
  NAND5_GATE U1066 ( .I1(n1011), .I2(n1010), .I3(n1009), .I4(n1008), .I5(n1007), .O(res[20]) );
  NAND_GATE U1067 ( .I1(res_add[21]), .I2(n1691), .O(n1050) );
  NAND_GATE U1068 ( .I1(hilo[21]), .I2(n178), .O(n1049) );
  NAND_GATE U1069 ( .I1(n131), .I2(n1694), .O(n1012) );
  NAND_GATE U1070 ( .I1(n99), .I2(n1012), .O(n1016) );
  AND_GATE U1076 ( .I1(op2[21]), .I2(n12), .O(n1014) );
  NAND_GATE U1077 ( .I1(n131), .I2(n74), .O(n1013) );
  NAND_GATE U1078 ( .I1(n1014), .I2(n1013), .O(n1015) );
  NAND_GATE U1079 ( .I1(n1016), .I2(n1015), .O(n1048) );
  NAND_GATE U1080 ( .I1(n699), .I2(n17), .O(n1024) );
  NAND_GATE U1081 ( .I1(n311), .I2(n1635), .O(n1019) );
  NAND_GATE U1082 ( .I1(n555), .I2(n13), .O(n1018) );
  NAND_GATE U1083 ( .I1(hilo[53]), .I2(n1700), .O(n1017) );
  AND4_GATE U1084 ( .I1(n1024), .I2(n1019), .I3(n1018), .I4(n1017), .O(n1047)
         );
  NAND_GATE U1085 ( .I1(op2[5]), .I2(n1508), .O(n1041) );
  NAND_GATE U1086 ( .I1(n310), .I2(n1303), .O(n1040) );
  NAND_GATE U1087 ( .I1(n316), .I2(n51), .O(n1039) );
  NAND_GATE U1088 ( .I1(n99), .I2(n1452), .O(n1026) );
  NAND_GATE U1089 ( .I1(op2[21]), .I2(n1499), .O(n1025) );
  NAND_GATE U1090 ( .I1(n1026), .I2(n1025), .O(n1027) );
  NAND_GATE U1091 ( .I1(n1456), .I2(n1027), .O(n1028) );
  NAND_GATE U1092 ( .I1(op1[21]), .I2(n1028), .O(n1032) );
  NAND_GATE U1093 ( .I1(n698), .I2(n14), .O(n1030) );
  NAND_GATE U1094 ( .I1(n556), .I2(n15), .O(n1029) );
  AND_GATE U1104 ( .I1(n1030), .I2(n1029), .O(n1031) );
  AND3_GATE U1105 ( .I1(n2050), .I2(n1032), .I3(n1031), .O(n1038) );
  AND4_GATE U1106 ( .I1(n1041), .I2(n1040), .I3(n1039), .I4(n1038), .O(n1046)
         );
  NAND5_GATE U1107 ( .I1(n1050), .I2(n1049), .I3(n1048), .I4(n1047), .I5(n1046), .O(res[21]) );
  NAND_GATE U1108 ( .I1(res_add[22]), .I2(n1691), .O(n1088) );
  NAND_GATE U1109 ( .I1(hilo[22]), .I2(n178), .O(n1087) );
  NAND_GATE U1110 ( .I1(n132), .I2(n1694), .O(n1051) );
  NAND_GATE U1111 ( .I1(n100), .I2(n1051), .O(n1055) );
  AND_GATE U1112 ( .I1(op2[22]), .I2(n12), .O(n1053) );
  NAND_GATE U1113 ( .I1(n132), .I2(n74), .O(n1052) );
  NAND_GATE U1114 ( .I1(n1053), .I2(n1052), .O(n1054) );
  NAND_GATE U1124 ( .I1(n1055), .I2(n1054), .O(n1086) );
  NAND_GATE U1125 ( .I1(n657), .I2(n17), .O(n1063) );
  NAND_GATE U1126 ( .I1(n281), .I2(n1635), .O(n1058) );
  NAND_GATE U1127 ( .I1(n467), .I2(n13), .O(n1057) );
  NAND_GATE U1128 ( .I1(hilo[54]), .I2(n1700), .O(n1056) );
  AND4_GATE U1129 ( .I1(n1063), .I2(n1058), .I3(n1057), .I4(n1056), .O(n1085)
         );
  NAND_GATE U1130 ( .I1(op2[6]), .I2(n1508), .O(n1079) );
  NAND_GATE U1131 ( .I1(n280), .I2(n1303), .O(n1078) );
  NAND_GATE U1132 ( .I1(n286), .I2(n51), .O(n1077) );
  NAND_GATE U1133 ( .I1(n100), .I2(n1452), .O(n1065) );
  NAND_GATE U1138 ( .I1(op2[22]), .I2(n1499), .O(n1064) );
  NAND_GATE U1139 ( .I1(n1065), .I2(n1064), .O(n1066) );
  NAND_GATE U1140 ( .I1(n1456), .I2(n1066), .O(n1067) );
  NAND_GATE U1141 ( .I1(op1[22]), .I2(n1067), .O(n1071) );
  NAND_GATE U1142 ( .I1(n823), .I2(n14), .O(n1069) );
  NAND_GATE U1150 ( .I1(n468), .I2(n15), .O(n1068) );
  AND_GATE U1154 ( .I1(n1069), .I2(n1068), .O(n1070) );
  AND3_GATE U1156 ( .I1(n2050), .I2(n1071), .I3(n1070), .O(n1076) );
  AND4_GATE U1160 ( .I1(n1079), .I2(n1078), .I3(n1077), .I4(n1076), .O(n1084)
         );
  NAND5_GATE U1161 ( .I1(n1088), .I2(n1087), .I3(n1086), .I4(n1085), .I5(n1084), .O(res[22]) );
  NAND_GATE U1162 ( .I1(res_add[23]), .I2(n1691), .O(n1118) );
  NAND_GATE U1163 ( .I1(hilo[23]), .I2(n178), .O(n1117) );
  NAND_GATE U1164 ( .I1(n133), .I2(n1694), .O(n1089) );
  NAND_GATE U1170 ( .I1(n101), .I2(n1089), .O(n1093) );
  AND_GATE U1171 ( .I1(op2[23]), .I2(n12), .O(n1091) );
  NAND_GATE U1172 ( .I1(n133), .I2(n74), .O(n1090) );
  NAND_GATE U1173 ( .I1(n1091), .I2(n1090), .O(n1092) );
  NAND_GATE U1174 ( .I1(n1093), .I2(n1092), .O(n1116) );
  NAND_GATE U1175 ( .I1(n619), .I2(n17), .O(n1101) );
  NAND_GATE U1176 ( .I1(n248), .I2(n1635), .O(n1100) );
  NAND_GATE U1177 ( .I1(n429), .I2(n13), .O(n1095) );
  NAND_GATE U1178 ( .I1(hilo[55]), .I2(n1700), .O(n1094) );
  AND4_GATE U1179 ( .I1(n1101), .I2(n1100), .I3(n1095), .I4(n1094), .O(n1115)
         );
  NAND_GATE U1180 ( .I1(op2[7]), .I2(n1508), .O(n1113) );
  NAND_GATE U1203 ( .I1(n247), .I2(n1303), .O(n1112) );
  NAND_GATE U1204 ( .I1(n253), .I2(n51), .O(n1111) );
  NAND_GATE U1205 ( .I1(n101), .I2(n1452), .O(n1103) );
  NAND_GATE U1206 ( .I1(op2[23]), .I2(n1499), .O(n1102) );
  NAND_GATE U1207 ( .I1(n1103), .I2(n1102), .O(n1104) );
  NAND_GATE U1208 ( .I1(n1456), .I2(n1104), .O(n1105) );
  NAND_GATE U1209 ( .I1(op1[23]), .I2(n1105), .O(n1109) );
  NAND_GATE U1210 ( .I1(n781), .I2(n14), .O(n1107) );
  NAND_GATE U1211 ( .I1(n430), .I2(n15), .O(n1106) );
  AND_GATE U1212 ( .I1(n1107), .I2(n1106), .O(n1108) );
  AND3_GATE U1234 ( .I1(n2050), .I2(n1109), .I3(n1108), .O(n1110) );
  AND4_GATE U1235 ( .I1(n1113), .I2(n1112), .I3(n1111), .I4(n1110), .O(n1114)
         );
  NAND5_GATE U1236 ( .I1(n1118), .I2(n1117), .I3(n1116), .I4(n1115), .I5(n1114), .O(res[23]) );
  NAND_GATE U1239 ( .I1(res_add[24]), .I2(n1691), .O(n1158) );
  NAND_GATE U1240 ( .I1(hilo[24]), .I2(n178), .O(n1157) );
  NAND_GATE U1241 ( .I1(n134), .I2(n1694), .O(n1119) );
  NAND_GATE U1246 ( .I1(n102), .I2(n1119), .O(n1123) );
  AND_GATE U1247 ( .I1(op2[24]), .I2(n12), .O(n1121) );
  NAND_GATE U1248 ( .I1(n134), .I2(n74), .O(n1120) );
  NAND_GATE U1249 ( .I1(n1121), .I2(n1120), .O(n1122) );
  NAND_GATE U1250 ( .I1(n1123), .I2(n1122), .O(n1156) );
  NAND_GATE U1251 ( .I1(n589), .I2(n17), .O(n1127) );
  NAND_GATE U1252 ( .I1(n216), .I2(n1635), .O(n1126) );
  NAND_GATE U1253 ( .I1(n590), .I2(n13), .O(n1125) );
  NAND_GATE U1254 ( .I1(hilo[56]), .I2(n1700), .O(n1124) );
  AND4_GATE U1255 ( .I1(n1127), .I2(n1126), .I3(n1125), .I4(n1124), .O(n1155)
         );
  NAND_GATE U1256 ( .I1(op2[8]), .I2(n1508), .O(n1153) );
  NAND_GATE U1257 ( .I1(n215), .I2(n1303), .O(n1152) );
  NAND_GATE U1258 ( .I1(n1128), .I2(n51), .O(n1151) );
  NAND_GATE U1259 ( .I1(n102), .I2(n1452), .O(n1138) );
  NAND_GATE U1260 ( .I1(op2[24]), .I2(n1499), .O(n1137) );
  NAND_GATE U1261 ( .I1(n1138), .I2(n1137), .O(n1139) );
  NAND_GATE U1262 ( .I1(n1456), .I2(n1139), .O(n1140) );
  NAND_GATE U1263 ( .I1(op1[24]), .I2(n1140), .O(n1144) );
  NAND_GATE U1264 ( .I1(n741), .I2(n14), .O(n1142) );
  NAND_GATE U1265 ( .I1(n588), .I2(n15), .O(n1141) );
  AND_GATE U1268 ( .I1(n1142), .I2(n1141), .O(n1143) );
  AND3_GATE U1269 ( .I1(n2050), .I2(n1144), .I3(n1143), .O(n1150) );
  AND4_GATE U1270 ( .I1(n1153), .I2(n1152), .I3(n1151), .I4(n1150), .O(n1154)
         );
  NAND5_GATE U1271 ( .I1(n1158), .I2(n1157), .I3(n1156), .I4(n1155), .I5(n1154), .O(res[24]) );
  NAND_GATE U1272 ( .I1(res_add[25]), .I2(n1691), .O(n1212) );
  NAND_GATE U1285 ( .I1(hilo[25]), .I2(n178), .O(n1202) );
  NAND_GATE U1287 ( .I1(n135), .I2(n1694), .O(n1159) );
  NAND_GATE U1288 ( .I1(n103), .I2(n1159), .O(n1163) );
  AND_GATE U1289 ( .I1(op2[25]), .I2(n12), .O(n1161) );
  NAND_GATE U1291 ( .I1(n135), .I2(n74), .O(n1160) );
  NAND_GATE U1292 ( .I1(n1161), .I2(n1160), .O(n1162) );
  NAND_GATE U1293 ( .I1(n1163), .I2(n1162), .O(n1201) );
  NAND_GATE U1294 ( .I1(n556), .I2(n17), .O(n1177) );
  NAND_GATE U1295 ( .I1(n177), .I2(n1635), .O(n1176) );
  NAND_GATE U1306 ( .I1(n557), .I2(n13), .O(n1165) );
  NAND_GATE U1307 ( .I1(hilo[57]), .I2(n1700), .O(n1164) );
  AND4_GATE U1308 ( .I1(n1177), .I2(n1176), .I3(n1165), .I4(n1164), .O(n1200)
         );
  NAND_GATE U1309 ( .I1(n103), .I2(n1452), .O(n1179) );
  NAND_GATE U1310 ( .I1(op2[25]), .I2(n1499), .O(n1178) );
  NAND_GATE U1311 ( .I1(n1179), .I2(n1178), .O(n1180) );
  NAND_GATE U1312 ( .I1(n1456), .I2(n1180), .O(n1181) );
  NAND_GATE U1313 ( .I1(op1[25]), .I2(n1181), .O(n1198) );
  NAND_GATE U1314 ( .I1(n699), .I2(n14), .O(n1197) );
  NAND_GATE U1315 ( .I1(n1182), .I2(n51), .O(n1191) );
  AND_GATE U1316 ( .I1(n2050), .I2(n1191), .O(n1196) );
  NAND_GATE U1335 ( .I1(n555), .I2(n15), .O(n1193) );
  NAND_GATE U1336 ( .I1(op2[9]), .I2(n1508), .O(n1192) );
  AND_GATE U1337 ( .I1(n1193), .I2(n1192), .O(n1195) );
  NAND_GATE U1338 ( .I1(n174), .I2(n1303), .O(n1194) );
  AND5_GATE U1339 ( .I1(n1198), .I2(n1197), .I3(n1196), .I4(n1195), .I5(n1194), 
        .O(n1199) );
  NAND5_GATE U1340 ( .I1(n1212), .I2(n1202), .I3(n1201), .I4(n1200), .I5(n1199), .O(res[25]) );
  NAND_GATE U1341 ( .I1(res_add[26]), .I2(n1691), .O(n1269) );
  NAND_GATE U1342 ( .I1(hilo[26]), .I2(n178), .O(n1268) );
  NAND_GATE U1343 ( .I1(n136), .I2(n1694), .O(n1213) );
  NAND_GATE U1344 ( .I1(n104), .I2(n1213), .O(n1226) );
  AND_GATE U1348 ( .I1(op2[26]), .I2(n12), .O(n1215) );
  NAND_GATE U1349 ( .I1(n136), .I2(n74), .O(n1214) );
  NAND_GATE U1350 ( .I1(n1215), .I2(n1214), .O(n1220) );
  NAND_GATE U1351 ( .I1(n1226), .I2(n1220), .O(n1267) );
  NAND_GATE U1352 ( .I1(n468), .I2(n17), .O(n1233) );
  NAND_GATE U1354 ( .I1(n672), .I2(n1635), .O(n1229) );
  NAND_GATE U1355 ( .I1(n469), .I2(n13), .O(n1228) );
  NAND_GATE U1356 ( .I1(hilo[58]), .I2(n1700), .O(n1227) );
  AND4_GATE U1357 ( .I1(n1233), .I2(n1229), .I3(n1228), .I4(n1227), .O(n1266)
         );
  NAND_GATE U1358 ( .I1(n104), .I2(n1452), .O(n1235) );
  NAND_GATE U1372 ( .I1(op2[26]), .I2(n1499), .O(n1234) );
  NAND_GATE U1374 ( .I1(n1235), .I2(n1234), .O(n1236) );
  NAND_GATE U1375 ( .I1(n1456), .I2(n1236), .O(n1237) );
  NAND_GATE U1376 ( .I1(op1[26]), .I2(n1237), .O(n1264) );
  NAND_GATE U1377 ( .I1(n657), .I2(n14), .O(n1263) );
  NAND_GATE U1378 ( .I1(n1238), .I2(n51), .O(n1239) );
  AND_GATE U1380 ( .I1(n2050), .I2(n1239), .O(n1262) );
  NAND_GATE U1389 ( .I1(n467), .I2(n15), .O(n1259) );
  NAND_GATE U1390 ( .I1(op2[10]), .I2(n1508), .O(n1258) );
  AND_GATE U1391 ( .I1(n1259), .I2(n1258), .O(n1261) );
  NAND_GATE U1392 ( .I1(n667), .I2(n1303), .O(n1260) );
  AND5_GATE U1393 ( .I1(n1264), .I2(n1263), .I3(n1262), .I4(n1261), .I5(n1260), 
        .O(n1265) );
  NAND5_GATE U1394 ( .I1(n1269), .I2(n1268), .I3(n1267), .I4(n1266), .I5(n1265), .O(res[26]) );
  NAND_GATE U1395 ( .I1(res_add[27]), .I2(n1691), .O(n1326) );
  NAND_GATE U1396 ( .I1(hilo[27]), .I2(n178), .O(n1325) );
  NAND_GATE U1397 ( .I1(n137), .I2(n1694), .O(n1287) );
  NAND_GATE U1398 ( .I1(n105), .I2(n1287), .O(n1297) );
  AND_GATE U1399 ( .I1(op2[27]), .I2(n12), .O(n1289) );
  NAND_GATE U1400 ( .I1(n137), .I2(n74), .O(n1288) );
  NAND_GATE U1401 ( .I1(n1289), .I2(n1288), .O(n1296) );
  NAND_GATE U1419 ( .I1(n1297), .I2(n1296), .O(n1324) );
  NAND_GATE U1420 ( .I1(n430), .I2(n17), .O(n1301) );
  NAND_GATE U1421 ( .I1(n631), .I2(n1635), .O(n1300) );
  NAND_GATE U1422 ( .I1(n431), .I2(n13), .O(n1299) );
  NAND_GATE U1423 ( .I1(hilo[59]), .I2(n1700), .O(n1298) );
  AND4_GATE U1424 ( .I1(n1301), .I2(n1300), .I3(n1299), .I4(n1298), .O(n1317)
         );
  AND_GATE U1425 ( .I1(n632), .I2(n113), .O(n1302) );
  NAND_GATE U1426 ( .I1(n1303), .I2(n1302), .O(n1315) );
  NAND_GATE U1427 ( .I1(n1304), .I2(n51), .O(n1314) );
  NAND_GATE U1428 ( .I1(n105), .I2(n1452), .O(n1306) );
  NAND_GATE U1429 ( .I1(op2[27]), .I2(n1499), .O(n1305) );
  NAND_GATE U1430 ( .I1(n1306), .I2(n1305), .O(n1307) );
  NAND_GATE U1431 ( .I1(n1456), .I2(n1307), .O(n1308) );
  NAND_GATE U1432 ( .I1(op1[27]), .I2(n1308), .O(n1313) );
  NAND_GATE U1434 ( .I1(n619), .I2(n14), .O(n1311) );
  NAND_GATE U1435 ( .I1(n429), .I2(n15), .O(n1310) );
  NAND_GATE U1436 ( .I1(op2[11]), .I2(n1508), .O(n1309) );
  AND3_GATE U1437 ( .I1(n1311), .I2(n1310), .I3(n1309), .O(n1312) );
  AND5_GATE U1438 ( .I1(n2050), .I2(n1315), .I3(n1314), .I4(n1313), .I5(n1312), 
        .O(n1316) );
  NAND5_GATE U1451 ( .I1(n1326), .I2(n1325), .I3(n1324), .I4(n1317), .I5(n1316), .O(res[27]) );
  NAND_GATE U1452 ( .I1(hilo[60]), .I2(n1700), .O(n1336) );
  NAND_GATE U1453 ( .I1(op2[12]), .I2(n1508), .O(n1335) );
  NAND_GATE U1454 ( .I1(res_add[28]), .I2(n1691), .O(n1327) );
  AND3_GATE U1455 ( .I1(n1336), .I2(n1335), .I3(n1327), .O(n1381) );
  NAND_GATE U1459 ( .I1(n106), .I2(n1452), .O(n1339) );
  NAND_GATE U1460 ( .I1(op2[28]), .I2(n1499), .O(n1337) );
  NAND_GATE U1461 ( .I1(n1339), .I2(n1337), .O(n1340) );
  NAND_GATE U1462 ( .I1(n1456), .I2(n1340), .O(n1341) );
  NAND_GATE U1463 ( .I1(op1[28]), .I2(n1341), .O(n1379) );
  NAND4_GATE U1466 ( .I1(n581), .I2(n580), .I3(n582), .I4(n583), .O(n1342) );
  NAND_GATE U1467 ( .I1(n1507), .I2(n1342), .O(n1378) );
  INV_GATE U1468 ( .I1(n175), .O(n1349) );
  NAND_GATE U1469 ( .I1(n1349), .I2(n1635), .O(n1476) );
  NAND_GATE U1470 ( .I1(n1350), .I2(n51), .O(n1368) );
  INV_GATE U1488 ( .I1(n760), .O(n2049) );
  NAND_GATE U1489 ( .I1(n175), .I2(n6), .O(n1417) );
  NAND_GATE U1490 ( .I1(n1512), .I2(n1417), .O(n1351) );
  NAND_GATE U1491 ( .I1(n2049), .I2(n1351), .O(n1352) );
  AND_GATE U1492 ( .I1(n1368), .I2(n1352), .O(n1377) );
  NAND_GATE U1494 ( .I1(n138), .I2(n1694), .O(n1369) );
  NAND_GATE U1499 ( .I1(n106), .I2(n1369), .O(n1373) );
  AND_GATE U1501 ( .I1(op2[28]), .I2(n12), .O(n1371) );
  NAND_GATE U1503 ( .I1(n138), .I2(n74), .O(n1370) );
  NAND_GATE U1504 ( .I1(n1371), .I2(n1370), .O(n1372) );
  NAND_GATE U1505 ( .I1(n1373), .I2(n1372), .O(n1375) );
  NAND_GATE U1506 ( .I1(hilo[28]), .I2(n178), .O(n1374) );
  AND_GATE U1507 ( .I1(n1375), .I2(n1374), .O(n1376) );
  AND5_GATE U1508 ( .I1(n1379), .I2(n1378), .I3(n1476), .I4(n1377), .I5(n1376), 
        .O(n1380) );
  NAND_GATE U1509 ( .I1(n1381), .I2(n1380), .O(res[28]) );
  NAND_GATE U1510 ( .I1(n1225), .I2(n1224), .O(n563) );
  NAND_GATE U1511 ( .I1(n139), .I2(n1694), .O(n1382) );
  NAND_GATE U1512 ( .I1(n107), .I2(n1382), .O(n1394) );
  AND_GATE U1513 ( .I1(op2[29]), .I2(n12), .O(n1392) );
  NAND_GATE U1515 ( .I1(n139), .I2(n74), .O(n1391) );
  NAND_GATE U1518 ( .I1(n1392), .I2(n1391), .O(n1393) );
  NAND_GATE U1519 ( .I1(n1394), .I2(n1393), .O(n1396) );
  NAND_GATE U1520 ( .I1(hilo[29]), .I2(n178), .O(n1395) );
  AND_GATE U1521 ( .I1(n1396), .I2(n1395), .O(n1443) );
  NAND_GATE U1522 ( .I1(n107), .I2(n1452), .O(n1398) );
  NAND_GATE U1523 ( .I1(op2[29]), .I2(n1499), .O(n1397) );
  NAND_GATE U1524 ( .I1(n1398), .I2(n1397), .O(n1407) );
  NAND_GATE U1525 ( .I1(n1456), .I2(n1407), .O(n1408) );
  NAND_GATE U1526 ( .I1(op1[29]), .I2(n1408), .O(n1437) );
  NAND4_GATE U1527 ( .I1(n548), .I2(n547), .I3(n549), .I4(n550), .O(n1409) );
  NAND_GATE U1528 ( .I1(n1507), .I2(n1409), .O(n1436) );
  NAND_GATE U1529 ( .I1(op2[13]), .I2(n1508), .O(n1421) );
  NAND_GATE U1530 ( .I1(n1410), .I2(n51), .O(n1419) );
  INV_GATE U1531 ( .I1(n1417), .O(n1461) );
  NAND_GATE U1532 ( .I1(n562), .I2(n1461), .O(n1418) );
  AND_GATE U1533 ( .I1(n1419), .I2(n1418), .O(n1420) );
  AND5_GATE U1534 ( .I1(n1437), .I2(n1436), .I3(n1421), .I4(n1476), .I5(n1420), 
        .O(n1442) );
  NAND_GATE U1535 ( .I1(hilo[61]), .I2(n1700), .O(n1440) );
  OR_GATE U1536 ( .I1(n1512), .I2(n563), .O(n1439) );
  NAND_GATE U1537 ( .I1(res_add[29]), .I2(n1691), .O(n1438) );
  AND3_GATE U1538 ( .I1(n1440), .I2(n1439), .I3(n1438), .O(n1441) );
  NAND3_GATE U1539 ( .I1(n1443), .I2(n1442), .I3(n1441), .O(res[29]) );
  NAND_GATE U1540 ( .I1(n140), .I2(n1694), .O(n1444) );
  NAND_GATE U1541 ( .I1(n108), .I2(n1444), .O(n1449) );
  AND_GATE U1542 ( .I1(op2[30]), .I2(n12), .O(n1447) );
  NAND_GATE U1543 ( .I1(n140), .I2(n74), .O(n1445) );
  NAND_GATE U1544 ( .I1(n1447), .I2(n1445), .O(n1448) );
  NAND_GATE U1545 ( .I1(n1449), .I2(n1448), .O(n1451) );
  NAND_GATE U1546 ( .I1(hilo[30]), .I2(n178), .O(n1450) );
  AND_GATE U1547 ( .I1(n1451), .I2(n1450), .O(n1485) );
  NAND_GATE U1548 ( .I1(n108), .I2(n1452), .O(n1454) );
  NAND_GATE U1549 ( .I1(op2[30]), .I2(n1499), .O(n1453) );
  NAND_GATE U1550 ( .I1(n1454), .I2(n1453), .O(n1455) );
  NAND_GATE U1551 ( .I1(n1456), .I2(n1455), .O(n1458) );
  NAND_GATE U1552 ( .I1(op1[30]), .I2(n1458), .O(n1479) );
  NAND4_GATE U1553 ( .I1(n460), .I2(n459), .I3(n461), .I4(n462), .O(n1459) );
  NAND_GATE U1554 ( .I1(n1507), .I2(n1459), .O(n1478) );
  NAND_GATE U1555 ( .I1(n399), .I2(n108), .O(n1535) );
  NAND_GATE U1556 ( .I1(n1635), .I2(n1535), .O(n1477) );
  NAND_GATE U1557 ( .I1(n1460), .I2(n51), .O(n1463) );
  NAND_GATE U1558 ( .I1(n479), .I2(n1461), .O(n1462) );
  AND_GATE U1559 ( .I1(n1463), .I2(n1462), .O(n1475) );
  AND5_GATE U1560 ( .I1(n1479), .I2(n1478), .I3(n1477), .I4(n1476), .I5(n1475), 
        .O(n1484) );
  NAND_GATE U1561 ( .I1(hilo[62]), .I2(n1700), .O(n1482) );
  NAND_GATE U1562 ( .I1(op2[14]), .I2(n1508), .O(n1481) );
  NAND_GATE U1563 ( .I1(res_add[30]), .I2(n1691), .O(n1480) );
  AND3_GATE U1564 ( .I1(n1482), .I2(n1481), .I3(n1480), .O(n1483) );
  NAND3_GATE U1565 ( .I1(n1485), .I2(n1484), .I3(n1483), .O(res[30]) );
  NAND_GATE U1566 ( .I1(n141), .I2(n1694), .O(n1486) );
  NAND_GATE U1567 ( .I1(n109), .I2(n1486), .O(n1504) );
  AND_GATE U1568 ( .I1(op2[31]), .I2(n12), .O(n1502) );
  NAND_GATE U1569 ( .I1(op1[31]), .I2(n75), .O(n1501) );
  NAND_GATE U1570 ( .I1(n374), .I2(n1701), .O(n1500) );
  NAND3_GATE U1571 ( .I1(n1502), .I2(n1501), .I3(n1500), .O(n1503) );
  NAND_GATE U1572 ( .I1(n1504), .I2(n1503), .O(n1520) );
  NAND_GATE U1573 ( .I1(hilo[31]), .I2(n178), .O(n1519) );
  NAND_GATE U1574 ( .I1(hilo[63]), .I2(n1700), .O(n1514) );
  NAND_GATE U1575 ( .I1(n419), .I2(n1507), .O(n1513) );
  NAND_GATE U1576 ( .I1(op2[15]), .I2(n1508), .O(n1511) );
  NAND_GATE U1577 ( .I1(op1[31]), .I2(n1509), .O(n1510) );
  AND5_GATE U1578 ( .I1(n1514), .I2(n1513), .I3(n1512), .I4(n1511), .I5(n1510), 
        .O(n1518) );
  NAND_GATE U1579 ( .I1(n417), .I2(n74), .O(n1516) );
  NAND_GATE U1580 ( .I1(res_add[31]), .I2(n1691), .O(n1515) );
  AND_GATE U1581 ( .I1(n1516), .I2(n1515), .O(n1517) );
  NAND4_GATE U1582 ( .I1(n1520), .I2(n1519), .I3(n1518), .I4(n1517), .O(
        res[31]) );
  INV_GATE U1583 ( .I1(efct_op2[31]), .O(n2058) );
  INV_GATE U1584 ( .I1(n1523), .O(n1521) );
  NAND3_GATE U1585 ( .I1(n1525), .I2(n1619), .I3(n8), .O(n1839) );
  INV_GATE U1586 ( .I1(n1524), .O(n1522) );
  NAND_GATE U1587 ( .I1(n1522), .I2(n5), .O(n1840) );
  NAND_GATE U1588 ( .I1(n1839), .I2(n1840), .O(n1697) );
  NAND3_GATE U1589 ( .I1(n1524), .I2(n5), .I3(n1525), .O(n1838) );
  INV_GATE U1590 ( .I1(n1838), .O(n2037) );
  INV_GATE U1591 ( .I1(n1525), .O(n1526) );
  NAND_GATE U1592 ( .I1(n399), .I2(n98), .O(n1528) );
  NAND_GATE U1593 ( .I1(n398), .I2(n99), .O(n1527) );
  NAND4_GATE U1594 ( .I1(n1506), .I2(n1505), .I3(n1528), .I4(n1527), .O(n214)
         );
  NAND_GATE U1595 ( .I1(n398), .I2(n95), .O(n1532) );
  NAND_GATE U1596 ( .I1(n399), .I2(n94), .O(n1531) );
  NAND_GATE U1597 ( .I1(n396), .I2(n97), .O(n1530) );
  NAND_GATE U1598 ( .I1(n397), .I2(n96), .O(n1529) );
  AND4_GATE U1599 ( .I1(n1532), .I2(n1531), .I3(n1530), .I4(n1529), .O(n2035)
         );
  INV_GATE U1600 ( .I1(n1533), .O(n2044) );
  INV_GATE U1601 ( .I1(n1534), .O(n2045) );
  INV_GATE U1602 ( .I1(n1535), .O(n2038) );
  NAND_GATE U1603 ( .I1(n399), .I2(n88), .O(n1539) );
  NAND_GATE U1604 ( .I1(n398), .I2(n89), .O(n1538) );
  NAND_GATE U1605 ( .I1(n397), .I2(n90), .O(n1537) );
  NAND_GATE U1606 ( .I1(n396), .I2(n91), .O(n1536) );
  NAND4_GATE U1607 ( .I1(n1539), .I2(n1538), .I3(n1537), .I4(n1536), .O(n1599)
         );
  INV_GATE U1608 ( .I1(n1599), .O(n2034) );
  NAND_GATE U1609 ( .I1(n399), .I2(n96), .O(n1543) );
  NAND_GATE U1610 ( .I1(n398), .I2(n97), .O(n1542) );
  NAND_GATE U1611 ( .I1(n397), .I2(n98), .O(n1541) );
  NAND_GATE U1612 ( .I1(n396), .I2(n99), .O(n1540) );
  NAND4_GATE U1613 ( .I1(n1543), .I2(n1542), .I3(n1541), .I4(n1540), .O(n279)
         );
  INV_GATE U1614 ( .I1(n279), .O(n2033) );
  NAND_GATE U1615 ( .I1(n399), .I2(n92), .O(n1547) );
  NAND_GATE U1616 ( .I1(n398), .I2(n93), .O(n1546) );
  NAND_GATE U1617 ( .I1(n397), .I2(n94), .O(n1545) );
  NAND_GATE U1618 ( .I1(n396), .I2(n95), .O(n1544) );
  NAND4_GATE U1619 ( .I1(n1547), .I2(n1546), .I3(n1545), .I4(n1544), .O(n278)
         );
  INV_GATE U1620 ( .I1(n278), .O(n2032) );
  INV_GATE U1621 ( .I1(n245), .O(n2039) );
  INV_GATE U1622 ( .I1(n246), .O(n2040) );
  NAND_GATE U1623 ( .I1(n399), .I2(n89), .O(n1551) );
  NAND_GATE U1624 ( .I1(n398), .I2(n90), .O(n1550) );
  NAND_GATE U1625 ( .I1(n397), .I2(n91), .O(n1549) );
  NAND_GATE U1626 ( .I1(n396), .I2(n92), .O(n1548) );
  NAND4_GATE U1627 ( .I1(n1551), .I2(n1550), .I3(n1549), .I4(n1548), .O(n391)
         );
  INV_GATE U1628 ( .I1(n391), .O(n2031) );
  INV_GATE U1629 ( .I1(n214), .O(n2036) );
  NAND_GATE U1630 ( .I1(n399), .I2(n91), .O(n1555) );
  NAND_GATE U1631 ( .I1(n398), .I2(n92), .O(n1554) );
  NAND_GATE U1632 ( .I1(n397), .I2(n93), .O(n1553) );
  NAND_GATE U1633 ( .I1(n396), .I2(n94), .O(n1552) );
  NAND4_GATE U1634 ( .I1(n1555), .I2(n1554), .I3(n1553), .I4(n1552), .O(n1573)
         );
  INV_GATE U1635 ( .I1(n1573), .O(n2030) );
  NAND_GATE U1636 ( .I1(n399), .I2(n99), .O(n1556) );
  NAND4_GATE U1637 ( .I1(n1223), .I2(n1222), .I3(n1221), .I4(n1556), .O(n172)
         );
  INV_GATE U1638 ( .I1(n172), .O(n2029) );
  NAND_GATE U1639 ( .I1(n399), .I2(n95), .O(n1560) );
  NAND_GATE U1640 ( .I1(n398), .I2(n96), .O(n1559) );
  NAND_GATE U1641 ( .I1(n397), .I2(n97), .O(n1558) );
  NAND_GATE U1642 ( .I1(n396), .I2(n98), .O(n1557) );
  NAND4_GATE U1643 ( .I1(n1560), .I2(n1559), .I3(n1558), .I4(n1557), .O(n170)
         );
  INV_GATE U1644 ( .I1(n170), .O(n2028) );
  NAND_GATE U1645 ( .I1(n79), .I2(n74), .O(n1561) );
  NAND_GATE U1646 ( .I1(n1619), .I2(n1561), .O(n967) );
  NAND_GATE U1647 ( .I1(n111), .I2(n74), .O(n1562) );
  NAND_GATE U1648 ( .I1(n1696), .I2(n1562), .O(n965) );
  NAND_GATE U1649 ( .I1(n399), .I2(n83), .O(n1566) );
  NAND_GATE U1650 ( .I1(n398), .I2(n84), .O(n1565) );
  NAND_GATE U1651 ( .I1(n397), .I2(n85), .O(n1564) );
  NAND_GATE U1652 ( .I1(n396), .I2(n86), .O(n1563) );
  NAND4_GATE U1653 ( .I1(n1566), .I2(n1565), .I3(n1564), .I4(n1563), .O(n1572)
         );
  INV_GATE U1654 ( .I1(n1572), .O(n2027) );
  NAND_GATE U1655 ( .I1(n399), .I2(n87), .O(n1570) );
  NAND_GATE U1656 ( .I1(n398), .I2(n88), .O(n1569) );
  NAND_GATE U1657 ( .I1(n397), .I2(n89), .O(n1568) );
  NAND_GATE U1658 ( .I1(n396), .I2(n90), .O(n1567) );
  NAND4_GATE U1659 ( .I1(n1570), .I2(n1569), .I3(n1568), .I4(n1567), .O(n1571)
         );
  INV_GATE U1660 ( .I1(n1571), .O(n2026) );
  NAND_GATE U1661 ( .I1(n2046), .I2(n1571), .O(n1582) );
  NAND_GATE U1662 ( .I1(n167), .I2(n1572), .O(n1575) );
  NAND_GATE U1663 ( .I1(n2047), .I2(n1573), .O(n1574) );
  AND_GATE U1664 ( .I1(n1575), .I2(n1574), .O(n1581) );
  NAND_GATE U1665 ( .I1(n374), .I2(n79), .O(n1579) );
  NAND_GATE U1666 ( .I1(n375), .I2(n80), .O(n1578) );
  NAND_GATE U1667 ( .I1(n377), .I2(n81), .O(n1577) );
  NAND_GATE U1668 ( .I1(n376), .I2(n82), .O(n1576) );
  AND4_GATE U1669 ( .I1(n1579), .I2(n1578), .I3(n1577), .I4(n1576), .O(n1580)
         );
  NAND5_GATE U1670 ( .I1(n934), .I2(n1635), .I3(n1582), .I4(n1581), .I5(n1580), 
        .O(n933) );
  NAND_GATE U1671 ( .I1(hilo[33]), .I2(n1700), .O(n920) );
  NAND_GATE U1672 ( .I1(n111), .I2(n79), .O(n1584) );
  INV_GATE U1673 ( .I1(n1584), .O(n1583) );
  NAND_GATE U1674 ( .I1(n1637), .I2(n1583), .O(n1586) );
  NAND_GATE U1675 ( .I1(n1688), .I2(n1584), .O(n1585) );
  NAND_GATE U1676 ( .I1(n1586), .I2(n1585), .O(n1591) );
  NAND_GATE U1677 ( .I1(res_add[1]), .I2(n1691), .O(n1590) );
  NAND_GATE U1678 ( .I1(n696), .I2(n13), .O(n1588) );
  NAND3_GATE U1679 ( .I1(op1[1]), .I2(op2[1]), .I3(n75), .O(n1587) );
  AND_GATE U1680 ( .I1(n1588), .I2(n1587), .O(n1589) );
  AND3_GATE U1681 ( .I1(n1591), .I2(n1590), .I3(n1589), .O(n923) );
  NAND_GATE U1682 ( .I1(n80), .I2(n74), .O(n1592) );
  NAND_GATE U1683 ( .I1(n1619), .I2(n1592), .O(n525) );
  NAND_GATE U1684 ( .I1(n112), .I2(n74), .O(n1593) );
  NAND_GATE U1685 ( .I1(n1696), .I2(n1593), .O(n523) );
  NAND_GATE U1686 ( .I1(n399), .I2(n84), .O(n1597) );
  NAND_GATE U1687 ( .I1(n398), .I2(n85), .O(n1596) );
  NAND_GATE U1688 ( .I1(n397), .I2(n86), .O(n1595) );
  NAND_GATE U1689 ( .I1(n396), .I2(n87), .O(n1594) );
  NAND4_GATE U1690 ( .I1(n1597), .I2(n1596), .I3(n1595), .I4(n1594), .O(n1598)
         );
  INV_GATE U1691 ( .I1(n1598), .O(n2025) );
  NAND_GATE U1692 ( .I1(n167), .I2(n1598), .O(n1608) );
  NAND_GATE U1693 ( .I1(n2046), .I2(n1599), .O(n1601) );
  NAND_GATE U1694 ( .I1(n2047), .I2(n278), .O(n1600) );
  AND_GATE U1695 ( .I1(n1601), .I2(n1600), .O(n1607) );
  NAND_GATE U1696 ( .I1(n374), .I2(n80), .O(n1605) );
  NAND_GATE U1697 ( .I1(n375), .I2(n81), .O(n1604) );
  NAND_GATE U1698 ( .I1(n377), .I2(n82), .O(n1603) );
  NAND_GATE U1699 ( .I1(n376), .I2(n83), .O(n1602) );
  AND4_GATE U1700 ( .I1(n1605), .I2(n1604), .I3(n1603), .I4(n1602), .O(n1606)
         );
  NAND5_GATE U1701 ( .I1(n497), .I2(n1635), .I3(n1608), .I4(n1607), .I5(n1606), 
        .O(n496) );
  NAND_GATE U1702 ( .I1(hilo[34]), .I2(n1700), .O(n482) );
  NAND_GATE U1703 ( .I1(n112), .I2(n80), .O(n1610) );
  INV_GATE U1704 ( .I1(n1610), .O(n1609) );
  NAND_GATE U1705 ( .I1(n1637), .I2(n1609), .O(n1612) );
  NAND_GATE U1706 ( .I1(n1688), .I2(n1610), .O(n1611) );
  NAND_GATE U1707 ( .I1(n1612), .I2(n1611), .O(n1617) );
  NAND_GATE U1708 ( .I1(res_add[2]), .I2(n1691), .O(n1616) );
  NAND_GATE U1709 ( .I1(n493), .I2(n13), .O(n1614) );
  NAND3_GATE U1710 ( .I1(op1[2]), .I2(op2[2]), .I3(n75), .O(n1613) );
  AND_GATE U1711 ( .I1(n1614), .I2(n1613), .O(n1615) );
  AND3_GATE U1712 ( .I1(n1617), .I2(n1616), .I3(n1615), .O(n485) );
  NAND_GATE U1713 ( .I1(n81), .I2(n74), .O(n1618) );
  NAND_GATE U1714 ( .I1(n1619), .I2(n1618), .O(n403) );
  NAND_GATE U1715 ( .I1(n113), .I2(n74), .O(n1620) );
  NAND_GATE U1716 ( .I1(n1696), .I2(n1620), .O(n401) );
  NAND_GATE U1717 ( .I1(n399), .I2(n85), .O(n1624) );
  NAND_GATE U1718 ( .I1(n398), .I2(n86), .O(n1623) );
  NAND_GATE U1719 ( .I1(n397), .I2(n87), .O(n1622) );
  NAND_GATE U1720 ( .I1(n396), .I2(n88), .O(n1621) );
  NAND4_GATE U1721 ( .I1(n1624), .I2(n1623), .I3(n1622), .I4(n1621), .O(n1625)
         );
  INV_GATE U1722 ( .I1(n1625), .O(n2024) );
  NAND_GATE U1723 ( .I1(n167), .I2(n1625), .O(n1634) );
  NAND_GATE U1724 ( .I1(n2046), .I2(n391), .O(n1627) );
  NAND_GATE U1725 ( .I1(n2047), .I2(n245), .O(n1626) );
  AND_GATE U1726 ( .I1(n1627), .I2(n1626), .O(n1633) );
  NAND_GATE U1727 ( .I1(n374), .I2(n81), .O(n1631) );
  NAND_GATE U1728 ( .I1(n375), .I2(n82), .O(n1630) );
  NAND_GATE U1729 ( .I1(n377), .I2(n83), .O(n1629) );
  NAND_GATE U1730 ( .I1(n376), .I2(n84), .O(n1628) );
  AND4_GATE U1731 ( .I1(n1631), .I2(n1630), .I3(n1629), .I4(n1628), .O(n1632)
         );
  NAND5_GATE U1732 ( .I1(n365), .I2(n1635), .I3(n1634), .I4(n1633), .I5(n1632), 
        .O(n364) );
  NAND_GATE U1733 ( .I1(hilo[35]), .I2(n1700), .O(n349) );
  OR_GATE U1734 ( .I1(op2[3]), .I2(op1[3]), .O(n1638) );
  INV_GATE U1735 ( .I1(n1638), .O(n1636) );
  NAND_GATE U1736 ( .I1(n1637), .I2(n1636), .O(n1640) );
  NAND_GATE U1737 ( .I1(n1688), .I2(n1638), .O(n1639) );
  NAND_GATE U1738 ( .I1(n1640), .I2(n1639), .O(n1645) );
  NAND_GATE U1739 ( .I1(res_add[3]), .I2(n1691), .O(n1644) );
  NAND_GATE U1740 ( .I1(n361), .I2(n13), .O(n1642) );
  NAND3_GATE U1741 ( .I1(op1[3]), .I2(op2[3]), .I3(n75), .O(n1641) );
  AND_GATE U1742 ( .I1(n1642), .I2(n1641), .O(n1643) );
  AND3_GATE U1743 ( .I1(n1645), .I2(n1644), .I3(n1643), .O(n352) );
  NAND_GATE U1744 ( .I1(n114), .I2(n74), .O(n1646) );
  NAND_GATE U1745 ( .I1(n1696), .I2(n1646), .O(n346) );
  NAND_GATE U1746 ( .I1(op1[4]), .I2(n75), .O(n1647) );
  NAND_GATE U1747 ( .I1(n1688), .I2(n1647), .O(n344) );
  NAND_GATE U1748 ( .I1(op1[4]), .I2(n1689), .O(n317) );
  INV_GATE U1749 ( .I1(n1688), .O(n1690) );
  NAND_GATE U1750 ( .I1(op1[4]), .I2(n1690), .O(n1649) );
  NAND_GATE U1751 ( .I1(res_add[4]), .I2(n1691), .O(n1648) );
  AND_GATE U1752 ( .I1(n1649), .I2(n1648), .O(n320) );
  NAND_GATE U1753 ( .I1(n114), .I2(n1694), .O(n1651) );
  NAND_GATE U1754 ( .I1(op1[4]), .I2(n74), .O(n1650) );
  NAND_GATE U1755 ( .I1(n1651), .I2(n1650), .O(n1652) );
  NAND_GATE U1756 ( .I1(n82), .I2(n1652), .O(n1658) );
  NAND_GATE U1757 ( .I1(n52), .I2(n7), .O(n1657) );
  NAND_GATE U1758 ( .I1(hilo[4]), .I2(n178), .O(n1655) );
  NAND_GATE U1759 ( .I1(hilo[36]), .I2(n1700), .O(n1654) );
  NAND_GATE U1760 ( .I1(n331), .I2(n1701), .O(n1653) );
  AND3_GATE U1761 ( .I1(n1655), .I2(n1654), .I3(n1653), .O(n1656) );
  AND3_GATE U1762 ( .I1(n1658), .I2(n1657), .I3(n1656), .O(n321) );
  NAND_GATE U1763 ( .I1(op1[5]), .I2(n75), .O(n1659) );
  NAND_GATE U1764 ( .I1(n1688), .I2(n1659), .O(n314) );
  NAND_GATE U1765 ( .I1(op1[5]), .I2(n1689), .O(n288) );
  NAND_GATE U1766 ( .I1(op1[5]), .I2(n1690), .O(n1661) );
  NAND_GATE U1767 ( .I1(res_add[5]), .I2(n1691), .O(n1660) );
  AND_GATE U1768 ( .I1(n1661), .I2(n1660), .O(n290) );
  NAND_GATE U1769 ( .I1(n115), .I2(n1694), .O(n1662) );
  NAND_GATE U1770 ( .I1(n83), .I2(n1662), .O(n1664) );
  NAND_GATE U1771 ( .I1(op2[5]), .I2(n1696), .O(n1663) );
  NAND_GATE U1772 ( .I1(n1664), .I2(n1663), .O(n1672) );
  NAND_GATE U1773 ( .I1(hilo[5]), .I2(n178), .O(n1671) );
  NAND_GATE U1774 ( .I1(hilo[37]), .I2(n1700), .O(n1670) );
  NAND_GATE U1775 ( .I1(n302), .I2(n1701), .O(n1669) );
  NAND_GATE U1776 ( .I1(op1[5]), .I2(n83), .O(n1666) );
  NAND_GATE U1777 ( .I1(n115), .I2(op2[5]), .O(n1665) );
  NAND_GATE U1778 ( .I1(n1666), .I2(n1665), .O(n1667) );
  NAND_GATE U1779 ( .I1(n74), .I2(n1667), .O(n1668) );
  AND5_GATE U1780 ( .I1(n1672), .I2(n1671), .I3(n1670), .I4(n1669), .I5(n1668), 
        .O(n291) );
  NAND_GATE U1781 ( .I1(op1[6]), .I2(n75), .O(n1673) );
  NAND_GATE U1782 ( .I1(n1688), .I2(n1673), .O(n284) );
  NAND_GATE U1783 ( .I1(op1[6]), .I2(n1689), .O(n255) );
  NAND_GATE U1784 ( .I1(op1[6]), .I2(n1690), .O(n1675) );
  NAND_GATE U1785 ( .I1(res_add[6]), .I2(n1691), .O(n1674) );
  AND_GATE U1786 ( .I1(n1675), .I2(n1674), .O(n257) );
  NAND_GATE U1787 ( .I1(n116), .I2(n1694), .O(n1676) );
  NAND_GATE U1788 ( .I1(n84), .I2(n1676), .O(n1678) );
  NAND_GATE U1789 ( .I1(op2[6]), .I2(n1696), .O(n1677) );
  NAND_GATE U1790 ( .I1(n1678), .I2(n1677), .O(n1686) );
  NAND_GATE U1791 ( .I1(hilo[6]), .I2(n178), .O(n1685) );
  NAND_GATE U1792 ( .I1(hilo[38]), .I2(n1700), .O(n1684) );
  NAND_GATE U1793 ( .I1(n269), .I2(n1701), .O(n1683) );
  NAND_GATE U1794 ( .I1(op1[6]), .I2(n84), .O(n1680) );
  NAND_GATE U1795 ( .I1(n116), .I2(op2[6]), .O(n1679) );
  NAND_GATE U1796 ( .I1(n1680), .I2(n1679), .O(n1681) );
  NAND_GATE U1797 ( .I1(n74), .I2(n1681), .O(n1682) );
  AND5_GATE U1798 ( .I1(n1686), .I2(n1685), .I3(n1684), .I4(n1683), .I5(n1682), 
        .O(n258) );
  NAND_GATE U1799 ( .I1(op1[7]), .I2(n75), .O(n1687) );
  NAND_GATE U1800 ( .I1(n1688), .I2(n1687), .O(n251) );
  NAND_GATE U1801 ( .I1(op1[7]), .I2(n1689), .O(n223) );
  NAND_GATE U1802 ( .I1(op1[7]), .I2(n1690), .O(n1693) );
  NAND_GATE U1803 ( .I1(res_add[7]), .I2(n1691), .O(n1692) );
  AND_GATE U1804 ( .I1(n1693), .I2(n1692), .O(n225) );
  NAND_GATE U1805 ( .I1(n117), .I2(n1694), .O(n1695) );
  NAND_GATE U1806 ( .I1(n85), .I2(n1695), .O(n1699) );
  NAND_GATE U1807 ( .I1(op2[7]), .I2(n1696), .O(n1698) );
  NAND_GATE U1808 ( .I1(n1699), .I2(n1698), .O(n1709) );
  NAND_GATE U1809 ( .I1(hilo[7]), .I2(n178), .O(n1708) );
  NAND_GATE U1810 ( .I1(hilo[39]), .I2(n1700), .O(n1707) );
  NAND_GATE U1811 ( .I1(n237), .I2(n1701), .O(n1706) );
  NAND_GATE U1812 ( .I1(op1[7]), .I2(n85), .O(n1703) );
  NAND_GATE U1813 ( .I1(n117), .I2(op2[7]), .O(n1702) );
  NAND_GATE U1871 ( .I1(n1703), .I2(n1702), .O(n1704) );
  NAND_GATE U1873 ( .I1(n74), .I2(n1704), .O(n1705) );
  AND5_GATE U1875 ( .I1(n1709), .I2(n1708), .I3(n1707), .I4(n1706), .I5(n1705), 
        .O(n226) );
  NAND_GATE U1877 ( .I1(N787), .I2(n9), .O(n1713) );
  NAND_GATE U1878 ( .I1(op1[12]), .I2(n2037), .O(n1712) );
  NAND_GATE U1879 ( .I1(N722), .I2(n10), .O(n1711) );
  NAND_GATE U1880 ( .I1(hilo[12]), .I2(n1697), .O(n1710) );
  NAND4_GATE U1881 ( .I1(n1713), .I2(n1712), .I3(n1711), .I4(n1710), .O(n1977)
         );
  NAND_GATE U1882 ( .I1(N788), .I2(n9), .O(n1717) );
  NAND_GATE U1883 ( .I1(op1[13]), .I2(n2037), .O(n1716) );
  NAND_GATE U1884 ( .I1(N723), .I2(n10), .O(n1715) );
  NAND_GATE U1885 ( .I1(hilo[13]), .I2(n1697), .O(n1714) );
  NAND4_GATE U1886 ( .I1(n1717), .I2(n1716), .I3(n1715), .I4(n1714), .O(n1976)
         );
  NAND_GATE U1887 ( .I1(N789), .I2(n9), .O(n1721) );
  NAND_GATE U1888 ( .I1(op1[14]), .I2(n2037), .O(n1720) );
  NAND_GATE U1889 ( .I1(N724), .I2(n10), .O(n1719) );
  NAND_GATE U1890 ( .I1(hilo[14]), .I2(n1697), .O(n1718) );
  NAND4_GATE U1891 ( .I1(n1721), .I2(n1720), .I3(n1719), .I4(n1718), .O(n1975)
         );
  NAND_GATE U1892 ( .I1(N790), .I2(n9), .O(n1725) );
  NAND_GATE U1893 ( .I1(op1[15]), .I2(n2037), .O(n1724) );
  NAND_GATE U1894 ( .I1(N725), .I2(n10), .O(n1723) );
  NAND_GATE U1895 ( .I1(hilo[15]), .I2(n1697), .O(n1722) );
  NAND4_GATE U1896 ( .I1(n1725), .I2(n1724), .I3(n1723), .I4(n1722), .O(n1974)
         );
  NAND_GATE U1897 ( .I1(N791), .I2(n9), .O(n1729) );
  NAND_GATE U1898 ( .I1(op1[16]), .I2(n2037), .O(n1728) );
  NAND_GATE U1899 ( .I1(N726), .I2(n10), .O(n1727) );
  NAND_GATE U1900 ( .I1(hilo[16]), .I2(n1697), .O(n1726) );
  NAND4_GATE U1901 ( .I1(n1729), .I2(n1728), .I3(n1727), .I4(n1726), .O(n1973)
         );
  NAND_GATE U1902 ( .I1(N792), .I2(n9), .O(n1733) );
  NAND_GATE U1903 ( .I1(op1[17]), .I2(n2037), .O(n1732) );
  NAND_GATE U1904 ( .I1(N727), .I2(n10), .O(n1731) );
  NAND_GATE U1905 ( .I1(hilo[17]), .I2(n1697), .O(n1730) );
  NAND4_GATE U1906 ( .I1(n1733), .I2(n1732), .I3(n1731), .I4(n1730), .O(n1972)
         );
  NAND_GATE U1907 ( .I1(N793), .I2(n9), .O(n1737) );
  NAND_GATE U1908 ( .I1(op1[18]), .I2(n2037), .O(n1736) );
  NAND_GATE U1909 ( .I1(N728), .I2(n10), .O(n1735) );
  NAND_GATE U1910 ( .I1(hilo[18]), .I2(n1697), .O(n1734) );
  NAND4_GATE U1911 ( .I1(n1737), .I2(n1736), .I3(n1735), .I4(n1734), .O(n1971)
         );
  NAND_GATE U1912 ( .I1(N794), .I2(n9), .O(n1741) );
  NAND_GATE U1913 ( .I1(op1[19]), .I2(n2037), .O(n1740) );
  NAND_GATE U1914 ( .I1(N729), .I2(n10), .O(n1739) );
  NAND_GATE U1915 ( .I1(hilo[19]), .I2(n1697), .O(n1738) );
  NAND4_GATE U1916 ( .I1(n1741), .I2(n1740), .I3(n1739), .I4(n1738), .O(n1970)
         );
  NAND_GATE U1917 ( .I1(N795), .I2(n9), .O(n1745) );
  NAND_GATE U1918 ( .I1(op1[20]), .I2(n2037), .O(n1744) );
  NAND_GATE U1919 ( .I1(N730), .I2(n10), .O(n1743) );
  NAND_GATE U1920 ( .I1(hilo[20]), .I2(n1697), .O(n1742) );
  NAND4_GATE U1921 ( .I1(n1745), .I2(n1744), .I3(n1743), .I4(n1742), .O(n1969)
         );
  NAND_GATE U1922 ( .I1(N796), .I2(n9), .O(n1749) );
  NAND_GATE U1923 ( .I1(op1[21]), .I2(n2037), .O(n1748) );
  NAND_GATE U1924 ( .I1(N731), .I2(n10), .O(n1747) );
  NAND_GATE U1925 ( .I1(hilo[21]), .I2(n1697), .O(n1746) );
  NAND4_GATE U1926 ( .I1(n1749), .I2(n1748), .I3(n1747), .I4(n1746), .O(n1968)
         );
  NAND_GATE U1927 ( .I1(N797), .I2(n9), .O(n1753) );
  NAND_GATE U1928 ( .I1(op1[22]), .I2(n2037), .O(n1752) );
  NAND_GATE U1929 ( .I1(N732), .I2(n10), .O(n1751) );
  NAND_GATE U1930 ( .I1(hilo[22]), .I2(n1697), .O(n1750) );
  NAND4_GATE U1931 ( .I1(n1753), .I2(n1752), .I3(n1751), .I4(n1750), .O(n1967)
         );
  NAND_GATE U1932 ( .I1(op1[23]), .I2(n2037), .O(n1757) );
  NAND_GATE U1933 ( .I1(N798), .I2(n9), .O(n1756) );
  NAND_GATE U1934 ( .I1(hilo[23]), .I2(n1697), .O(n1755) );
  NAND_GATE U1935 ( .I1(N733), .I2(n10), .O(n1754) );
  NAND4_GATE U1936 ( .I1(n1757), .I2(n1756), .I3(n1755), .I4(n1754), .O(n1966)
         );
  NAND_GATE U1937 ( .I1(N799), .I2(n9), .O(n1761) );
  NAND_GATE U1938 ( .I1(op1[24]), .I2(n2037), .O(n1760) );
  NAND_GATE U1939 ( .I1(N734), .I2(n10), .O(n1759) );
  NAND_GATE U1940 ( .I1(hilo[24]), .I2(n1697), .O(n1758) );
  NAND4_GATE U1941 ( .I1(n1761), .I2(n1760), .I3(n1759), .I4(n1758), .O(n1965)
         );
  NAND_GATE U1942 ( .I1(N800), .I2(n9), .O(n1765) );
  NAND_GATE U1943 ( .I1(op1[25]), .I2(n2037), .O(n1764) );
  NAND_GATE U1944 ( .I1(N735), .I2(n10), .O(n1763) );
  NAND_GATE U1945 ( .I1(hilo[25]), .I2(n1697), .O(n1762) );
  NAND4_GATE U1946 ( .I1(n1765), .I2(n1764), .I3(n1763), .I4(n1762), .O(n1964)
         );
  NAND_GATE U1947 ( .I1(N801), .I2(n9), .O(n1769) );
  NAND_GATE U1948 ( .I1(op1[26]), .I2(n2037), .O(n1768) );
  NAND_GATE U1949 ( .I1(N736), .I2(n10), .O(n1767) );
  NAND_GATE U1950 ( .I1(hilo[26]), .I2(n1697), .O(n1766) );
  NAND4_GATE U1951 ( .I1(n1769), .I2(n1768), .I3(n1767), .I4(n1766), .O(n1963)
         );
  NAND_GATE U1952 ( .I1(hilo[27]), .I2(n1697), .O(n1773) );
  NAND_GATE U1953 ( .I1(N737), .I2(n10), .O(n1772) );
  NAND_GATE U1954 ( .I1(op1[27]), .I2(n2037), .O(n1771) );
  NAND_GATE U1955 ( .I1(N802), .I2(n9), .O(n1770) );
  NAND4_GATE U1956 ( .I1(n1773), .I2(n1772), .I3(n1771), .I4(n1770), .O(n1962)
         );
  NAND_GATE U1957 ( .I1(N803), .I2(n9), .O(n1825) );
  NAND_GATE U1958 ( .I1(op1[28]), .I2(n2037), .O(n1824) );
  NAND_GATE U1959 ( .I1(N738), .I2(n10), .O(n1823) );
  NAND_GATE U1960 ( .I1(hilo[28]), .I2(n1697), .O(n1822) );
  NAND4_GATE U1961 ( .I1(n1825), .I2(n1824), .I3(n1823), .I4(n1822), .O(n1961)
         );
  NAND_GATE U1962 ( .I1(hilo[29]), .I2(n1697), .O(n1829) );
  NAND_GATE U1963 ( .I1(N739), .I2(n10), .O(n1828) );
  NAND_GATE U1964 ( .I1(op1[29]), .I2(n2037), .O(n1827) );
  NAND_GATE U1965 ( .I1(N804), .I2(n9), .O(n1826) );
  NAND4_GATE U1966 ( .I1(n1829), .I2(n1828), .I3(n1827), .I4(n1826), .O(n1960)
         );
  NAND_GATE U1967 ( .I1(hilo[30]), .I2(n1697), .O(n1833) );
  NAND_GATE U1968 ( .I1(N740), .I2(n10), .O(n1832) );
  NAND_GATE U1969 ( .I1(op1[30]), .I2(n2037), .O(n1831) );
  NAND_GATE U1970 ( .I1(N805), .I2(n9), .O(n1830) );
  NAND4_GATE U1971 ( .I1(n1833), .I2(n1832), .I3(n1831), .I4(n1830), .O(n1959)
         );
  NAND_GATE U1972 ( .I1(hilo[31]), .I2(n1697), .O(n1837) );
  NAND_GATE U1973 ( .I1(N741), .I2(n10), .O(n1836) );
  NAND_GATE U1974 ( .I1(op1[31]), .I2(n2037), .O(n1835) );
  NAND_GATE U1975 ( .I1(N806), .I2(n9), .O(n1834) );
  NAND4_GATE U1976 ( .I1(n1837), .I2(n1836), .I3(n1835), .I4(n1834), .O(n1958)
         );
  NAND_GATE U1977 ( .I1(N807), .I2(n9), .O(n1844) );
  NAND_GATE U1978 ( .I1(n1839), .I2(n1838), .O(n2020) );
  NAND_GATE U1979 ( .I1(hilo[32]), .I2(n2020), .O(n1843) );
  INV_GATE U1980 ( .I1(n1840), .O(n2021) );
  NAND_GATE U1981 ( .I1(op1[0]), .I2(n2021), .O(n1842) );
  NAND_GATE U1982 ( .I1(N742), .I2(n10), .O(n1841) );
  NAND4_GATE U1983 ( .I1(n1844), .I2(n1843), .I3(n1842), .I4(n1841), .O(n1957)
         );
  NAND_GATE U1984 ( .I1(N808), .I2(n9), .O(n1848) );
  NAND_GATE U1985 ( .I1(hilo[33]), .I2(n2020), .O(n1847) );
  NAND_GATE U1986 ( .I1(op1[1]), .I2(n2021), .O(n1846) );
  NAND_GATE U1987 ( .I1(N743), .I2(n10), .O(n1845) );
  NAND4_GATE U1988 ( .I1(n1848), .I2(n1847), .I3(n1846), .I4(n1845), .O(n1956)
         );
  NAND_GATE U1989 ( .I1(N809), .I2(n9), .O(n1852) );
  NAND_GATE U1990 ( .I1(hilo[34]), .I2(n2020), .O(n1851) );
  NAND_GATE U1991 ( .I1(op1[2]), .I2(n2021), .O(n1850) );
  NAND_GATE U1992 ( .I1(N744), .I2(n10), .O(n1849) );
  NAND4_GATE U1993 ( .I1(n1852), .I2(n1851), .I3(n1850), .I4(n1849), .O(n1955)
         );
  NAND_GATE U1994 ( .I1(N810), .I2(n9), .O(n1856) );
  NAND_GATE U1995 ( .I1(hilo[35]), .I2(n2020), .O(n1855) );
  NAND_GATE U1996 ( .I1(op1[3]), .I2(n2021), .O(n1854) );
  NAND_GATE U1997 ( .I1(N745), .I2(n10), .O(n1853) );
  NAND4_GATE U1998 ( .I1(n1856), .I2(n1855), .I3(n1854), .I4(n1853), .O(n1954)
         );
  NAND_GATE U1999 ( .I1(N811), .I2(n9), .O(n1860) );
  NAND_GATE U2000 ( .I1(hilo[36]), .I2(n2020), .O(n1859) );
  NAND_GATE U2004 ( .I1(op1[4]), .I2(n2021), .O(n1858) );
  NAND_GATE U2005 ( .I1(N746), .I2(n10), .O(n1857) );
  NAND4_GATE U2006 ( .I1(n1860), .I2(n1859), .I3(n1858), .I4(n1857), .O(n1953)
         );
  NAND_GATE U2007 ( .I1(hilo[37]), .I2(n2020), .O(n1864) );
  NAND_GATE U2008 ( .I1(op1[5]), .I2(n2021), .O(n1863) );
  NAND_GATE U2009 ( .I1(N812), .I2(n9), .O(n1862) );
  NAND_GATE U2010 ( .I1(N747), .I2(n10), .O(n1861) );
  NAND4_GATE U2011 ( .I1(n1864), .I2(n1863), .I3(n1862), .I4(n1861), .O(n1952)
         );
  NAND_GATE U2012 ( .I1(N813), .I2(n9), .O(n1868) );
  NAND_GATE U2013 ( .I1(hilo[38]), .I2(n2020), .O(n1867) );
  NAND_GATE U2014 ( .I1(op1[6]), .I2(n2021), .O(n1866) );
  NAND_GATE U2015 ( .I1(N748), .I2(n10), .O(n1865) );
  NAND4_GATE U2016 ( .I1(n1868), .I2(n1867), .I3(n1866), .I4(n1865), .O(n1951)
         );
  NAND_GATE U2017 ( .I1(N814), .I2(n9), .O(n1872) );
  NAND_GATE U2018 ( .I1(hilo[39]), .I2(n2020), .O(n1871) );
  NAND_GATE U2019 ( .I1(op1[7]), .I2(n2021), .O(n1870) );
  NAND_GATE U2020 ( .I1(N749), .I2(n10), .O(n1869) );
  NAND4_GATE U2021 ( .I1(n1872), .I2(n1871), .I3(n1870), .I4(n1869), .O(n1950)
         );
  NAND_GATE U2022 ( .I1(N815), .I2(n9), .O(n1876) );
  NAND_GATE U2023 ( .I1(N750), .I2(n10), .O(n1875) );
  NAND_GATE U2024 ( .I1(hilo[40]), .I2(n2020), .O(n1874) );
  NAND_GATE U2025 ( .I1(op1[8]), .I2(n2021), .O(n1873) );
  NAND4_GATE U2026 ( .I1(n1876), .I2(n1875), .I3(n1874), .I4(n1873), .O(n1949)
         );
  NAND_GATE U2027 ( .I1(hilo[41]), .I2(n2020), .O(n1878) );
  NAND_GATE U2028 ( .I1(op1[9]), .I2(n2021), .O(n1877) );
  NAND_GATE U2029 ( .I1(N817), .I2(n9), .O(n1882) );
  NAND_GATE U2030 ( .I1(hilo[42]), .I2(n2020), .O(n1881) );
  NAND_GATE U2031 ( .I1(op1[10]), .I2(n2021), .O(n1880) );
  NAND_GATE U2032 ( .I1(N752), .I2(n10), .O(n1879) );
  NAND4_GATE U2033 ( .I1(n1882), .I2(n1881), .I3(n1880), .I4(n1879), .O(n1947)
         );
  NAND_GATE U2034 ( .I1(N818), .I2(n9), .O(n1886) );
  NAND_GATE U2035 ( .I1(hilo[43]), .I2(n2020), .O(n1885) );
  NAND_GATE U2036 ( .I1(op1[11]), .I2(n2021), .O(n1884) );
  NAND_GATE U2037 ( .I1(N753), .I2(n10), .O(n1883) );
  NAND4_GATE U2038 ( .I1(n1886), .I2(n1885), .I3(n1884), .I4(n1883), .O(n1946)
         );
  NAND_GATE U2039 ( .I1(hilo[44]), .I2(n2020), .O(n1890) );
  NAND_GATE U2040 ( .I1(op1[12]), .I2(n2021), .O(n1889) );
  NAND_GATE U2041 ( .I1(N819), .I2(n9), .O(n1888) );
  NAND_GATE U2045 ( .I1(N754), .I2(n10), .O(n1887) );
  NAND4_GATE U2046 ( .I1(n1890), .I2(n1889), .I3(n1888), .I4(n1887), .O(n1945)
         );
  NAND_GATE U2047 ( .I1(op1[13]), .I2(n2021), .O(n1892) );
  NAND_GATE U2048 ( .I1(hilo[45]), .I2(n2020), .O(n1891) );
  NAND_GATE U2049 ( .I1(N821), .I2(n9), .O(n1896) );
  NAND_GATE U2050 ( .I1(hilo[46]), .I2(n2020), .O(n1895) );
  NAND_GATE U2051 ( .I1(op1[14]), .I2(n2021), .O(n1894) );
  NAND_GATE U2052 ( .I1(N756), .I2(n10), .O(n1893) );
  NAND4_GATE U2053 ( .I1(n1896), .I2(n1895), .I3(n1894), .I4(n1893), .O(n1943)
         );
  NAND_GATE U2054 ( .I1(hilo[47]), .I2(n2020), .O(n1900) );
  NAND_GATE U2055 ( .I1(op1[15]), .I2(n2021), .O(n1899) );
  NAND_GATE U2056 ( .I1(N822), .I2(n9), .O(n1898) );
  NAND_GATE U2057 ( .I1(N757), .I2(n10), .O(n1897) );
  NAND4_GATE U2058 ( .I1(n1900), .I2(n1899), .I3(n1898), .I4(n1897), .O(n1942)
         );
  NAND_GATE U2059 ( .I1(hilo[48]), .I2(n2020), .O(n1902) );
  NAND_GATE U2060 ( .I1(op1[16]), .I2(n2021), .O(n1901) );
  NAND_GATE U2061 ( .I1(op1[17]), .I2(n2021), .O(n1906) );
  NAND_GATE U2062 ( .I1(hilo[49]), .I2(n2020), .O(n1905) );
  NAND_GATE U2063 ( .I1(N824), .I2(n9), .O(n1904) );
  NAND_GATE U2064 ( .I1(N759), .I2(n10), .O(n1903) );
  NAND4_GATE U2065 ( .I1(n1906), .I2(n1905), .I3(n1904), .I4(n1903), .O(n1940)
         );
  NAND_GATE U2066 ( .I1(N825), .I2(n9), .O(n1913) );
  NAND_GATE U2067 ( .I1(N760), .I2(n10), .O(n1912) );
  NAND_GATE U2068 ( .I1(hilo[50]), .I2(n2020), .O(n1908) );
  NAND_GATE U2069 ( .I1(op1[18]), .I2(n2021), .O(n1907) );
  NAND4_GATE U2070 ( .I1(n1913), .I2(n1912), .I3(n1908), .I4(n1907), .O(n1939)
         );
  NAND_GATE U2071 ( .I1(hilo[51]), .I2(n2020), .O(n1917) );
  NAND_GATE U2072 ( .I1(op1[19]), .I2(n2021), .O(n1916) );
  NAND_GATE U2073 ( .I1(N826), .I2(n9), .O(n1915) );
  NAND_GATE U2074 ( .I1(N761), .I2(n10), .O(n1914) );
  NAND4_GATE U2075 ( .I1(n1917), .I2(n1916), .I3(n1915), .I4(n1914), .O(n1938)
         );
  NAND_GATE U2076 ( .I1(hilo[52]), .I2(n2020), .O(n1921) );
  NAND_GATE U2077 ( .I1(op1[20]), .I2(n2021), .O(n1920) );
  NAND_GATE U2078 ( .I1(N827), .I2(n9), .O(n1919) );
  NAND_GATE U2079 ( .I1(N762), .I2(n10), .O(n1918) );
  NAND4_GATE U2080 ( .I1(n1921), .I2(n1920), .I3(n1919), .I4(n1918), .O(n1937)
         );
  NAND_GATE U2081 ( .I1(hilo[53]), .I2(n2020), .O(n1991) );
  NAND_GATE U2082 ( .I1(op1[21]), .I2(n2021), .O(n1990) );
  NAND_GATE U2083 ( .I1(N828), .I2(n9), .O(n1925) );
  NAND_GATE U2084 ( .I1(N763), .I2(n10), .O(n1924) );
  NAND4_GATE U2085 ( .I1(n1991), .I2(n1990), .I3(n1925), .I4(n1924), .O(n1936)
         );
  NAND_GATE U2086 ( .I1(hilo[54]), .I2(n2020), .O(n1995) );
  NAND_GATE U2087 ( .I1(op1[22]), .I2(n2021), .O(n1994) );
  NAND_GATE U2088 ( .I1(N829), .I2(n9), .O(n1993) );
  NAND_GATE U2089 ( .I1(N764), .I2(n10), .O(n1992) );
  NAND4_GATE U2090 ( .I1(n1995), .I2(n1994), .I3(n1993), .I4(n1992), .O(n1935)
         );
  NAND_GATE U2091 ( .I1(hilo[55]), .I2(n2020), .O(n1999) );
  NAND_GATE U2092 ( .I1(op1[23]), .I2(n2021), .O(n1998) );
  NAND_GATE U2093 ( .I1(N830), .I2(n9), .O(n1997) );
  NAND_GATE U2094 ( .I1(N765), .I2(n10), .O(n1996) );
  NAND4_GATE U2095 ( .I1(n1999), .I2(n1998), .I3(n1997), .I4(n1996), .O(n1934)
         );
  NAND_GATE U2096 ( .I1(hilo[56]), .I2(n2020), .O(n2001) );
  NAND_GATE U2097 ( .I1(op1[24]), .I2(n2021), .O(n2000) );
  NAND_GATE U2098 ( .I1(hilo[57]), .I2(n2020), .O(n2005) );
  NAND_GATE U2099 ( .I1(op1[25]), .I2(n2021), .O(n2004) );
  NAND_GATE U2100 ( .I1(N832), .I2(n9), .O(n2003) );
  NAND_GATE U2101 ( .I1(N767), .I2(n10), .O(n2002) );
  NAND4_GATE U2102 ( .I1(n2005), .I2(n2004), .I3(n2003), .I4(n2002), .O(n1932)
         );
  NAND_GATE U2103 ( .I1(hilo[58]), .I2(n2020), .O(n2009) );
  NAND_GATE U2104 ( .I1(op1[26]), .I2(n2021), .O(n2008) );
  NAND_GATE U2105 ( .I1(N833), .I2(n9), .O(n2007) );
  NAND_GATE U2106 ( .I1(N768), .I2(n10), .O(n2006) );
  NAND4_GATE U2107 ( .I1(n2009), .I2(n2008), .I3(n2007), .I4(n2006), .O(n1931)
         );
  NAND_GATE U2108 ( .I1(hilo[59]), .I2(n2020), .O(n2013) );
  NAND_GATE U2109 ( .I1(op1[27]), .I2(n2021), .O(n2012) );
  NAND_GATE U2110 ( .I1(N834), .I2(n9), .O(n2011) );
  NAND_GATE U2111 ( .I1(N769), .I2(n10), .O(n2010) );
  NAND4_GATE U2112 ( .I1(n2013), .I2(n2012), .I3(n2011), .I4(n2010), .O(n1930)
         );
  NAND_GATE U2113 ( .I1(hilo[60]), .I2(n2020), .O(n2015) );
  NAND_GATE U2114 ( .I1(op1[28]), .I2(n2021), .O(n2014) );
  NAND_GATE U2115 ( .I1(hilo[61]), .I2(n2020), .O(n2017) );
  NAND_GATE U2116 ( .I1(op1[29]), .I2(n2021), .O(n2016) );
  NAND_GATE U2117 ( .I1(hilo[62]), .I2(n2020), .O(n2019) );
  NAND_GATE U2118 ( .I1(op1[30]), .I2(n2021), .O(n2018) );
  NAND_GATE U2119 ( .I1(hilo[63]), .I2(n2020), .O(n2023) );
  NAND_GATE U2120 ( .I1(op1[31]), .I2(n2021), .O(n2022) );
  INV_GATE U2121 ( .I1(n759), .O(n2052) );
  INV_GATE U2122 ( .I1(n843), .O(n2053) );
  INV_GATE U2123 ( .I1(n844), .O(n2054) );
  INV_GATE U2124 ( .I1(n802), .O(n2055) );
  INV_GATE U2125 ( .I1(n801), .O(n2056) );
  INV_GATE U2126 ( .I1(n717), .O(n2057) );
endmodule


module predict_nb_record3_1 ( clock, reset, PF_pc, DI_bra, DI_adr, 
        EX_bra_confirm, EX_adr, EX_adresse, EX_uncleared, PR_bra_cmd, 
        PR_bra_bad, PR_bra_adr, PR_clear );
  input [31:0] PF_pc;
  input [31:0] DI_adr;
  input [31:0] EX_adr;
  input [31:0] EX_adresse;
  output [31:0] PR_bra_adr;
  input clock, reset, DI_bra, EX_bra_confirm, EX_uncleared;
  output PR_bra_cmd, PR_bra_bad, PR_clear;
  wire   \pre_pred_tab[1][IS_AFFECTED] , \pre_pred_tab[2][IS_AFFECTED] ,
         \pre_pred_tab[3][IS_AFFECTED] , \pred_tab[1][IS_AFFECTED] ,
         \pred_tab[1][LAST_BRA] , \pred_tab[1][CODE_ADR][31] ,
         \pred_tab[1][CODE_ADR][30] , \pred_tab[1][CODE_ADR][29] ,
         \pred_tab[1][CODE_ADR][28] , \pred_tab[1][CODE_ADR][27] ,
         \pred_tab[1][CODE_ADR][26] , \pred_tab[1][CODE_ADR][25] ,
         \pred_tab[1][CODE_ADR][24] , \pred_tab[1][CODE_ADR][23] ,
         \pred_tab[1][CODE_ADR][22] , \pred_tab[1][CODE_ADR][21] ,
         \pred_tab[1][CODE_ADR][20] , \pred_tab[1][CODE_ADR][19] ,
         \pred_tab[1][CODE_ADR][18] , \pred_tab[1][CODE_ADR][17] ,
         \pred_tab[1][CODE_ADR][16] , \pred_tab[1][CODE_ADR][15] ,
         \pred_tab[1][CODE_ADR][14] , \pred_tab[1][CODE_ADR][13] ,
         \pred_tab[1][CODE_ADR][12] , \pred_tab[1][CODE_ADR][11] ,
         \pred_tab[1][CODE_ADR][10] , \pred_tab[1][CODE_ADR][9] ,
         \pred_tab[1][CODE_ADR][8] , \pred_tab[1][CODE_ADR][7] ,
         \pred_tab[1][CODE_ADR][6] , \pred_tab[1][CODE_ADR][5] ,
         \pred_tab[1][CODE_ADR][4] , \pred_tab[1][CODE_ADR][3] ,
         \pred_tab[1][CODE_ADR][2] , \pred_tab[1][CODE_ADR][1] ,
         \pred_tab[1][CODE_ADR][0] , \pred_tab[1][BRA_ADR][31] ,
         \pred_tab[1][BRA_ADR][30] , \pred_tab[1][BRA_ADR][29] ,
         \pred_tab[1][BRA_ADR][28] , \pred_tab[1][BRA_ADR][27] ,
         \pred_tab[1][BRA_ADR][26] , \pred_tab[1][BRA_ADR][25] ,
         \pred_tab[1][BRA_ADR][24] , \pred_tab[1][BRA_ADR][23] ,
         \pred_tab[1][BRA_ADR][22] , \pred_tab[1][BRA_ADR][21] ,
         \pred_tab[1][BRA_ADR][20] , \pred_tab[1][BRA_ADR][19] ,
         \pred_tab[1][BRA_ADR][18] , \pred_tab[1][BRA_ADR][17] ,
         \pred_tab[1][BRA_ADR][16] , \pred_tab[1][BRA_ADR][15] ,
         \pred_tab[1][BRA_ADR][14] , \pred_tab[1][BRA_ADR][13] ,
         \pred_tab[1][BRA_ADR][12] , \pred_tab[1][BRA_ADR][11] ,
         \pred_tab[1][BRA_ADR][10] , \pred_tab[1][BRA_ADR][9] ,
         \pred_tab[1][BRA_ADR][8] , \pred_tab[1][BRA_ADR][7] ,
         \pred_tab[1][BRA_ADR][6] , \pred_tab[1][BRA_ADR][5] ,
         \pred_tab[1][BRA_ADR][4] , \pred_tab[1][BRA_ADR][3] ,
         \pred_tab[1][BRA_ADR][2] , \pred_tab[1][BRA_ADR][1] ,
         \pred_tab[1][BRA_ADR][0] , \pred_tab[2][IS_AFFECTED] ,
         \pred_tab[2][LAST_BRA] , \pred_tab[2][CODE_ADR][31] ,
         \pred_tab[2][CODE_ADR][30] , \pred_tab[2][CODE_ADR][29] ,
         \pred_tab[2][CODE_ADR][28] , \pred_tab[2][CODE_ADR][27] ,
         \pred_tab[2][CODE_ADR][26] , \pred_tab[2][CODE_ADR][25] ,
         \pred_tab[2][CODE_ADR][24] , \pred_tab[2][CODE_ADR][23] ,
         \pred_tab[2][CODE_ADR][22] , \pred_tab[2][CODE_ADR][21] ,
         \pred_tab[2][CODE_ADR][20] , \pred_tab[2][CODE_ADR][19] ,
         \pred_tab[2][CODE_ADR][18] , \pred_tab[2][CODE_ADR][17] ,
         \pred_tab[2][CODE_ADR][16] , \pred_tab[2][CODE_ADR][15] ,
         \pred_tab[2][CODE_ADR][14] , \pred_tab[2][CODE_ADR][13] ,
         \pred_tab[2][CODE_ADR][12] , \pred_tab[2][CODE_ADR][11] ,
         \pred_tab[2][CODE_ADR][10] , \pred_tab[2][CODE_ADR][9] ,
         \pred_tab[2][CODE_ADR][8] , \pred_tab[2][CODE_ADR][7] ,
         \pred_tab[2][CODE_ADR][6] , \pred_tab[2][CODE_ADR][5] ,
         \pred_tab[2][CODE_ADR][4] , \pred_tab[2][CODE_ADR][3] ,
         \pred_tab[2][CODE_ADR][2] , \pred_tab[2][CODE_ADR][1] ,
         \pred_tab[2][CODE_ADR][0] , \pred_tab[2][BRA_ADR][31] ,
         \pred_tab[2][BRA_ADR][30] , \pred_tab[2][BRA_ADR][29] ,
         \pred_tab[2][BRA_ADR][28] , \pred_tab[2][BRA_ADR][27] ,
         \pred_tab[2][BRA_ADR][26] , \pred_tab[2][BRA_ADR][25] ,
         \pred_tab[2][BRA_ADR][24] , \pred_tab[2][BRA_ADR][23] ,
         \pred_tab[2][BRA_ADR][22] , \pred_tab[2][BRA_ADR][21] ,
         \pred_tab[2][BRA_ADR][20] , \pred_tab[2][BRA_ADR][19] ,
         \pred_tab[2][BRA_ADR][18] , \pred_tab[2][BRA_ADR][17] ,
         \pred_tab[2][BRA_ADR][16] , \pred_tab[2][BRA_ADR][15] ,
         \pred_tab[2][BRA_ADR][14] , \pred_tab[2][BRA_ADR][13] ,
         \pred_tab[2][BRA_ADR][12] , \pred_tab[2][BRA_ADR][11] ,
         \pred_tab[2][BRA_ADR][10] , \pred_tab[2][BRA_ADR][9] ,
         \pred_tab[2][BRA_ADR][8] , \pred_tab[2][BRA_ADR][7] ,
         \pred_tab[2][BRA_ADR][6] , \pred_tab[2][BRA_ADR][5] ,
         \pred_tab[2][BRA_ADR][4] , \pred_tab[2][BRA_ADR][3] ,
         \pred_tab[2][BRA_ADR][2] , \pred_tab[2][BRA_ADR][1] ,
         \pred_tab[2][BRA_ADR][0] , \pred_tab[3][IS_AFFECTED] ,
         \pred_tab[3][LAST_BRA] , \pred_tab[3][CODE_ADR][31] ,
         \pred_tab[3][CODE_ADR][30] , \pred_tab[3][CODE_ADR][29] ,
         \pred_tab[3][CODE_ADR][28] , \pred_tab[3][CODE_ADR][27] ,
         \pred_tab[3][CODE_ADR][26] , \pred_tab[3][CODE_ADR][25] ,
         \pred_tab[3][CODE_ADR][24] , \pred_tab[3][CODE_ADR][23] ,
         \pred_tab[3][CODE_ADR][22] , \pred_tab[3][CODE_ADR][21] ,
         \pred_tab[3][CODE_ADR][20] , \pred_tab[3][CODE_ADR][19] ,
         \pred_tab[3][CODE_ADR][18] , \pred_tab[3][CODE_ADR][17] ,
         \pred_tab[3][CODE_ADR][16] , \pred_tab[3][CODE_ADR][15] ,
         \pred_tab[3][CODE_ADR][14] , \pred_tab[3][CODE_ADR][13] ,
         \pred_tab[3][CODE_ADR][12] , \pred_tab[3][CODE_ADR][11] ,
         \pred_tab[3][CODE_ADR][10] , \pred_tab[3][CODE_ADR][9] ,
         \pred_tab[3][CODE_ADR][8] , \pred_tab[3][CODE_ADR][7] ,
         \pred_tab[3][CODE_ADR][6] , \pred_tab[3][CODE_ADR][5] ,
         \pred_tab[3][CODE_ADR][4] , \pred_tab[3][CODE_ADR][3] ,
         \pred_tab[3][CODE_ADR][2] , \pred_tab[3][CODE_ADR][1] ,
         \pred_tab[3][CODE_ADR][0] , \pred_tab[3][BRA_ADR][31] ,
         \pred_tab[3][BRA_ADR][30] , \pred_tab[3][BRA_ADR][29] ,
         \pred_tab[3][BRA_ADR][28] , \pred_tab[3][BRA_ADR][27] ,
         \pred_tab[3][BRA_ADR][26] , \pred_tab[3][BRA_ADR][25] ,
         \pred_tab[3][BRA_ADR][24] , \pred_tab[3][BRA_ADR][23] ,
         \pred_tab[3][BRA_ADR][22] , \pred_tab[3][BRA_ADR][21] ,
         \pred_tab[3][BRA_ADR][20] , \pred_tab[3][BRA_ADR][19] ,
         \pred_tab[3][BRA_ADR][18] , \pred_tab[3][BRA_ADR][17] ,
         \pred_tab[3][BRA_ADR][16] , \pred_tab[3][BRA_ADR][15] ,
         \pred_tab[3][BRA_ADR][14] , \pred_tab[3][BRA_ADR][13] ,
         \pred_tab[3][BRA_ADR][12] , \pred_tab[3][BRA_ADR][11] ,
         \pred_tab[3][BRA_ADR][10] , \pred_tab[3][BRA_ADR][9] ,
         \pred_tab[3][BRA_ADR][8] , \pred_tab[3][BRA_ADR][7] ,
         \pred_tab[3][BRA_ADR][6] , \pred_tab[3][BRA_ADR][5] ,
         \pred_tab[3][BRA_ADR][4] , \pred_tab[3][BRA_ADR][3] ,
         \pred_tab[3][BRA_ADR][2] , \pred_tab[3][BRA_ADR][1] ,
         \pred_tab[3][BRA_ADR][0] , N69, N70, N71, N76, N79, N82, N92, N96,
         N100, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589,
         N590, N591, N592, N593, N594, N595, N596, N597, N598, N599,
         \next_out[1] , \next_out[0] , N1244, N1245, N1246, N1247, N1248,
         N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258,
         N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268,
         N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1579, N1582, N1614,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n428, n429,
         n430, n431, n432, n433, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n643,
         n644, n645, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1221, n1222, n1224, n1225, n1226, n1228, n1230,
         n1231, n1232, n1234, n1235, n1236, n1237, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1640, n1641, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n427, n434,
         n447, n512, n577, n642, n646, PR_clear, n1223, n1227, n1229, n1233,
         n1238;
  assign PR_bra_cmd = N1579;
  assign PR_bra_bad = PR_clear;

  FLIP_FLOP_D_PRESET \next_out_reg[0]  ( .D(n1641), .CK(clock), .PRESET(n434), 
        .Q(\next_out[0] ) );
  FLIP_FLOP_D_RESET \pred_tab_reg[2][IS_AFFECTED]  ( .D(
        \pre_pred_tab[2][IS_AFFECTED] ), .CK(clock), .RESET(n434), .Q(
        \pred_tab[2][IS_AFFECTED] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][0]  ( .D(n1637), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][0] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][10]  ( .D(n1636), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][10] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][11]  ( .D(n1635), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][11] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][12]  ( .D(n1634), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][12] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][13]  ( .D(n1633), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][13] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][14]  ( .D(n1632), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][14] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][15]  ( .D(n1631), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][15] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][16]  ( .D(n1630), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][16] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][17]  ( .D(n1629), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][17] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][18]  ( .D(n1628), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][18] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][19]  ( .D(n1627), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][19] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][1]  ( .D(n1626), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][1] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][20]  ( .D(n1625), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][20] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][21]  ( .D(n1624), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][21] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][22]  ( .D(n1623), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][22] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][23]  ( .D(n1622), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][23] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][24]  ( .D(n1621), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][24] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][25]  ( .D(n1620), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][25] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][26]  ( .D(n1619), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][26] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][27]  ( .D(n1618), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][27] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][28]  ( .D(n1617), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][28] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][29]  ( .D(n1616), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][29] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][2]  ( .D(n1615), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][2] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][30]  ( .D(n1614), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][30] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][31]  ( .D(n1613), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][31] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][3]  ( .D(n1612), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][3] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][4]  ( .D(n1611), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][4] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][5]  ( .D(n1610), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][5] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][6]  ( .D(n1609), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][6] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][7]  ( .D(n1608), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][7] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][8]  ( .D(n1607), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][8] ) );
  FLIP_FLOP_D \pred_tab_reg[2][CODE_ADR][9]  ( .D(n1606), .CK(clock), .Q(
        \pred_tab[2][CODE_ADR][9] ) );
  FLIP_FLOP_D_RESET \next_out_reg[1]  ( .D(n1640), .CK(clock), .RESET(n434), 
        .Q(\next_out[1] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][0]  ( .D(n1605), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][0] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][10]  ( .D(n1604), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][10] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][11]  ( .D(n1603), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][11] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][12]  ( .D(n1602), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][12] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][13]  ( .D(n1601), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][13] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][14]  ( .D(n1600), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][14] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][15]  ( .D(n1599), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][15] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][16]  ( .D(n1598), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][16] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][17]  ( .D(n1597), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][17] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][18]  ( .D(n1596), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][18] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][19]  ( .D(n1595), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][19] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][1]  ( .D(n1594), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][1] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][20]  ( .D(n1593), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][20] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][21]  ( .D(n1592), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][21] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][22]  ( .D(n1591), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][22] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][23]  ( .D(n1590), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][23] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][24]  ( .D(n1589), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][24] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][25]  ( .D(n1588), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][25] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][26]  ( .D(n1587), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][26] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][27]  ( .D(n1586), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][27] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][28]  ( .D(n1585), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][28] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][29]  ( .D(n1584), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][29] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][2]  ( .D(n1583), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][2] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][30]  ( .D(n1582), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][30] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][31]  ( .D(n1581), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][31] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][3]  ( .D(n1580), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][3] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][4]  ( .D(n1579), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][4] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][5]  ( .D(n1578), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][5] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][6]  ( .D(n1577), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][6] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][7]  ( .D(n1576), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][7] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][8]  ( .D(n1575), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][8] ) );
  FLIP_FLOP_D \pred_tab_reg[3][CODE_ADR][9]  ( .D(n1574), .CK(clock), .Q(
        \pred_tab[3][CODE_ADR][9] ) );
  FLIP_FLOP_D_RESET \pred_tab_reg[3][IS_AFFECTED]  ( .D(
        \pre_pred_tab[3][IS_AFFECTED] ), .CK(clock), .RESET(n434), .Q(
        \pred_tab[3][IS_AFFECTED] ) );
  FLIP_FLOP_D_RESET \pred_tab_reg[1][IS_AFFECTED]  ( .D(
        \pre_pred_tab[1][IS_AFFECTED] ), .CK(clock), .RESET(n434), .Q(
        \pred_tab[1][IS_AFFECTED] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][0]  ( .D(n1573), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][0] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][10]  ( .D(n1572), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][10] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][11]  ( .D(n1571), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][11] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][12]  ( .D(n1570), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][12] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][13]  ( .D(n1569), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][13] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][14]  ( .D(n1568), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][14] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][15]  ( .D(n1567), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][15] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][16]  ( .D(n1566), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][16] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][17]  ( .D(n1565), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][17] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][18]  ( .D(n1564), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][18] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][19]  ( .D(n1563), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][19] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][1]  ( .D(n1562), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][1] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][20]  ( .D(n1561), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][20] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][21]  ( .D(n1560), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][21] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][22]  ( .D(n1559), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][22] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][23]  ( .D(n1558), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][23] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][24]  ( .D(n1557), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][24] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][25]  ( .D(n1556), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][25] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][26]  ( .D(n1555), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][26] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][27]  ( .D(n1554), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][27] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][28]  ( .D(n1553), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][28] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][29]  ( .D(n1552), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][29] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][2]  ( .D(n1551), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][2] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][30]  ( .D(n1550), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][30] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][31]  ( .D(n1549), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][31] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][3]  ( .D(n1548), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][3] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][4]  ( .D(n1547), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][4] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][5]  ( .D(n1546), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][5] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][6]  ( .D(n1545), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][6] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][7]  ( .D(n1544), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][7] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][8]  ( .D(n1543), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][8] ) );
  FLIP_FLOP_D \pred_tab_reg[1][CODE_ADR][9]  ( .D(n1542), .CK(clock), .Q(
        \pred_tab[1][CODE_ADR][9] ) );
  FLIP_FLOP_D \pred_tab_reg[3][LAST_BRA]  ( .D(n1541), .CK(clock), .Q(
        \pred_tab[3][LAST_BRA] ) );
  FLIP_FLOP_D \pred_tab_reg[1][LAST_BRA]  ( .D(n1540), .CK(clock), .Q(
        \pred_tab[1][LAST_BRA] ) );
  FLIP_FLOP_D \pred_tab_reg[2][LAST_BRA]  ( .D(n1539), .CK(clock), .Q(
        \pred_tab[2][LAST_BRA] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][0]  ( .D(n1538), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][0] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][9]  ( .D(n1537), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][9] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][8]  ( .D(n1536), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][8] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][7]  ( .D(n1535), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][7] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][6]  ( .D(n1534), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][6] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][5]  ( .D(n1533), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][5] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][4]  ( .D(n1532), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][4] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][3]  ( .D(n1531), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][3] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][31]  ( .D(n1530), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][31] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][30]  ( .D(n1529), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][30] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][2]  ( .D(n1528), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][2] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][29]  ( .D(n1527), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][29] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][28]  ( .D(n1526), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][28] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][27]  ( .D(n1525), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][27] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][26]  ( .D(n1524), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][26] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][25]  ( .D(n1523), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][25] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][24]  ( .D(n1522), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][24] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][23]  ( .D(n1521), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][23] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][22]  ( .D(n1520), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][22] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][21]  ( .D(n1519), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][21] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][20]  ( .D(n1518), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][20] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][1]  ( .D(n1517), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][1] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][19]  ( .D(n1516), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][19] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][18]  ( .D(n1515), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][18] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][17]  ( .D(n1514), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][17] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][16]  ( .D(n1513), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][16] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][15]  ( .D(n1512), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][15] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][14]  ( .D(n1511), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][14] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][13]  ( .D(n1510), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][13] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][12]  ( .D(n1509), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][12] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][11]  ( .D(n1508), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][11] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][10]  ( .D(n1507), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][10] ) );
  FLIP_FLOP_D \pred_tab_reg[3][BRA_ADR][0]  ( .D(n1506), .CK(clock), .Q(
        \pred_tab[3][BRA_ADR][0] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][9]  ( .D(n1505), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][9] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][8]  ( .D(n1504), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][8] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][7]  ( .D(n1503), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][7] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][6]  ( .D(n1502), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][6] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][5]  ( .D(n1501), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][5] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][4]  ( .D(n1500), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][4] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][3]  ( .D(n1499), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][3] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][31]  ( .D(n1498), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][31] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][30]  ( .D(n1497), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][30] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][2]  ( .D(n1496), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][2] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][29]  ( .D(n1495), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][29] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][28]  ( .D(n1494), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][28] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][27]  ( .D(n1493), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][27] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][26]  ( .D(n1492), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][26] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][25]  ( .D(n1491), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][25] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][24]  ( .D(n1490), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][24] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][23]  ( .D(n1489), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][23] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][22]  ( .D(n1488), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][22] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][21]  ( .D(n1487), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][21] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][20]  ( .D(n1486), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][20] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][1]  ( .D(n1485), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][1] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][19]  ( .D(n1484), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][19] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][18]  ( .D(n1483), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][18] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][17]  ( .D(n1482), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][17] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][16]  ( .D(n1481), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][16] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][15]  ( .D(n1480), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][15] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][14]  ( .D(n1479), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][14] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][13]  ( .D(n1478), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][13] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][12]  ( .D(n1477), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][12] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][11]  ( .D(n1476), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][11] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][10]  ( .D(n1475), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][10] ) );
  FLIP_FLOP_D \pred_tab_reg[2][BRA_ADR][0]  ( .D(n1474), .CK(clock), .Q(
        \pred_tab[2][BRA_ADR][0] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][9]  ( .D(n1473), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][9] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][8]  ( .D(n1472), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][8] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][7]  ( .D(n1471), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][7] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][6]  ( .D(n1470), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][6] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][5]  ( .D(n1469), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][5] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][4]  ( .D(n1468), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][4] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][3]  ( .D(n1467), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][3] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][31]  ( .D(n1466), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][31] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][30]  ( .D(n1465), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][30] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][2]  ( .D(n1464), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][2] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][29]  ( .D(n1463), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][29] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][28]  ( .D(n1462), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][28] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][27]  ( .D(n1461), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][27] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][26]  ( .D(n1460), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][26] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][25]  ( .D(n1459), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][25] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][24]  ( .D(n1458), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][24] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][23]  ( .D(n1457), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][23] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][22]  ( .D(n1456), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][22] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][21]  ( .D(n1455), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][21] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][20]  ( .D(n1454), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][20] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][1]  ( .D(n1453), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][1] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][19]  ( .D(n1452), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][19] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][18]  ( .D(n1451), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][18] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][17]  ( .D(n1450), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][17] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][16]  ( .D(n1449), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][16] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][15]  ( .D(n1448), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][15] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][14]  ( .D(n1447), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][14] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][13]  ( .D(n1446), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][13] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][12]  ( .D(n1445), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][12] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][11]  ( .D(n1444), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][11] ) );
  FLIP_FLOP_D \pred_tab_reg[1][BRA_ADR][10]  ( .D(n1443), .CK(clock), .Q(
        \pred_tab[1][BRA_ADR][10] ) );
  OR_GATE U3 ( .I1(\pred_tab[3][IS_AFFECTED] ), .I2(n642), .O(
        \pre_pred_tab[3][IS_AFFECTED] ) );
  OR_GATE U4 ( .I1(\pred_tab[2][IS_AFFECTED] ), .I2(n28), .O(
        \pre_pred_tab[2][IS_AFFECTED] ) );
  OR_GATE U5 ( .I1(\pred_tab[1][IS_AFFECTED] ), .I2(n29), .O(
        \pre_pred_tab[1][IS_AFFECTED] ) );
  NAND3_GATE U6 ( .I1(n30), .I2(n31), .I3(n32), .O(n1443) );
  NAND_GATE U7 ( .I1(\pred_tab[1][BRA_ADR][10] ), .I2(n33), .O(n32) );
  NAND_GATE U8 ( .I1(n34), .I2(n35), .O(n31) );
  NAND_GATE U9 ( .I1(N1254), .I2(n36), .O(n30) );
  NAND3_GATE U10 ( .I1(n37), .I2(n38), .I3(n39), .O(n1444) );
  NAND_GATE U11 ( .I1(\pred_tab[1][BRA_ADR][11] ), .I2(n33), .O(n39) );
  NAND_GATE U12 ( .I1(n34), .I2(n40), .O(n38) );
  NAND_GATE U13 ( .I1(N1255), .I2(n36), .O(n37) );
  NAND3_GATE U14 ( .I1(n41), .I2(n42), .I3(n43), .O(n1445) );
  NAND_GATE U15 ( .I1(\pred_tab[1][BRA_ADR][12] ), .I2(n33), .O(n43) );
  NAND_GATE U16 ( .I1(n34), .I2(n44), .O(n42) );
  NAND_GATE U29 ( .I1(N1256), .I2(n36), .O(n41) );
  NAND3_GATE U30 ( .I1(n45), .I2(n46), .I3(n47), .O(n1446) );
  NAND_GATE U31 ( .I1(\pred_tab[1][BRA_ADR][13] ), .I2(n33), .O(n47) );
  NAND_GATE U32 ( .I1(n34), .I2(n48), .O(n46) );
  NAND_GATE U33 ( .I1(N1257), .I2(n36), .O(n45) );
  NAND3_GATE U34 ( .I1(n49), .I2(n50), .I3(n51), .O(n1447) );
  NAND_GATE U35 ( .I1(\pred_tab[1][BRA_ADR][14] ), .I2(n33), .O(n51) );
  NAND_GATE U36 ( .I1(n34), .I2(n52), .O(n50) );
  NAND_GATE U37 ( .I1(N1258), .I2(n36), .O(n49) );
  NAND3_GATE U38 ( .I1(n53), .I2(n54), .I3(n55), .O(n1448) );
  NAND_GATE U39 ( .I1(\pred_tab[1][BRA_ADR][15] ), .I2(n33), .O(n55) );
  NAND_GATE U40 ( .I1(n34), .I2(n56), .O(n54) );
  NAND_GATE U41 ( .I1(N1259), .I2(n36), .O(n53) );
  NAND3_GATE U42 ( .I1(n57), .I2(n58), .I3(n59), .O(n1449) );
  NAND_GATE U43 ( .I1(\pred_tab[1][BRA_ADR][16] ), .I2(n33), .O(n59) );
  NAND_GATE U44 ( .I1(n34), .I2(n60), .O(n58) );
  NAND_GATE U45 ( .I1(N1260), .I2(n36), .O(n57) );
  NAND3_GATE U46 ( .I1(n61), .I2(n62), .I3(n63), .O(n1450) );
  NAND_GATE U47 ( .I1(\pred_tab[1][BRA_ADR][17] ), .I2(n33), .O(n63) );
  NAND_GATE U48 ( .I1(n34), .I2(n64), .O(n62) );
  NAND_GATE U49 ( .I1(N1261), .I2(n36), .O(n61) );
  NAND3_GATE U50 ( .I1(n65), .I2(n66), .I3(n67), .O(n1451) );
  NAND_GATE U51 ( .I1(\pred_tab[1][BRA_ADR][18] ), .I2(n33), .O(n67) );
  NAND_GATE U52 ( .I1(n34), .I2(n68), .O(n66) );
  NAND_GATE U53 ( .I1(N1262), .I2(n36), .O(n65) );
  NAND3_GATE U54 ( .I1(n69), .I2(n70), .I3(n71), .O(n1452) );
  NAND_GATE U55 ( .I1(\pred_tab[1][BRA_ADR][19] ), .I2(n33), .O(n71) );
  NAND_GATE U56 ( .I1(n34), .I2(n72), .O(n70) );
  NAND_GATE U57 ( .I1(N1263), .I2(n26), .O(n69) );
  NAND3_GATE U58 ( .I1(n73), .I2(n74), .I3(n75), .O(n1453) );
  NAND_GATE U59 ( .I1(\pred_tab[1][BRA_ADR][1] ), .I2(n33), .O(n75) );
  NAND_GATE U60 ( .I1(n34), .I2(n76), .O(n74) );
  NAND_GATE U61 ( .I1(N1245), .I2(n27), .O(n73) );
  NAND3_GATE U62 ( .I1(n77), .I2(n78), .I3(n79), .O(n1454) );
  NAND_GATE U63 ( .I1(\pred_tab[1][BRA_ADR][20] ), .I2(n33), .O(n79) );
  NAND_GATE U64 ( .I1(n34), .I2(n80), .O(n78) );
  NAND_GATE U65 ( .I1(N1264), .I2(n24), .O(n77) );
  NAND3_GATE U66 ( .I1(n81), .I2(n82), .I3(n83), .O(n1455) );
  NAND_GATE U67 ( .I1(\pred_tab[1][BRA_ADR][21] ), .I2(n33), .O(n83) );
  NAND_GATE U68 ( .I1(n34), .I2(n84), .O(n82) );
  NAND_GATE U69 ( .I1(N1265), .I2(n25), .O(n81) );
  NAND3_GATE U70 ( .I1(n85), .I2(n86), .I3(n87), .O(n1456) );
  NAND_GATE U71 ( .I1(\pred_tab[1][BRA_ADR][22] ), .I2(n33), .O(n87) );
  NAND_GATE U72 ( .I1(n34), .I2(n88), .O(n86) );
  NAND_GATE U73 ( .I1(N1266), .I2(n36), .O(n85) );
  NAND3_GATE U74 ( .I1(n89), .I2(n90), .I3(n91), .O(n1457) );
  NAND_GATE U75 ( .I1(\pred_tab[1][BRA_ADR][23] ), .I2(n33), .O(n91) );
  NAND_GATE U76 ( .I1(n34), .I2(n92), .O(n90) );
  NAND_GATE U77 ( .I1(N1267), .I2(n36), .O(n89) );
  NAND3_GATE U78 ( .I1(n93), .I2(n94), .I3(n95), .O(n1458) );
  NAND_GATE U79 ( .I1(\pred_tab[1][BRA_ADR][24] ), .I2(n33), .O(n95) );
  NAND_GATE U80 ( .I1(n34), .I2(n96), .O(n94) );
  NAND_GATE U81 ( .I1(N1268), .I2(n26), .O(n93) );
  NAND3_GATE U82 ( .I1(n97), .I2(n98), .I3(n99), .O(n1459) );
  NAND_GATE U83 ( .I1(\pred_tab[1][BRA_ADR][25] ), .I2(n33), .O(n99) );
  NAND_GATE U84 ( .I1(n34), .I2(n100), .O(n98) );
  NAND_GATE U85 ( .I1(N1269), .I2(n27), .O(n97) );
  NAND3_GATE U86 ( .I1(n101), .I2(n102), .I3(n103), .O(n1460) );
  NAND_GATE U87 ( .I1(\pred_tab[1][BRA_ADR][26] ), .I2(n33), .O(n103) );
  NAND_GATE U88 ( .I1(n34), .I2(n104), .O(n102) );
  NAND_GATE U89 ( .I1(N1270), .I2(n24), .O(n101) );
  NAND3_GATE U90 ( .I1(n105), .I2(n106), .I3(n107), .O(n1461) );
  NAND_GATE U91 ( .I1(\pred_tab[1][BRA_ADR][27] ), .I2(n33), .O(n107) );
  NAND_GATE U92 ( .I1(n34), .I2(n108), .O(n106) );
  NAND_GATE U93 ( .I1(N1271), .I2(n25), .O(n105) );
  NAND3_GATE U94 ( .I1(n109), .I2(n110), .I3(n111), .O(n1462) );
  NAND_GATE U95 ( .I1(\pred_tab[1][BRA_ADR][28] ), .I2(n33), .O(n111) );
  NAND_GATE U96 ( .I1(n34), .I2(n112), .O(n110) );
  NAND_GATE U97 ( .I1(N1272), .I2(n27), .O(n109) );
  NAND3_GATE U98 ( .I1(n113), .I2(n114), .I3(n115), .O(n1463) );
  NAND_GATE U99 ( .I1(\pred_tab[1][BRA_ADR][29] ), .I2(n33), .O(n115) );
  NAND_GATE U100 ( .I1(n34), .I2(n116), .O(n114) );
  NAND_GATE U101 ( .I1(N1273), .I2(n27), .O(n113) );
  NAND3_GATE U102 ( .I1(n117), .I2(n118), .I3(n119), .O(n1464) );
  NAND_GATE U103 ( .I1(\pred_tab[1][BRA_ADR][2] ), .I2(n33), .O(n119) );
  NAND_GATE U104 ( .I1(n34), .I2(n120), .O(n118) );
  NAND_GATE U105 ( .I1(N1246), .I2(n27), .O(n117) );
  NAND3_GATE U106 ( .I1(n121), .I2(n122), .I3(n123), .O(n1465) );
  NAND_GATE U107 ( .I1(\pred_tab[1][BRA_ADR][30] ), .I2(n33), .O(n123) );
  NAND_GATE U108 ( .I1(n34), .I2(n124), .O(n122) );
  NAND_GATE U109 ( .I1(N1274), .I2(n27), .O(n121) );
  NAND3_GATE U110 ( .I1(n125), .I2(n126), .I3(n127), .O(n1466) );
  NAND_GATE U111 ( .I1(\pred_tab[1][BRA_ADR][31] ), .I2(n33), .O(n127) );
  NAND_GATE U112 ( .I1(n34), .I2(n128), .O(n126) );
  NAND_GATE U113 ( .I1(N1275), .I2(n27), .O(n125) );
  NAND3_GATE U114 ( .I1(n129), .I2(n130), .I3(n131), .O(n1467) );
  NAND_GATE U115 ( .I1(\pred_tab[1][BRA_ADR][3] ), .I2(n33), .O(n131) );
  NAND_GATE U116 ( .I1(n34), .I2(n132), .O(n130) );
  NAND_GATE U117 ( .I1(N1247), .I2(n27), .O(n129) );
  NAND3_GATE U118 ( .I1(n133), .I2(n134), .I3(n135), .O(n1468) );
  NAND_GATE U119 ( .I1(\pred_tab[1][BRA_ADR][4] ), .I2(n33), .O(n135) );
  NAND_GATE U120 ( .I1(n34), .I2(n136), .O(n134) );
  NAND_GATE U121 ( .I1(N1248), .I2(n27), .O(n133) );
  NAND3_GATE U122 ( .I1(n137), .I2(n138), .I3(n139), .O(n1469) );
  NAND_GATE U123 ( .I1(\pred_tab[1][BRA_ADR][5] ), .I2(n33), .O(n139) );
  NAND_GATE U124 ( .I1(n34), .I2(n140), .O(n138) );
  NAND_GATE U125 ( .I1(N1249), .I2(n27), .O(n137) );
  NAND3_GATE U126 ( .I1(n141), .I2(n142), .I3(n143), .O(n1470) );
  NAND_GATE U127 ( .I1(\pred_tab[1][BRA_ADR][6] ), .I2(n33), .O(n143) );
  NAND_GATE U128 ( .I1(n34), .I2(n144), .O(n142) );
  NAND_GATE U129 ( .I1(N1250), .I2(n27), .O(n141) );
  NAND3_GATE U130 ( .I1(n145), .I2(n146), .I3(n147), .O(n1471) );
  NAND_GATE U131 ( .I1(\pred_tab[1][BRA_ADR][7] ), .I2(n33), .O(n147) );
  NAND_GATE U132 ( .I1(n34), .I2(n148), .O(n146) );
  NAND_GATE U133 ( .I1(N1251), .I2(n26), .O(n145) );
  NAND3_GATE U134 ( .I1(n149), .I2(n150), .I3(n151), .O(n1472) );
  NAND_GATE U135 ( .I1(\pred_tab[1][BRA_ADR][8] ), .I2(n33), .O(n151) );
  NAND_GATE U136 ( .I1(n34), .I2(n152), .O(n150) );
  NAND_GATE U137 ( .I1(N1252), .I2(n26), .O(n149) );
  NAND3_GATE U138 ( .I1(n153), .I2(n154), .I3(n155), .O(n1473) );
  NAND_GATE U139 ( .I1(\pred_tab[1][BRA_ADR][9] ), .I2(n33), .O(n155) );
  NAND_GATE U140 ( .I1(n34), .I2(n156), .O(n154) );
  NAND_GATE U141 ( .I1(N1253), .I2(n26), .O(n153) );
  NAND3_GATE U142 ( .I1(n157), .I2(n158), .I3(n159), .O(n1474) );
  NAND_GATE U143 ( .I1(\pred_tab[2][BRA_ADR][0] ), .I2(n160), .O(n159) );
  NAND_GATE U144 ( .I1(n161), .I2(n162), .O(n158) );
  NAND_GATE U145 ( .I1(N1244), .I2(n163), .O(n157) );
  NAND3_GATE U146 ( .I1(n164), .I2(n165), .I3(n166), .O(n1475) );
  NAND_GATE U147 ( .I1(\pred_tab[2][BRA_ADR][10] ), .I2(n160), .O(n166) );
  NAND_GATE U148 ( .I1(n161), .I2(n167), .O(n165) );
  NAND_GATE U149 ( .I1(n163), .I2(N1254), .O(n164) );
  NAND3_GATE U150 ( .I1(n168), .I2(n169), .I3(n170), .O(n1476) );
  NAND_GATE U151 ( .I1(\pred_tab[2][BRA_ADR][11] ), .I2(n160), .O(n170) );
  NAND_GATE U152 ( .I1(n161), .I2(n171), .O(n169) );
  NAND_GATE U153 ( .I1(n163), .I2(N1255), .O(n168) );
  NAND3_GATE U154 ( .I1(n172), .I2(n173), .I3(n174), .O(n1477) );
  NAND_GATE U155 ( .I1(\pred_tab[2][BRA_ADR][12] ), .I2(n160), .O(n174) );
  NAND_GATE U156 ( .I1(n161), .I2(n175), .O(n173) );
  NAND_GATE U157 ( .I1(n163), .I2(N1256), .O(n172) );
  NAND3_GATE U158 ( .I1(n176), .I2(n177), .I3(n178), .O(n1478) );
  NAND_GATE U159 ( .I1(\pred_tab[2][BRA_ADR][13] ), .I2(n160), .O(n178) );
  NAND_GATE U160 ( .I1(n161), .I2(n179), .O(n177) );
  NAND_GATE U161 ( .I1(n163), .I2(N1257), .O(n176) );
  NAND3_GATE U162 ( .I1(n180), .I2(n181), .I3(n182), .O(n1479) );
  NAND_GATE U163 ( .I1(\pred_tab[2][BRA_ADR][14] ), .I2(n160), .O(n182) );
  NAND_GATE U164 ( .I1(n161), .I2(n183), .O(n181) );
  NAND_GATE U165 ( .I1(n163), .I2(N1258), .O(n180) );
  NAND3_GATE U166 ( .I1(n184), .I2(n185), .I3(n186), .O(n1480) );
  NAND_GATE U167 ( .I1(\pred_tab[2][BRA_ADR][15] ), .I2(n160), .O(n186) );
  NAND_GATE U168 ( .I1(n161), .I2(n187), .O(n185) );
  NAND_GATE U169 ( .I1(n163), .I2(N1259), .O(n184) );
  NAND3_GATE U170 ( .I1(n188), .I2(n189), .I3(n190), .O(n1481) );
  NAND_GATE U171 ( .I1(\pred_tab[2][BRA_ADR][16] ), .I2(n160), .O(n190) );
  NAND_GATE U172 ( .I1(n161), .I2(n191), .O(n189) );
  NAND_GATE U173 ( .I1(n163), .I2(N1260), .O(n188) );
  NAND3_GATE U174 ( .I1(n192), .I2(n193), .I3(n194), .O(n1482) );
  NAND_GATE U175 ( .I1(\pred_tab[2][BRA_ADR][17] ), .I2(n160), .O(n194) );
  NAND_GATE U176 ( .I1(n161), .I2(n195), .O(n193) );
  NAND_GATE U177 ( .I1(n163), .I2(N1261), .O(n192) );
  NAND3_GATE U178 ( .I1(n196), .I2(n197), .I3(n198), .O(n1483) );
  NAND_GATE U179 ( .I1(\pred_tab[2][BRA_ADR][18] ), .I2(n160), .O(n198) );
  NAND_GATE U180 ( .I1(n161), .I2(n199), .O(n197) );
  NAND_GATE U181 ( .I1(n21), .I2(N1262), .O(n196) );
  NAND3_GATE U182 ( .I1(n200), .I2(n201), .I3(n202), .O(n1484) );
  NAND_GATE U183 ( .I1(\pred_tab[2][BRA_ADR][19] ), .I2(n160), .O(n202) );
  NAND_GATE U184 ( .I1(n161), .I2(n203), .O(n201) );
  NAND_GATE U185 ( .I1(n22), .I2(N1263), .O(n200) );
  NAND3_GATE U186 ( .I1(n204), .I2(n205), .I3(n206), .O(n1485) );
  NAND_GATE U187 ( .I1(\pred_tab[2][BRA_ADR][1] ), .I2(n160), .O(n206) );
  NAND_GATE U188 ( .I1(n161), .I2(n207), .O(n205) );
  NAND_GATE U189 ( .I1(n19), .I2(N1245), .O(n204) );
  NAND3_GATE U190 ( .I1(n208), .I2(n209), .I3(n210), .O(n1486) );
  NAND_GATE U191 ( .I1(\pred_tab[2][BRA_ADR][20] ), .I2(n160), .O(n210) );
  NAND_GATE U192 ( .I1(n161), .I2(n211), .O(n209) );
  NAND_GATE U193 ( .I1(n20), .I2(N1264), .O(n208) );
  NAND3_GATE U194 ( .I1(n212), .I2(n213), .I3(n214), .O(n1487) );
  NAND_GATE U195 ( .I1(\pred_tab[2][BRA_ADR][21] ), .I2(n160), .O(n214) );
  NAND_GATE U196 ( .I1(n161), .I2(n215), .O(n213) );
  NAND_GATE U197 ( .I1(n163), .I2(N1265), .O(n212) );
  NAND3_GATE U198 ( .I1(n216), .I2(n217), .I3(n218), .O(n1488) );
  NAND_GATE U199 ( .I1(\pred_tab[2][BRA_ADR][22] ), .I2(n160), .O(n218) );
  NAND_GATE U200 ( .I1(n161), .I2(n219), .O(n217) );
  NAND_GATE U201 ( .I1(n163), .I2(N1266), .O(n216) );
  NAND3_GATE U202 ( .I1(n220), .I2(n221), .I3(n222), .O(n1489) );
  NAND_GATE U203 ( .I1(\pred_tab[2][BRA_ADR][23] ), .I2(n160), .O(n222) );
  NAND_GATE U204 ( .I1(n161), .I2(n223), .O(n221) );
  NAND_GATE U205 ( .I1(n21), .I2(N1267), .O(n220) );
  NAND3_GATE U206 ( .I1(n224), .I2(n225), .I3(n226), .O(n1490) );
  NAND_GATE U207 ( .I1(\pred_tab[2][BRA_ADR][24] ), .I2(n160), .O(n226) );
  NAND_GATE U208 ( .I1(n161), .I2(n227), .O(n225) );
  NAND_GATE U209 ( .I1(n22), .I2(N1268), .O(n224) );
  NAND3_GATE U210 ( .I1(n228), .I2(n229), .I3(n230), .O(n1491) );
  NAND_GATE U211 ( .I1(\pred_tab[2][BRA_ADR][25] ), .I2(n160), .O(n230) );
  NAND_GATE U212 ( .I1(n161), .I2(n231), .O(n229) );
  NAND_GATE U213 ( .I1(n19), .I2(N1269), .O(n228) );
  NAND3_GATE U214 ( .I1(n232), .I2(n233), .I3(n234), .O(n1492) );
  NAND_GATE U215 ( .I1(\pred_tab[2][BRA_ADR][26] ), .I2(n160), .O(n234) );
  NAND_GATE U216 ( .I1(n161), .I2(n235), .O(n233) );
  NAND_GATE U217 ( .I1(n20), .I2(N1270), .O(n232) );
  NAND3_GATE U218 ( .I1(n236), .I2(n237), .I3(n238), .O(n1493) );
  NAND_GATE U219 ( .I1(\pred_tab[2][BRA_ADR][27] ), .I2(n160), .O(n238) );
  NAND_GATE U220 ( .I1(n161), .I2(n239), .O(n237) );
  NAND_GATE U221 ( .I1(n22), .I2(N1271), .O(n236) );
  NAND3_GATE U222 ( .I1(n240), .I2(n241), .I3(n242), .O(n1494) );
  NAND_GATE U223 ( .I1(\pred_tab[2][BRA_ADR][28] ), .I2(n160), .O(n242) );
  NAND_GATE U224 ( .I1(n161), .I2(n243), .O(n241) );
  NAND_GATE U225 ( .I1(n22), .I2(N1272), .O(n240) );
  NAND3_GATE U226 ( .I1(n244), .I2(n245), .I3(n246), .O(n1495) );
  NAND_GATE U227 ( .I1(\pred_tab[2][BRA_ADR][29] ), .I2(n160), .O(n246) );
  NAND_GATE U228 ( .I1(n161), .I2(n247), .O(n245) );
  NAND_GATE U229 ( .I1(n22), .I2(N1273), .O(n244) );
  NAND3_GATE U230 ( .I1(n248), .I2(n249), .I3(n250), .O(n1496) );
  NAND_GATE U231 ( .I1(\pred_tab[2][BRA_ADR][2] ), .I2(n160), .O(n250) );
  NAND_GATE U232 ( .I1(n161), .I2(n251), .O(n249) );
  NAND_GATE U233 ( .I1(n22), .I2(N1246), .O(n248) );
  NAND3_GATE U234 ( .I1(n252), .I2(n253), .I3(n254), .O(n1497) );
  NAND_GATE U235 ( .I1(\pred_tab[2][BRA_ADR][30] ), .I2(n160), .O(n254) );
  NAND_GATE U236 ( .I1(n161), .I2(n255), .O(n253) );
  NAND_GATE U237 ( .I1(n22), .I2(N1274), .O(n252) );
  NAND3_GATE U238 ( .I1(n256), .I2(n257), .I3(n258), .O(n1498) );
  NAND_GATE U239 ( .I1(\pred_tab[2][BRA_ADR][31] ), .I2(n160), .O(n258) );
  NAND_GATE U240 ( .I1(n161), .I2(n259), .O(n257) );
  NAND_GATE U241 ( .I1(n22), .I2(N1275), .O(n256) );
  NAND3_GATE U242 ( .I1(n260), .I2(n261), .I3(n262), .O(n1499) );
  NAND_GATE U243 ( .I1(\pred_tab[2][BRA_ADR][3] ), .I2(n160), .O(n262) );
  NAND_GATE U244 ( .I1(n161), .I2(n263), .O(n261) );
  NAND_GATE U245 ( .I1(n22), .I2(N1247), .O(n260) );
  NAND3_GATE U246 ( .I1(n264), .I2(n265), .I3(n266), .O(n1500) );
  NAND_GATE U247 ( .I1(\pred_tab[2][BRA_ADR][4] ), .I2(n160), .O(n266) );
  NAND_GATE U248 ( .I1(n161), .I2(n267), .O(n265) );
  NAND_GATE U249 ( .I1(n22), .I2(N1248), .O(n264) );
  NAND3_GATE U250 ( .I1(n268), .I2(n269), .I3(n270), .O(n1501) );
  NAND_GATE U251 ( .I1(\pred_tab[2][BRA_ADR][5] ), .I2(n160), .O(n270) );
  NAND_GATE U252 ( .I1(n161), .I2(n271), .O(n269) );
  NAND_GATE U253 ( .I1(n22), .I2(N1249), .O(n268) );
  NAND3_GATE U254 ( .I1(n272), .I2(n273), .I3(n274), .O(n1502) );
  NAND_GATE U255 ( .I1(\pred_tab[2][BRA_ADR][6] ), .I2(n160), .O(n274) );
  NAND_GATE U256 ( .I1(n161), .I2(n275), .O(n273) );
  NAND_GATE U257 ( .I1(n21), .I2(N1250), .O(n272) );
  NAND3_GATE U258 ( .I1(n276), .I2(n277), .I3(n278), .O(n1503) );
  NAND_GATE U259 ( .I1(\pred_tab[2][BRA_ADR][7] ), .I2(n160), .O(n278) );
  NAND_GATE U260 ( .I1(n161), .I2(n279), .O(n277) );
  NAND_GATE U261 ( .I1(n21), .I2(N1251), .O(n276) );
  NAND3_GATE U262 ( .I1(n280), .I2(n281), .I3(n282), .O(n1504) );
  NAND_GATE U263 ( .I1(\pred_tab[2][BRA_ADR][8] ), .I2(n160), .O(n282) );
  NAND_GATE U264 ( .I1(n161), .I2(n283), .O(n281) );
  NAND_GATE U265 ( .I1(n21), .I2(N1252), .O(n280) );
  NAND3_GATE U266 ( .I1(n284), .I2(n285), .I3(n286), .O(n1505) );
  NAND_GATE U267 ( .I1(\pred_tab[2][BRA_ADR][9] ), .I2(n160), .O(n286) );
  NAND_GATE U268 ( .I1(n161), .I2(n287), .O(n285) );
  NAND_GATE U269 ( .I1(n21), .I2(N1253), .O(n284) );
  NAND3_GATE U270 ( .I1(n288), .I2(n289), .I3(n290), .O(n1506) );
  NAND_GATE U271 ( .I1(\pred_tab[3][BRA_ADR][0] ), .I2(n291), .O(n290) );
  NAND_GATE U272 ( .I1(n292), .I2(n293), .O(n289) );
  NAND_GATE U273 ( .I1(n294), .I2(N1244), .O(n288) );
  NAND3_GATE U274 ( .I1(n295), .I2(n296), .I3(n297), .O(n1507) );
  NAND_GATE U275 ( .I1(\pred_tab[3][BRA_ADR][10] ), .I2(n291), .O(n297) );
  NAND_GATE U276 ( .I1(n292), .I2(n298), .O(n296) );
  NAND_GATE U277 ( .I1(n294), .I2(N1254), .O(n295) );
  NAND3_GATE U278 ( .I1(n299), .I2(n300), .I3(n301), .O(n1508) );
  NAND_GATE U279 ( .I1(\pred_tab[3][BRA_ADR][11] ), .I2(n291), .O(n301) );
  NAND_GATE U280 ( .I1(n292), .I2(n302), .O(n300) );
  NAND_GATE U281 ( .I1(n294), .I2(N1255), .O(n299) );
  NAND3_GATE U282 ( .I1(n303), .I2(n304), .I3(n305), .O(n1509) );
  NAND_GATE U283 ( .I1(\pred_tab[3][BRA_ADR][12] ), .I2(n291), .O(n305) );
  NAND_GATE U284 ( .I1(n292), .I2(n306), .O(n304) );
  NAND_GATE U285 ( .I1(n294), .I2(N1256), .O(n303) );
  NAND3_GATE U286 ( .I1(n307), .I2(n308), .I3(n309), .O(n1510) );
  NAND_GATE U287 ( .I1(\pred_tab[3][BRA_ADR][13] ), .I2(n291), .O(n309) );
  NAND_GATE U288 ( .I1(n292), .I2(n310), .O(n308) );
  NAND_GATE U289 ( .I1(n294), .I2(N1257), .O(n307) );
  NAND3_GATE U290 ( .I1(n311), .I2(n312), .I3(n313), .O(n1511) );
  NAND_GATE U291 ( .I1(\pred_tab[3][BRA_ADR][14] ), .I2(n291), .O(n313) );
  NAND_GATE U292 ( .I1(n292), .I2(n314), .O(n312) );
  NAND_GATE U293 ( .I1(n294), .I2(N1258), .O(n311) );
  NAND3_GATE U294 ( .I1(n315), .I2(n316), .I3(n317), .O(n1512) );
  NAND_GATE U295 ( .I1(\pred_tab[3][BRA_ADR][15] ), .I2(n291), .O(n317) );
  NAND_GATE U296 ( .I1(n292), .I2(n318), .O(n316) );
  NAND_GATE U297 ( .I1(n294), .I2(N1259), .O(n315) );
  NAND3_GATE U298 ( .I1(n319), .I2(n320), .I3(n321), .O(n1513) );
  NAND_GATE U299 ( .I1(\pred_tab[3][BRA_ADR][16] ), .I2(n291), .O(n321) );
  NAND_GATE U300 ( .I1(n292), .I2(n322), .O(n320) );
  NAND_GATE U301 ( .I1(n294), .I2(N1260), .O(n319) );
  NAND3_GATE U302 ( .I1(n323), .I2(n324), .I3(n325), .O(n1514) );
  NAND_GATE U303 ( .I1(\pred_tab[3][BRA_ADR][17] ), .I2(n291), .O(n325) );
  NAND_GATE U304 ( .I1(n292), .I2(n326), .O(n324) );
  NAND_GATE U305 ( .I1(n294), .I2(N1261), .O(n323) );
  NAND3_GATE U306 ( .I1(n327), .I2(n328), .I3(n329), .O(n1515) );
  NAND_GATE U307 ( .I1(\pred_tab[3][BRA_ADR][18] ), .I2(n291), .O(n329) );
  NAND_GATE U308 ( .I1(n292), .I2(n330), .O(n328) );
  NAND_GATE U309 ( .I1(n16), .I2(N1262), .O(n327) );
  NAND3_GATE U310 ( .I1(n331), .I2(n332), .I3(n333), .O(n1516) );
  NAND_GATE U311 ( .I1(\pred_tab[3][BRA_ADR][19] ), .I2(n291), .O(n333) );
  NAND_GATE U312 ( .I1(n292), .I2(n334), .O(n332) );
  NAND_GATE U313 ( .I1(n17), .I2(N1263), .O(n331) );
  NAND3_GATE U314 ( .I1(n335), .I2(n336), .I3(n337), .O(n1517) );
  NAND_GATE U315 ( .I1(\pred_tab[3][BRA_ADR][1] ), .I2(n291), .O(n337) );
  NAND_GATE U316 ( .I1(n292), .I2(n338), .O(n336) );
  NAND_GATE U317 ( .I1(n14), .I2(N1245), .O(n335) );
  NAND3_GATE U318 ( .I1(n339), .I2(n340), .I3(n341), .O(n1518) );
  NAND_GATE U319 ( .I1(\pred_tab[3][BRA_ADR][20] ), .I2(n291), .O(n341) );
  NAND_GATE U320 ( .I1(n292), .I2(n342), .O(n340) );
  NAND_GATE U321 ( .I1(n15), .I2(N1264), .O(n339) );
  NAND3_GATE U322 ( .I1(n343), .I2(n344), .I3(n345), .O(n1519) );
  NAND_GATE U323 ( .I1(\pred_tab[3][BRA_ADR][21] ), .I2(n291), .O(n345) );
  NAND_GATE U324 ( .I1(n292), .I2(n346), .O(n344) );
  NAND_GATE U325 ( .I1(n294), .I2(N1265), .O(n343) );
  NAND3_GATE U326 ( .I1(n347), .I2(n348), .I3(n349), .O(n1520) );
  NAND_GATE U327 ( .I1(\pred_tab[3][BRA_ADR][22] ), .I2(n291), .O(n349) );
  NAND_GATE U328 ( .I1(n292), .I2(n350), .O(n348) );
  NAND_GATE U329 ( .I1(n294), .I2(N1266), .O(n347) );
  NAND3_GATE U330 ( .I1(n351), .I2(n352), .I3(n353), .O(n1521) );
  NAND_GATE U331 ( .I1(\pred_tab[3][BRA_ADR][23] ), .I2(n291), .O(n353) );
  NAND_GATE U332 ( .I1(n292), .I2(n354), .O(n352) );
  NAND_GATE U333 ( .I1(n16), .I2(N1267), .O(n351) );
  NAND3_GATE U334 ( .I1(n355), .I2(n356), .I3(n357), .O(n1522) );
  NAND_GATE U335 ( .I1(\pred_tab[3][BRA_ADR][24] ), .I2(n291), .O(n357) );
  NAND_GATE U336 ( .I1(n292), .I2(n358), .O(n356) );
  NAND_GATE U337 ( .I1(n17), .I2(N1268), .O(n355) );
  NAND3_GATE U338 ( .I1(n359), .I2(n360), .I3(n361), .O(n1523) );
  NAND_GATE U339 ( .I1(\pred_tab[3][BRA_ADR][25] ), .I2(n291), .O(n361) );
  NAND_GATE U340 ( .I1(n292), .I2(n362), .O(n360) );
  NAND_GATE U341 ( .I1(n14), .I2(N1269), .O(n359) );
  NAND3_GATE U342 ( .I1(n363), .I2(n364), .I3(n365), .O(n1524) );
  NAND_GATE U343 ( .I1(\pred_tab[3][BRA_ADR][26] ), .I2(n291), .O(n365) );
  NAND_GATE U344 ( .I1(n292), .I2(n366), .O(n364) );
  NAND_GATE U345 ( .I1(n15), .I2(N1270), .O(n363) );
  NAND3_GATE U346 ( .I1(n367), .I2(n368), .I3(n369), .O(n1525) );
  NAND_GATE U347 ( .I1(\pred_tab[3][BRA_ADR][27] ), .I2(n291), .O(n369) );
  NAND_GATE U348 ( .I1(n292), .I2(n370), .O(n368) );
  NAND_GATE U349 ( .I1(n17), .I2(N1271), .O(n367) );
  NAND3_GATE U350 ( .I1(n371), .I2(n372), .I3(n373), .O(n1526) );
  NAND_GATE U351 ( .I1(\pred_tab[3][BRA_ADR][28] ), .I2(n291), .O(n373) );
  NAND_GATE U352 ( .I1(n292), .I2(n374), .O(n372) );
  NAND_GATE U353 ( .I1(n17), .I2(N1272), .O(n371) );
  NAND3_GATE U354 ( .I1(n375), .I2(n376), .I3(n377), .O(n1527) );
  NAND_GATE U355 ( .I1(\pred_tab[3][BRA_ADR][29] ), .I2(n291), .O(n377) );
  NAND_GATE U356 ( .I1(n292), .I2(n378), .O(n376) );
  NAND_GATE U357 ( .I1(n17), .I2(N1273), .O(n375) );
  NAND3_GATE U358 ( .I1(n379), .I2(n380), .I3(n381), .O(n1528) );
  NAND_GATE U359 ( .I1(\pred_tab[3][BRA_ADR][2] ), .I2(n291), .O(n381) );
  NAND_GATE U360 ( .I1(n292), .I2(n382), .O(n380) );
  NAND_GATE U361 ( .I1(n17), .I2(N1246), .O(n379) );
  NAND3_GATE U362 ( .I1(n383), .I2(n384), .I3(n385), .O(n1529) );
  NAND_GATE U363 ( .I1(\pred_tab[3][BRA_ADR][30] ), .I2(n291), .O(n385) );
  NAND_GATE U364 ( .I1(n292), .I2(n386), .O(n384) );
  NAND_GATE U365 ( .I1(n17), .I2(N1274), .O(n383) );
  NAND3_GATE U366 ( .I1(n387), .I2(n388), .I3(n389), .O(n1530) );
  NAND_GATE U367 ( .I1(\pred_tab[3][BRA_ADR][31] ), .I2(n291), .O(n389) );
  NAND_GATE U368 ( .I1(n292), .I2(n390), .O(n388) );
  NAND_GATE U369 ( .I1(n17), .I2(N1275), .O(n387) );
  NAND3_GATE U370 ( .I1(n391), .I2(n392), .I3(n393), .O(n1531) );
  NAND_GATE U371 ( .I1(\pred_tab[3][BRA_ADR][3] ), .I2(n291), .O(n393) );
  NAND_GATE U372 ( .I1(n292), .I2(n394), .O(n392) );
  NAND_GATE U373 ( .I1(n17), .I2(N1247), .O(n391) );
  NAND3_GATE U374 ( .I1(n395), .I2(n396), .I3(n397), .O(n1532) );
  NAND_GATE U375 ( .I1(\pred_tab[3][BRA_ADR][4] ), .I2(n291), .O(n397) );
  NAND_GATE U376 ( .I1(n292), .I2(n398), .O(n396) );
  NAND_GATE U377 ( .I1(n17), .I2(N1248), .O(n395) );
  NAND3_GATE U378 ( .I1(n399), .I2(n400), .I3(n401), .O(n1533) );
  NAND_GATE U379 ( .I1(\pred_tab[3][BRA_ADR][5] ), .I2(n291), .O(n401) );
  NAND_GATE U380 ( .I1(n292), .I2(n402), .O(n400) );
  NAND_GATE U381 ( .I1(n17), .I2(N1249), .O(n399) );
  NAND3_GATE U382 ( .I1(n403), .I2(n404), .I3(n405), .O(n1534) );
  NAND_GATE U383 ( .I1(\pred_tab[3][BRA_ADR][6] ), .I2(n291), .O(n405) );
  NAND_GATE U384 ( .I1(n292), .I2(n406), .O(n404) );
  NAND_GATE U385 ( .I1(n16), .I2(N1250), .O(n403) );
  NAND3_GATE U386 ( .I1(n407), .I2(n408), .I3(n409), .O(n1535) );
  NAND_GATE U387 ( .I1(\pred_tab[3][BRA_ADR][7] ), .I2(n291), .O(n409) );
  NAND_GATE U388 ( .I1(n292), .I2(n410), .O(n408) );
  NAND_GATE U389 ( .I1(n16), .I2(N1251), .O(n407) );
  NAND3_GATE U390 ( .I1(n411), .I2(n412), .I3(n413), .O(n1536) );
  NAND_GATE U391 ( .I1(\pred_tab[3][BRA_ADR][8] ), .I2(n291), .O(n413) );
  NAND_GATE U392 ( .I1(n292), .I2(n414), .O(n412) );
  NAND_GATE U393 ( .I1(n16), .I2(N1252), .O(n411) );
  NAND3_GATE U394 ( .I1(n415), .I2(n416), .I3(n417), .O(n1537) );
  NAND_GATE U395 ( .I1(\pred_tab[3][BRA_ADR][9] ), .I2(n291), .O(n417) );
  NAND_GATE U396 ( .I1(n292), .I2(n418), .O(n416) );
  NAND_GATE U397 ( .I1(n16), .I2(N1253), .O(n415) );
  NAND3_GATE U398 ( .I1(n419), .I2(n420), .I3(n421), .O(n1538) );
  NAND_GATE U399 ( .I1(\pred_tab[1][BRA_ADR][0] ), .I2(n33), .O(n421) );
  NAND_GATE U400 ( .I1(n34), .I2(n422), .O(n420) );
  NAND_GATE U401 ( .I1(N1244), .I2(n26), .O(n419) );
  NAND_GATE U402 ( .I1(n423), .I2(n424), .O(n1539) );
  NAND3_GATE U403 ( .I1(n425), .I2(EX_bra_confirm), .I3(n161), .O(n424) );
  AND_GATE U404 ( .I1(n426), .I2(n447), .O(n161) );
  NAND_GATE U405 ( .I1(\pred_tab[2][LAST_BRA] ), .I2(n428), .O(n423) );
  OR_GATE U406 ( .I1(n160), .I2(n429), .O(n428) );
  NOR_GATE U407 ( .I1(n425), .I2(n28), .O(n429) );
  NAND_GATE U408 ( .I1(n434), .I2(n430), .O(n160) );
  OR_GATE U409 ( .I1(n28), .I2(EX_uncleared), .O(n430) );
  NAND_GATE U410 ( .I1(n431), .I2(n432), .O(n1540) );
  NAND3_GATE U411 ( .I1(n433), .I2(EX_bra_confirm), .I3(n34), .O(n432) );
  AND_GATE U412 ( .I1(n426), .I2(n577), .O(n34) );
  NAND_GATE U413 ( .I1(\pred_tab[1][LAST_BRA] ), .I2(n435), .O(n431) );
  OR_GATE U414 ( .I1(n33), .I2(n436), .O(n435) );
  NOR_GATE U415 ( .I1(n433), .I2(n29), .O(n436) );
  NAND_GATE U416 ( .I1(n434), .I2(n437), .O(n33) );
  OR_GATE U417 ( .I1(n29), .I2(EX_uncleared), .O(n437) );
  NAND_GATE U418 ( .I1(n438), .I2(n439), .O(n1541) );
  NAND3_GATE U419 ( .I1(EX_bra_confirm), .I2(n440), .I3(n292), .O(n439) );
  AND_GATE U420 ( .I1(n426), .I2(n441), .O(n292) );
  AND_GATE U421 ( .I1(EX_uncleared), .I2(n434), .O(n426) );
  NAND_GATE U422 ( .I1(\pred_tab[3][LAST_BRA] ), .I2(n442), .O(n438) );
  OR_GATE U423 ( .I1(n291), .I2(n443), .O(n442) );
  NOR_GATE U424 ( .I1(n642), .I2(n440), .O(n443) );
  NAND_GATE U425 ( .I1(n434), .I2(n444), .O(n291) );
  OR_GATE U426 ( .I1(n642), .I2(EX_uncleared), .O(n444) );
  NAND_GATE U427 ( .I1(n445), .I2(n446), .O(n1542) );
  NAND_GATE U428 ( .I1(DI_adr[9]), .I2(n26), .O(n446) );
  NAND_GATE U429 ( .I1(\pred_tab[1][CODE_ADR][9] ), .I2(n427), .O(n445) );
  NAND_GATE U430 ( .I1(n448), .I2(n449), .O(n1543) );
  NAND_GATE U431 ( .I1(DI_adr[8]), .I2(n26), .O(n449) );
  NAND_GATE U432 ( .I1(\pred_tab[1][CODE_ADR][8] ), .I2(n427), .O(n448) );
  NAND_GATE U433 ( .I1(n450), .I2(n451), .O(n1544) );
  NAND_GATE U434 ( .I1(DI_adr[7]), .I2(n26), .O(n451) );
  NAND_GATE U435 ( .I1(\pred_tab[1][CODE_ADR][7] ), .I2(n427), .O(n450) );
  NAND_GATE U436 ( .I1(n452), .I2(n453), .O(n1545) );
  NAND_GATE U437 ( .I1(DI_adr[6]), .I2(n26), .O(n453) );
  NAND_GATE U438 ( .I1(\pred_tab[1][CODE_ADR][6] ), .I2(n427), .O(n452) );
  NAND_GATE U439 ( .I1(n454), .I2(n455), .O(n1546) );
  NAND_GATE U440 ( .I1(DI_adr[5]), .I2(n26), .O(n455) );
  NAND_GATE U441 ( .I1(\pred_tab[1][CODE_ADR][5] ), .I2(n427), .O(n454) );
  NAND_GATE U442 ( .I1(n456), .I2(n457), .O(n1547) );
  NAND_GATE U443 ( .I1(DI_adr[4]), .I2(n26), .O(n457) );
  NAND_GATE U444 ( .I1(\pred_tab[1][CODE_ADR][4] ), .I2(n427), .O(n456) );
  NAND_GATE U445 ( .I1(n458), .I2(n459), .O(n1548) );
  NAND_GATE U446 ( .I1(DI_adr[3]), .I2(n27), .O(n459) );
  NAND_GATE U447 ( .I1(\pred_tab[1][CODE_ADR][3] ), .I2(n427), .O(n458) );
  NAND_GATE U448 ( .I1(n460), .I2(n461), .O(n1549) );
  NAND_GATE U449 ( .I1(DI_adr[31]), .I2(n24), .O(n461) );
  NAND_GATE U450 ( .I1(\pred_tab[1][CODE_ADR][31] ), .I2(n427), .O(n460) );
  NAND_GATE U451 ( .I1(n462), .I2(n463), .O(n1550) );
  NAND_GATE U452 ( .I1(DI_adr[30]), .I2(n25), .O(n463) );
  NAND_GATE U453 ( .I1(\pred_tab[1][CODE_ADR][30] ), .I2(n427), .O(n462) );
  NAND_GATE U454 ( .I1(n464), .I2(n465), .O(n1551) );
  NAND_GATE U455 ( .I1(DI_adr[2]), .I2(n36), .O(n465) );
  NAND_GATE U456 ( .I1(\pred_tab[1][CODE_ADR][2] ), .I2(n427), .O(n464) );
  NAND_GATE U457 ( .I1(n466), .I2(n467), .O(n1552) );
  NAND_GATE U458 ( .I1(DI_adr[29]), .I2(n26), .O(n467) );
  NAND_GATE U459 ( .I1(\pred_tab[1][CODE_ADR][29] ), .I2(n427), .O(n466) );
  NAND_GATE U460 ( .I1(n468), .I2(n469), .O(n1553) );
  NAND_GATE U461 ( .I1(DI_adr[28]), .I2(n27), .O(n469) );
  NAND_GATE U462 ( .I1(\pred_tab[1][CODE_ADR][28] ), .I2(n427), .O(n468) );
  NAND_GATE U463 ( .I1(n470), .I2(n471), .O(n1554) );
  NAND_GATE U464 ( .I1(DI_adr[27]), .I2(n24), .O(n471) );
  NAND_GATE U465 ( .I1(\pred_tab[1][CODE_ADR][27] ), .I2(n427), .O(n470) );
  NAND_GATE U466 ( .I1(n472), .I2(n473), .O(n1555) );
  NAND_GATE U467 ( .I1(DI_adr[26]), .I2(n25), .O(n473) );
  NAND_GATE U468 ( .I1(\pred_tab[1][CODE_ADR][26] ), .I2(n427), .O(n472) );
  NAND_GATE U469 ( .I1(n474), .I2(n475), .O(n1556) );
  NAND_GATE U470 ( .I1(DI_adr[25]), .I2(n25), .O(n475) );
  NAND_GATE U471 ( .I1(\pred_tab[1][CODE_ADR][25] ), .I2(n427), .O(n474) );
  NAND_GATE U472 ( .I1(n476), .I2(n477), .O(n1557) );
  NAND_GATE U473 ( .I1(DI_adr[24]), .I2(n25), .O(n477) );
  NAND_GATE U474 ( .I1(\pred_tab[1][CODE_ADR][24] ), .I2(n427), .O(n476) );
  NAND_GATE U475 ( .I1(n478), .I2(n479), .O(n1558) );
  NAND_GATE U476 ( .I1(DI_adr[23]), .I2(n25), .O(n479) );
  NAND_GATE U477 ( .I1(\pred_tab[1][CODE_ADR][23] ), .I2(n427), .O(n478) );
  NAND_GATE U478 ( .I1(n480), .I2(n481), .O(n1559) );
  NAND_GATE U479 ( .I1(DI_adr[22]), .I2(n25), .O(n481) );
  NAND_GATE U480 ( .I1(\pred_tab[1][CODE_ADR][22] ), .I2(n427), .O(n480) );
  NAND_GATE U481 ( .I1(n482), .I2(n483), .O(n1560) );
  NAND_GATE U482 ( .I1(DI_adr[21]), .I2(n25), .O(n483) );
  NAND_GATE U483 ( .I1(\pred_tab[1][CODE_ADR][21] ), .I2(n427), .O(n482) );
  NAND_GATE U484 ( .I1(n484), .I2(n485), .O(n1561) );
  NAND_GATE U485 ( .I1(DI_adr[20]), .I2(n25), .O(n485) );
  NAND_GATE U486 ( .I1(\pred_tab[1][CODE_ADR][20] ), .I2(n427), .O(n484) );
  NAND_GATE U487 ( .I1(n486), .I2(n487), .O(n1562) );
  NAND_GATE U488 ( .I1(DI_adr[1]), .I2(n25), .O(n487) );
  NAND_GATE U489 ( .I1(\pred_tab[1][CODE_ADR][1] ), .I2(n427), .O(n486) );
  NAND_GATE U490 ( .I1(n488), .I2(n489), .O(n1563) );
  NAND_GATE U491 ( .I1(DI_adr[19]), .I2(n25), .O(n489) );
  NAND_GATE U492 ( .I1(\pred_tab[1][CODE_ADR][19] ), .I2(n427), .O(n488) );
  NAND_GATE U493 ( .I1(n490), .I2(n491), .O(n1564) );
  NAND_GATE U494 ( .I1(DI_adr[18]), .I2(n25), .O(n491) );
  NAND_GATE U495 ( .I1(\pred_tab[1][CODE_ADR][18] ), .I2(n427), .O(n490) );
  NAND_GATE U496 ( .I1(n492), .I2(n493), .O(n1565) );
  NAND_GATE U497 ( .I1(DI_adr[17]), .I2(n24), .O(n493) );
  NAND_GATE U498 ( .I1(\pred_tab[1][CODE_ADR][17] ), .I2(n427), .O(n492) );
  NAND_GATE U499 ( .I1(n494), .I2(n495), .O(n1566) );
  NAND_GATE U500 ( .I1(DI_adr[16]), .I2(n24), .O(n495) );
  NAND_GATE U501 ( .I1(\pred_tab[1][CODE_ADR][16] ), .I2(n427), .O(n494) );
  NAND_GATE U502 ( .I1(n496), .I2(n497), .O(n1567) );
  NAND_GATE U503 ( .I1(DI_adr[15]), .I2(n24), .O(n497) );
  NAND_GATE U504 ( .I1(\pred_tab[1][CODE_ADR][15] ), .I2(n427), .O(n496) );
  NAND_GATE U505 ( .I1(n498), .I2(n499), .O(n1568) );
  NAND_GATE U506 ( .I1(DI_adr[14]), .I2(n24), .O(n499) );
  NAND_GATE U507 ( .I1(\pred_tab[1][CODE_ADR][14] ), .I2(n427), .O(n498) );
  NAND_GATE U508 ( .I1(n500), .I2(n501), .O(n1569) );
  NAND_GATE U509 ( .I1(DI_adr[13]), .I2(n24), .O(n501) );
  NAND_GATE U510 ( .I1(\pred_tab[1][CODE_ADR][13] ), .I2(n427), .O(n500) );
  NAND_GATE U511 ( .I1(n502), .I2(n503), .O(n1570) );
  NAND_GATE U512 ( .I1(DI_adr[12]), .I2(n24), .O(n503) );
  NAND_GATE U513 ( .I1(\pred_tab[1][CODE_ADR][12] ), .I2(n427), .O(n502) );
  NAND_GATE U514 ( .I1(n504), .I2(n505), .O(n1571) );
  NAND_GATE U515 ( .I1(DI_adr[11]), .I2(n24), .O(n505) );
  NAND_GATE U516 ( .I1(\pred_tab[1][CODE_ADR][11] ), .I2(n427), .O(n504) );
  NAND_GATE U517 ( .I1(n506), .I2(n507), .O(n1572) );
  NAND_GATE U518 ( .I1(DI_adr[10]), .I2(n24), .O(n507) );
  NAND_GATE U519 ( .I1(\pred_tab[1][CODE_ADR][10] ), .I2(n427), .O(n506) );
  NAND_GATE U520 ( .I1(n508), .I2(n509), .O(n1573) );
  NAND_GATE U521 ( .I1(DI_adr[0]), .I2(n24), .O(n509) );
  NAND_GATE U522 ( .I1(\pred_tab[1][CODE_ADR][0] ), .I2(n427), .O(n508) );
  AND_GATE U524 ( .I1(n29), .I2(n434), .O(n36) );
  NAND_GATE U525 ( .I1(n510), .I2(n511), .O(n1574) );
  NAND_GATE U526 ( .I1(DI_adr[9]), .I2(n16), .O(n511) );
  NAND_GATE U527 ( .I1(\pred_tab[3][CODE_ADR][9] ), .I2(n18), .O(n510) );
  NAND_GATE U528 ( .I1(n513), .I2(n514), .O(n1575) );
  NAND_GATE U529 ( .I1(DI_adr[8]), .I2(n16), .O(n514) );
  NAND_GATE U530 ( .I1(\pred_tab[3][CODE_ADR][8] ), .I2(n18), .O(n513) );
  NAND_GATE U531 ( .I1(n515), .I2(n516), .O(n1576) );
  NAND_GATE U532 ( .I1(DI_adr[7]), .I2(n16), .O(n516) );
  NAND_GATE U533 ( .I1(\pred_tab[3][CODE_ADR][7] ), .I2(n18), .O(n515) );
  NAND_GATE U534 ( .I1(n517), .I2(n518), .O(n1577) );
  NAND_GATE U535 ( .I1(DI_adr[6]), .I2(n16), .O(n518) );
  NAND_GATE U536 ( .I1(\pred_tab[3][CODE_ADR][6] ), .I2(n18), .O(n517) );
  NAND_GATE U537 ( .I1(n519), .I2(n520), .O(n1578) );
  NAND_GATE U538 ( .I1(DI_adr[5]), .I2(n16), .O(n520) );
  NAND_GATE U539 ( .I1(\pred_tab[3][CODE_ADR][5] ), .I2(n18), .O(n519) );
  NAND_GATE U540 ( .I1(n521), .I2(n522), .O(n1579) );
  NAND_GATE U541 ( .I1(DI_adr[4]), .I2(n16), .O(n522) );
  NAND_GATE U542 ( .I1(\pred_tab[3][CODE_ADR][4] ), .I2(n18), .O(n521) );
  NAND_GATE U543 ( .I1(n523), .I2(n524), .O(n1580) );
  NAND_GATE U544 ( .I1(DI_adr[3]), .I2(n17), .O(n524) );
  NAND_GATE U545 ( .I1(\pred_tab[3][CODE_ADR][3] ), .I2(n18), .O(n523) );
  NAND_GATE U546 ( .I1(n525), .I2(n526), .O(n1581) );
  NAND_GATE U547 ( .I1(DI_adr[31]), .I2(n14), .O(n526) );
  NAND_GATE U548 ( .I1(\pred_tab[3][CODE_ADR][31] ), .I2(n18), .O(n525) );
  NAND_GATE U549 ( .I1(n527), .I2(n528), .O(n1582) );
  NAND_GATE U550 ( .I1(DI_adr[30]), .I2(n15), .O(n528) );
  NAND_GATE U551 ( .I1(\pred_tab[3][CODE_ADR][30] ), .I2(n18), .O(n527) );
  NAND_GATE U552 ( .I1(n529), .I2(n530), .O(n1583) );
  NAND_GATE U553 ( .I1(DI_adr[2]), .I2(n294), .O(n530) );
  NAND_GATE U554 ( .I1(\pred_tab[3][CODE_ADR][2] ), .I2(n18), .O(n529) );
  NAND_GATE U555 ( .I1(n531), .I2(n532), .O(n1584) );
  NAND_GATE U556 ( .I1(DI_adr[29]), .I2(n16), .O(n532) );
  NAND_GATE U557 ( .I1(\pred_tab[3][CODE_ADR][29] ), .I2(n18), .O(n531) );
  NAND_GATE U558 ( .I1(n533), .I2(n534), .O(n1585) );
  NAND_GATE U559 ( .I1(DI_adr[28]), .I2(n17), .O(n534) );
  NAND_GATE U560 ( .I1(\pred_tab[3][CODE_ADR][28] ), .I2(n18), .O(n533) );
  NAND_GATE U561 ( .I1(n535), .I2(n536), .O(n1586) );
  NAND_GATE U562 ( .I1(DI_adr[27]), .I2(n14), .O(n536) );
  NAND_GATE U563 ( .I1(\pred_tab[3][CODE_ADR][27] ), .I2(n18), .O(n535) );
  NAND_GATE U564 ( .I1(n537), .I2(n538), .O(n1587) );
  NAND_GATE U565 ( .I1(DI_adr[26]), .I2(n15), .O(n538) );
  NAND_GATE U566 ( .I1(\pred_tab[3][CODE_ADR][26] ), .I2(n18), .O(n537) );
  NAND_GATE U567 ( .I1(n539), .I2(n540), .O(n1588) );
  NAND_GATE U568 ( .I1(DI_adr[25]), .I2(n15), .O(n540) );
  NAND_GATE U569 ( .I1(\pred_tab[3][CODE_ADR][25] ), .I2(n18), .O(n539) );
  NAND_GATE U570 ( .I1(n541), .I2(n542), .O(n1589) );
  NAND_GATE U571 ( .I1(DI_adr[24]), .I2(n15), .O(n542) );
  NAND_GATE U572 ( .I1(\pred_tab[3][CODE_ADR][24] ), .I2(n18), .O(n541) );
  NAND_GATE U573 ( .I1(n543), .I2(n544), .O(n1590) );
  NAND_GATE U574 ( .I1(DI_adr[23]), .I2(n15), .O(n544) );
  NAND_GATE U575 ( .I1(\pred_tab[3][CODE_ADR][23] ), .I2(n18), .O(n543) );
  NAND_GATE U576 ( .I1(n545), .I2(n546), .O(n1591) );
  NAND_GATE U577 ( .I1(DI_adr[22]), .I2(n15), .O(n546) );
  NAND_GATE U578 ( .I1(\pred_tab[3][CODE_ADR][22] ), .I2(n18), .O(n545) );
  NAND_GATE U579 ( .I1(n547), .I2(n548), .O(n1592) );
  NAND_GATE U580 ( .I1(DI_adr[21]), .I2(n15), .O(n548) );
  NAND_GATE U581 ( .I1(\pred_tab[3][CODE_ADR][21] ), .I2(n18), .O(n547) );
  NAND_GATE U582 ( .I1(n549), .I2(n550), .O(n1593) );
  NAND_GATE U583 ( .I1(DI_adr[20]), .I2(n15), .O(n550) );
  NAND_GATE U584 ( .I1(\pred_tab[3][CODE_ADR][20] ), .I2(n18), .O(n549) );
  NAND_GATE U585 ( .I1(n551), .I2(n552), .O(n1594) );
  NAND_GATE U586 ( .I1(DI_adr[1]), .I2(n15), .O(n552) );
  NAND_GATE U587 ( .I1(\pred_tab[3][CODE_ADR][1] ), .I2(n18), .O(n551) );
  NAND_GATE U588 ( .I1(n553), .I2(n554), .O(n1595) );
  NAND_GATE U589 ( .I1(DI_adr[19]), .I2(n15), .O(n554) );
  NAND_GATE U590 ( .I1(\pred_tab[3][CODE_ADR][19] ), .I2(n18), .O(n553) );
  NAND_GATE U591 ( .I1(n555), .I2(n556), .O(n1596) );
  NAND_GATE U592 ( .I1(DI_adr[18]), .I2(n15), .O(n556) );
  NAND_GATE U593 ( .I1(\pred_tab[3][CODE_ADR][18] ), .I2(n18), .O(n555) );
  NAND_GATE U594 ( .I1(n557), .I2(n558), .O(n1597) );
  NAND_GATE U595 ( .I1(DI_adr[17]), .I2(n14), .O(n558) );
  NAND_GATE U596 ( .I1(\pred_tab[3][CODE_ADR][17] ), .I2(n18), .O(n557) );
  NAND_GATE U597 ( .I1(n559), .I2(n560), .O(n1598) );
  NAND_GATE U598 ( .I1(DI_adr[16]), .I2(n14), .O(n560) );
  NAND_GATE U599 ( .I1(\pred_tab[3][CODE_ADR][16] ), .I2(n18), .O(n559) );
  NAND_GATE U600 ( .I1(n561), .I2(n562), .O(n1599) );
  NAND_GATE U601 ( .I1(DI_adr[15]), .I2(n14), .O(n562) );
  NAND_GATE U602 ( .I1(\pred_tab[3][CODE_ADR][15] ), .I2(n18), .O(n561) );
  NAND_GATE U603 ( .I1(n563), .I2(n564), .O(n1600) );
  NAND_GATE U604 ( .I1(DI_adr[14]), .I2(n14), .O(n564) );
  NAND_GATE U605 ( .I1(\pred_tab[3][CODE_ADR][14] ), .I2(n18), .O(n563) );
  NAND_GATE U606 ( .I1(n565), .I2(n566), .O(n1601) );
  NAND_GATE U607 ( .I1(DI_adr[13]), .I2(n14), .O(n566) );
  NAND_GATE U608 ( .I1(\pred_tab[3][CODE_ADR][13] ), .I2(n18), .O(n565) );
  NAND_GATE U609 ( .I1(n567), .I2(n568), .O(n1602) );
  NAND_GATE U610 ( .I1(DI_adr[12]), .I2(n14), .O(n568) );
  NAND_GATE U611 ( .I1(\pred_tab[3][CODE_ADR][12] ), .I2(n18), .O(n567) );
  NAND_GATE U612 ( .I1(n569), .I2(n570), .O(n1603) );
  NAND_GATE U613 ( .I1(DI_adr[11]), .I2(n14), .O(n570) );
  NAND_GATE U614 ( .I1(\pred_tab[3][CODE_ADR][11] ), .I2(n18), .O(n569) );
  NAND_GATE U615 ( .I1(n571), .I2(n572), .O(n1604) );
  NAND_GATE U616 ( .I1(DI_adr[10]), .I2(n14), .O(n572) );
  NAND_GATE U617 ( .I1(\pred_tab[3][CODE_ADR][10] ), .I2(n18), .O(n571) );
  NAND_GATE U618 ( .I1(n573), .I2(n574), .O(n1605) );
  NAND_GATE U619 ( .I1(DI_adr[0]), .I2(n14), .O(n574) );
  NAND_GATE U620 ( .I1(\pred_tab[3][CODE_ADR][0] ), .I2(n18), .O(n573) );
  AND_GATE U622 ( .I1(n642), .I2(n434), .O(n294) );
  NAND_GATE U623 ( .I1(n575), .I2(n576), .O(n1606) );
  NAND_GATE U624 ( .I1(DI_adr[9]), .I2(n21), .O(n576) );
  NAND_GATE U625 ( .I1(\pred_tab[2][CODE_ADR][9] ), .I2(n23), .O(n575) );
  NAND_GATE U626 ( .I1(n578), .I2(n579), .O(n1607) );
  NAND_GATE U627 ( .I1(DI_adr[8]), .I2(n21), .O(n579) );
  NAND_GATE U628 ( .I1(\pred_tab[2][CODE_ADR][8] ), .I2(n23), .O(n578) );
  NAND_GATE U629 ( .I1(n580), .I2(n581), .O(n1608) );
  NAND_GATE U630 ( .I1(DI_adr[7]), .I2(n21), .O(n581) );
  NAND_GATE U631 ( .I1(\pred_tab[2][CODE_ADR][7] ), .I2(n23), .O(n580) );
  NAND_GATE U632 ( .I1(n582), .I2(n583), .O(n1609) );
  NAND_GATE U633 ( .I1(DI_adr[6]), .I2(n21), .O(n583) );
  NAND_GATE U634 ( .I1(\pred_tab[2][CODE_ADR][6] ), .I2(n23), .O(n582) );
  NAND_GATE U635 ( .I1(n584), .I2(n585), .O(n1610) );
  NAND_GATE U636 ( .I1(DI_adr[5]), .I2(n21), .O(n585) );
  NAND_GATE U637 ( .I1(\pred_tab[2][CODE_ADR][5] ), .I2(n23), .O(n584) );
  NAND_GATE U638 ( .I1(n586), .I2(n587), .O(n1611) );
  NAND_GATE U639 ( .I1(DI_adr[4]), .I2(n21), .O(n587) );
  NAND_GATE U640 ( .I1(\pred_tab[2][CODE_ADR][4] ), .I2(n23), .O(n586) );
  NAND_GATE U641 ( .I1(n588), .I2(n589), .O(n1612) );
  NAND_GATE U642 ( .I1(DI_adr[3]), .I2(n22), .O(n589) );
  NAND_GATE U643 ( .I1(\pred_tab[2][CODE_ADR][3] ), .I2(n23), .O(n588) );
  NAND_GATE U644 ( .I1(n590), .I2(n591), .O(n1613) );
  NAND_GATE U645 ( .I1(DI_adr[31]), .I2(n19), .O(n591) );
  NAND_GATE U646 ( .I1(\pred_tab[2][CODE_ADR][31] ), .I2(n23), .O(n590) );
  NAND_GATE U647 ( .I1(n592), .I2(n593), .O(n1614) );
  NAND_GATE U648 ( .I1(DI_adr[30]), .I2(n20), .O(n593) );
  NAND_GATE U649 ( .I1(\pred_tab[2][CODE_ADR][30] ), .I2(n23), .O(n592) );
  NAND_GATE U650 ( .I1(n594), .I2(n595), .O(n1615) );
  NAND_GATE U651 ( .I1(DI_adr[2]), .I2(n163), .O(n595) );
  NAND_GATE U652 ( .I1(\pred_tab[2][CODE_ADR][2] ), .I2(n23), .O(n594) );
  NAND_GATE U653 ( .I1(n596), .I2(n597), .O(n1616) );
  NAND_GATE U654 ( .I1(DI_adr[29]), .I2(n21), .O(n597) );
  NAND_GATE U655 ( .I1(\pred_tab[2][CODE_ADR][29] ), .I2(n23), .O(n596) );
  NAND_GATE U656 ( .I1(n598), .I2(n599), .O(n1617) );
  NAND_GATE U657 ( .I1(DI_adr[28]), .I2(n22), .O(n599) );
  NAND_GATE U658 ( .I1(\pred_tab[2][CODE_ADR][28] ), .I2(n23), .O(n598) );
  NAND_GATE U659 ( .I1(n600), .I2(n601), .O(n1618) );
  NAND_GATE U660 ( .I1(DI_adr[27]), .I2(n19), .O(n601) );
  NAND_GATE U661 ( .I1(\pred_tab[2][CODE_ADR][27] ), .I2(n23), .O(n600) );
  NAND_GATE U662 ( .I1(n602), .I2(n603), .O(n1619) );
  NAND_GATE U663 ( .I1(DI_adr[26]), .I2(n20), .O(n603) );
  NAND_GATE U664 ( .I1(\pred_tab[2][CODE_ADR][26] ), .I2(n23), .O(n602) );
  NAND_GATE U665 ( .I1(n604), .I2(n605), .O(n1620) );
  NAND_GATE U666 ( .I1(DI_adr[25]), .I2(n20), .O(n605) );
  NAND_GATE U667 ( .I1(\pred_tab[2][CODE_ADR][25] ), .I2(n23), .O(n604) );
  NAND_GATE U668 ( .I1(n606), .I2(n607), .O(n1621) );
  NAND_GATE U669 ( .I1(DI_adr[24]), .I2(n20), .O(n607) );
  NAND_GATE U670 ( .I1(\pred_tab[2][CODE_ADR][24] ), .I2(n23), .O(n606) );
  NAND_GATE U671 ( .I1(n608), .I2(n609), .O(n1622) );
  NAND_GATE U672 ( .I1(DI_adr[23]), .I2(n20), .O(n609) );
  NAND_GATE U673 ( .I1(\pred_tab[2][CODE_ADR][23] ), .I2(n23), .O(n608) );
  NAND_GATE U674 ( .I1(n610), .I2(n611), .O(n1623) );
  NAND_GATE U675 ( .I1(DI_adr[22]), .I2(n20), .O(n611) );
  NAND_GATE U676 ( .I1(\pred_tab[2][CODE_ADR][22] ), .I2(n23), .O(n610) );
  NAND_GATE U677 ( .I1(n612), .I2(n613), .O(n1624) );
  NAND_GATE U678 ( .I1(DI_adr[21]), .I2(n20), .O(n613) );
  NAND_GATE U679 ( .I1(\pred_tab[2][CODE_ADR][21] ), .I2(n23), .O(n612) );
  NAND_GATE U680 ( .I1(n614), .I2(n615), .O(n1625) );
  NAND_GATE U681 ( .I1(DI_adr[20]), .I2(n20), .O(n615) );
  NAND_GATE U682 ( .I1(\pred_tab[2][CODE_ADR][20] ), .I2(n23), .O(n614) );
  NAND_GATE U683 ( .I1(n616), .I2(n617), .O(n1626) );
  NAND_GATE U684 ( .I1(DI_adr[1]), .I2(n20), .O(n617) );
  NAND_GATE U685 ( .I1(\pred_tab[2][CODE_ADR][1] ), .I2(n23), .O(n616) );
  NAND_GATE U686 ( .I1(n618), .I2(n619), .O(n1627) );
  NAND_GATE U687 ( .I1(DI_adr[19]), .I2(n20), .O(n619) );
  NAND_GATE U688 ( .I1(\pred_tab[2][CODE_ADR][19] ), .I2(n23), .O(n618) );
  NAND_GATE U689 ( .I1(n620), .I2(n621), .O(n1628) );
  NAND_GATE U690 ( .I1(DI_adr[18]), .I2(n20), .O(n621) );
  NAND_GATE U691 ( .I1(\pred_tab[2][CODE_ADR][18] ), .I2(n23), .O(n620) );
  NAND_GATE U692 ( .I1(n622), .I2(n623), .O(n1629) );
  NAND_GATE U693 ( .I1(DI_adr[17]), .I2(n19), .O(n623) );
  NAND_GATE U694 ( .I1(\pred_tab[2][CODE_ADR][17] ), .I2(n23), .O(n622) );
  NAND_GATE U695 ( .I1(n624), .I2(n625), .O(n1630) );
  NAND_GATE U696 ( .I1(DI_adr[16]), .I2(n19), .O(n625) );
  NAND_GATE U697 ( .I1(\pred_tab[2][CODE_ADR][16] ), .I2(n23), .O(n624) );
  NAND_GATE U698 ( .I1(n626), .I2(n627), .O(n1631) );
  NAND_GATE U699 ( .I1(DI_adr[15]), .I2(n19), .O(n627) );
  NAND_GATE U700 ( .I1(\pred_tab[2][CODE_ADR][15] ), .I2(n23), .O(n626) );
  NAND_GATE U701 ( .I1(n628), .I2(n629), .O(n1632) );
  NAND_GATE U702 ( .I1(DI_adr[14]), .I2(n19), .O(n629) );
  NAND_GATE U703 ( .I1(\pred_tab[2][CODE_ADR][14] ), .I2(n23), .O(n628) );
  NAND_GATE U704 ( .I1(n630), .I2(n631), .O(n1633) );
  NAND_GATE U705 ( .I1(DI_adr[13]), .I2(n19), .O(n631) );
  NAND_GATE U706 ( .I1(\pred_tab[2][CODE_ADR][13] ), .I2(n23), .O(n630) );
  NAND_GATE U707 ( .I1(n632), .I2(n633), .O(n1634) );
  NAND_GATE U708 ( .I1(DI_adr[12]), .I2(n19), .O(n633) );
  NAND_GATE U709 ( .I1(\pred_tab[2][CODE_ADR][12] ), .I2(n23), .O(n632) );
  NAND_GATE U710 ( .I1(n634), .I2(n635), .O(n1635) );
  NAND_GATE U711 ( .I1(DI_adr[11]), .I2(n19), .O(n635) );
  NAND_GATE U712 ( .I1(\pred_tab[2][CODE_ADR][11] ), .I2(n23), .O(n634) );
  NAND_GATE U713 ( .I1(n636), .I2(n637), .O(n1636) );
  NAND_GATE U714 ( .I1(DI_adr[10]), .I2(n19), .O(n637) );
  NAND_GATE U715 ( .I1(\pred_tab[2][CODE_ADR][10] ), .I2(n23), .O(n636) );
  NAND_GATE U716 ( .I1(n638), .I2(n639), .O(n1637) );
  NAND_GATE U717 ( .I1(DI_adr[0]), .I2(n19), .O(n639) );
  NAND_GATE U718 ( .I1(\pred_tab[2][CODE_ADR][0] ), .I2(n23), .O(n638) );
  AND_GATE U720 ( .I1(n28), .I2(n434), .O(n163) );
  NAND_GATE U722 ( .I1(n640), .I2(n641), .O(n1640) );
  NAND_GATE U723 ( .I1(n646), .I2(n643), .O(n641) );
  NAND_GATE U724 ( .I1(n644), .I2(n645), .O(n643) );
  NAND_GATE U725 ( .I1(N1614), .I2(n13), .O(n645) );
  OR_GATE U726 ( .I1(n13), .I2(N1614), .O(n644) );
  NAND_GATE U727 ( .I1(\next_out[1] ), .I2(n647), .O(n640) );
  NAND_GATE U728 ( .I1(n648), .I2(n649), .O(n1641) );
  NAND_GATE U729 ( .I1(n646), .I2(n13), .O(n649) );
  NAND_GATE U731 ( .I1(\next_out[0] ), .I2(n647), .O(n648) );
  NAND4_GATE U732 ( .I1(n650), .I2(n651), .I3(n652), .I4(n653), .O(
        PR_bra_adr[9]) );
  AND4_GATE U733 ( .I1(n654), .I2(n655), .I3(n656), .I4(n657), .O(n653) );
  NAND_GATE U734 ( .I1(n658), .I2(n418), .O(n657) );
  NAND3_GATE U735 ( .I1(n659), .I2(n660), .I3(n661), .O(n418) );
  NAND_GATE U736 ( .I1(n662), .I2(N343), .O(n661) );
  NAND_GATE U737 ( .I1(\pred_tab[3][BRA_ADR][9] ), .I2(n663), .O(n660) );
  NAND_GATE U738 ( .I1(n664), .I2(EX_adresse[9]), .O(n659) );
  NAND_GATE U739 ( .I1(n665), .I2(n287), .O(n656) );
  NAND3_GATE U740 ( .I1(n666), .I2(n667), .I3(n668), .O(n287) );
  NAND_GATE U741 ( .I1(n669), .I2(N343), .O(n668) );
  NAND_GATE U742 ( .I1(\pred_tab[2][BRA_ADR][9] ), .I2(n670), .O(n667) );
  NAND_GATE U743 ( .I1(n671), .I2(EX_adresse[9]), .O(n666) );
  NAND_GATE U744 ( .I1(n672), .I2(n156), .O(n655) );
  NAND3_GATE U745 ( .I1(n673), .I2(n674), .I3(n675), .O(n156) );
  NAND_GATE U746 ( .I1(N343), .I2(n676), .O(n675) );
  NAND_GATE U747 ( .I1(\pred_tab[1][BRA_ADR][9] ), .I2(n677), .O(n674) );
  NAND_GATE U748 ( .I1(EX_adresse[9]), .I2(n678), .O(n673) );
  NAND_GATE U749 ( .I1(\pred_tab[1][BRA_ADR][9] ), .I2(n679), .O(n654) );
  NAND_GATE U750 ( .I1(N1253), .I2(n680), .O(n652) );
  NAND_GATE U751 ( .I1(\pred_tab[2][BRA_ADR][9] ), .I2(n681), .O(n651) );
  NAND_GATE U752 ( .I1(\pred_tab[3][BRA_ADR][9] ), .I2(n682), .O(n650) );
  NAND4_GATE U753 ( .I1(n683), .I2(n684), .I3(n685), .I4(n686), .O(
        PR_bra_adr[8]) );
  AND4_GATE U754 ( .I1(n687), .I2(n688), .I3(n689), .I4(n690), .O(n686) );
  NAND_GATE U755 ( .I1(n658), .I2(n414), .O(n690) );
  NAND3_GATE U756 ( .I1(n691), .I2(n692), .I3(n693), .O(n414) );
  NAND_GATE U757 ( .I1(n662), .I2(N342), .O(n693) );
  NAND_GATE U758 ( .I1(\pred_tab[3][BRA_ADR][8] ), .I2(n663), .O(n692) );
  NAND_GATE U759 ( .I1(n664), .I2(EX_adresse[8]), .O(n691) );
  NAND_GATE U760 ( .I1(n665), .I2(n283), .O(n689) );
  NAND3_GATE U761 ( .I1(n694), .I2(n695), .I3(n696), .O(n283) );
  NAND_GATE U762 ( .I1(n669), .I2(N342), .O(n696) );
  NAND_GATE U763 ( .I1(\pred_tab[2][BRA_ADR][8] ), .I2(n670), .O(n695) );
  NAND_GATE U764 ( .I1(n671), .I2(EX_adresse[8]), .O(n694) );
  NAND_GATE U765 ( .I1(n672), .I2(n152), .O(n688) );
  NAND3_GATE U766 ( .I1(n697), .I2(n698), .I3(n699), .O(n152) );
  NAND_GATE U767 ( .I1(N342), .I2(n676), .O(n699) );
  NAND_GATE U768 ( .I1(\pred_tab[1][BRA_ADR][8] ), .I2(n677), .O(n698) );
  NAND_GATE U769 ( .I1(EX_adresse[8]), .I2(n678), .O(n697) );
  NAND_GATE U770 ( .I1(\pred_tab[1][BRA_ADR][8] ), .I2(n679), .O(n687) );
  NAND_GATE U771 ( .I1(N1252), .I2(n680), .O(n685) );
  NAND_GATE U772 ( .I1(\pred_tab[2][BRA_ADR][8] ), .I2(n681), .O(n684) );
  NAND_GATE U773 ( .I1(\pred_tab[3][BRA_ADR][8] ), .I2(n682), .O(n683) );
  NAND4_GATE U774 ( .I1(n700), .I2(n701), .I3(n702), .I4(n703), .O(
        PR_bra_adr[7]) );
  AND4_GATE U775 ( .I1(n704), .I2(n705), .I3(n706), .I4(n707), .O(n703) );
  NAND_GATE U776 ( .I1(n658), .I2(n410), .O(n707) );
  NAND3_GATE U777 ( .I1(n708), .I2(n709), .I3(n710), .O(n410) );
  NAND_GATE U778 ( .I1(n662), .I2(N341), .O(n710) );
  NAND_GATE U779 ( .I1(\pred_tab[3][BRA_ADR][7] ), .I2(n663), .O(n709) );
  NAND_GATE U780 ( .I1(n664), .I2(EX_adresse[7]), .O(n708) );
  NAND_GATE U781 ( .I1(n665), .I2(n279), .O(n706) );
  NAND3_GATE U782 ( .I1(n711), .I2(n712), .I3(n713), .O(n279) );
  NAND_GATE U783 ( .I1(n669), .I2(N341), .O(n713) );
  NAND_GATE U784 ( .I1(\pred_tab[2][BRA_ADR][7] ), .I2(n670), .O(n712) );
  NAND_GATE U785 ( .I1(n671), .I2(EX_adresse[7]), .O(n711) );
  NAND_GATE U786 ( .I1(n672), .I2(n148), .O(n705) );
  NAND3_GATE U787 ( .I1(n714), .I2(n715), .I3(n716), .O(n148) );
  NAND_GATE U788 ( .I1(N341), .I2(n676), .O(n716) );
  NAND_GATE U789 ( .I1(\pred_tab[1][BRA_ADR][7] ), .I2(n677), .O(n715) );
  NAND_GATE U790 ( .I1(EX_adresse[7]), .I2(n678), .O(n714) );
  NAND_GATE U791 ( .I1(\pred_tab[1][BRA_ADR][7] ), .I2(n679), .O(n704) );
  NAND_GATE U792 ( .I1(N1251), .I2(n680), .O(n702) );
  NAND_GATE U793 ( .I1(\pred_tab[2][BRA_ADR][7] ), .I2(n681), .O(n701) );
  NAND_GATE U794 ( .I1(\pred_tab[3][BRA_ADR][7] ), .I2(n682), .O(n700) );
  NAND4_GATE U795 ( .I1(n717), .I2(n718), .I3(n719), .I4(n720), .O(
        PR_bra_adr[6]) );
  AND4_GATE U796 ( .I1(n721), .I2(n722), .I3(n723), .I4(n724), .O(n720) );
  NAND_GATE U797 ( .I1(n658), .I2(n406), .O(n724) );
  NAND3_GATE U798 ( .I1(n725), .I2(n726), .I3(n727), .O(n406) );
  NAND_GATE U799 ( .I1(n662), .I2(N340), .O(n727) );
  NAND_GATE U800 ( .I1(\pred_tab[3][BRA_ADR][6] ), .I2(n663), .O(n726) );
  NAND_GATE U801 ( .I1(n664), .I2(EX_adresse[6]), .O(n725) );
  NAND_GATE U802 ( .I1(n665), .I2(n275), .O(n723) );
  NAND3_GATE U803 ( .I1(n728), .I2(n729), .I3(n730), .O(n275) );
  NAND_GATE U804 ( .I1(n669), .I2(N340), .O(n730) );
  NAND_GATE U805 ( .I1(\pred_tab[2][BRA_ADR][6] ), .I2(n670), .O(n729) );
  NAND_GATE U806 ( .I1(n671), .I2(EX_adresse[6]), .O(n728) );
  NAND_GATE U807 ( .I1(n672), .I2(n144), .O(n722) );
  NAND3_GATE U808 ( .I1(n731), .I2(n732), .I3(n733), .O(n144) );
  NAND_GATE U809 ( .I1(N340), .I2(n676), .O(n733) );
  NAND_GATE U810 ( .I1(\pred_tab[1][BRA_ADR][6] ), .I2(n677), .O(n732) );
  NAND_GATE U811 ( .I1(EX_adresse[6]), .I2(n678), .O(n731) );
  NAND_GATE U812 ( .I1(\pred_tab[1][BRA_ADR][6] ), .I2(n679), .O(n721) );
  NAND_GATE U813 ( .I1(N1250), .I2(n680), .O(n719) );
  NAND_GATE U814 ( .I1(\pred_tab[2][BRA_ADR][6] ), .I2(n681), .O(n718) );
  NAND_GATE U815 ( .I1(\pred_tab[3][BRA_ADR][6] ), .I2(n682), .O(n717) );
  NAND4_GATE U816 ( .I1(n734), .I2(n735), .I3(n736), .I4(n737), .O(
        PR_bra_adr[5]) );
  AND4_GATE U817 ( .I1(n738), .I2(n739), .I3(n740), .I4(n741), .O(n737) );
  NAND_GATE U818 ( .I1(n658), .I2(n402), .O(n741) );
  NAND3_GATE U819 ( .I1(n742), .I2(n743), .I3(n744), .O(n402) );
  NAND_GATE U820 ( .I1(n662), .I2(N339), .O(n744) );
  NAND_GATE U821 ( .I1(\pred_tab[3][BRA_ADR][5] ), .I2(n663), .O(n743) );
  NAND_GATE U822 ( .I1(n664), .I2(EX_adresse[5]), .O(n742) );
  NAND_GATE U823 ( .I1(n665), .I2(n271), .O(n740) );
  NAND3_GATE U824 ( .I1(n745), .I2(n746), .I3(n747), .O(n271) );
  NAND_GATE U825 ( .I1(n669), .I2(N339), .O(n747) );
  NAND_GATE U826 ( .I1(\pred_tab[2][BRA_ADR][5] ), .I2(n670), .O(n746) );
  NAND_GATE U827 ( .I1(n671), .I2(EX_adresse[5]), .O(n745) );
  NAND_GATE U828 ( .I1(n672), .I2(n140), .O(n739) );
  NAND3_GATE U829 ( .I1(n748), .I2(n749), .I3(n750), .O(n140) );
  NAND_GATE U830 ( .I1(N339), .I2(n676), .O(n750) );
  NAND_GATE U831 ( .I1(\pred_tab[1][BRA_ADR][5] ), .I2(n677), .O(n749) );
  NAND_GATE U832 ( .I1(EX_adresse[5]), .I2(n678), .O(n748) );
  NAND_GATE U833 ( .I1(\pred_tab[1][BRA_ADR][5] ), .I2(n679), .O(n738) );
  NAND_GATE U834 ( .I1(N1249), .I2(n680), .O(n736) );
  NAND_GATE U835 ( .I1(\pred_tab[2][BRA_ADR][5] ), .I2(n681), .O(n735) );
  NAND_GATE U836 ( .I1(\pred_tab[3][BRA_ADR][5] ), .I2(n682), .O(n734) );
  NAND4_GATE U837 ( .I1(n751), .I2(n752), .I3(n753), .I4(n754), .O(
        PR_bra_adr[4]) );
  AND4_GATE U838 ( .I1(n755), .I2(n756), .I3(n757), .I4(n758), .O(n754) );
  NAND_GATE U839 ( .I1(n658), .I2(n398), .O(n758) );
  NAND3_GATE U840 ( .I1(n759), .I2(n760), .I3(n761), .O(n398) );
  NAND_GATE U841 ( .I1(n662), .I2(N338), .O(n761) );
  NAND_GATE U842 ( .I1(\pred_tab[3][BRA_ADR][4] ), .I2(n663), .O(n760) );
  NAND_GATE U843 ( .I1(n664), .I2(EX_adresse[4]), .O(n759) );
  NAND_GATE U844 ( .I1(n665), .I2(n267), .O(n757) );
  NAND3_GATE U845 ( .I1(n762), .I2(n763), .I3(n764), .O(n267) );
  NAND_GATE U846 ( .I1(n669), .I2(N338), .O(n764) );
  NAND_GATE U847 ( .I1(\pred_tab[2][BRA_ADR][4] ), .I2(n670), .O(n763) );
  NAND_GATE U848 ( .I1(n671), .I2(EX_adresse[4]), .O(n762) );
  NAND_GATE U849 ( .I1(n672), .I2(n136), .O(n756) );
  NAND3_GATE U850 ( .I1(n765), .I2(n766), .I3(n767), .O(n136) );
  NAND_GATE U851 ( .I1(N338), .I2(n676), .O(n767) );
  NAND_GATE U852 ( .I1(\pred_tab[1][BRA_ADR][4] ), .I2(n677), .O(n766) );
  NAND_GATE U853 ( .I1(EX_adresse[4]), .I2(n678), .O(n765) );
  NAND_GATE U854 ( .I1(\pred_tab[1][BRA_ADR][4] ), .I2(n679), .O(n755) );
  NAND_GATE U855 ( .I1(N1248), .I2(n680), .O(n753) );
  NAND_GATE U856 ( .I1(\pred_tab[2][BRA_ADR][4] ), .I2(n681), .O(n752) );
  NAND_GATE U857 ( .I1(\pred_tab[3][BRA_ADR][4] ), .I2(n682), .O(n751) );
  NAND4_GATE U858 ( .I1(n768), .I2(n769), .I3(n770), .I4(n771), .O(
        PR_bra_adr[3]) );
  AND4_GATE U859 ( .I1(n772), .I2(n773), .I3(n774), .I4(n775), .O(n771) );
  NAND_GATE U860 ( .I1(n658), .I2(n394), .O(n775) );
  NAND3_GATE U861 ( .I1(n776), .I2(n777), .I3(n778), .O(n394) );
  NAND_GATE U862 ( .I1(n662), .I2(N337), .O(n778) );
  NAND_GATE U863 ( .I1(\pred_tab[3][BRA_ADR][3] ), .I2(n663), .O(n777) );
  NAND_GATE U864 ( .I1(n664), .I2(EX_adresse[3]), .O(n776) );
  NAND_GATE U865 ( .I1(n665), .I2(n263), .O(n774) );
  NAND3_GATE U866 ( .I1(n779), .I2(n780), .I3(n781), .O(n263) );
  NAND_GATE U867 ( .I1(n669), .I2(N337), .O(n781) );
  NAND_GATE U868 ( .I1(\pred_tab[2][BRA_ADR][3] ), .I2(n670), .O(n780) );
  NAND_GATE U869 ( .I1(n671), .I2(EX_adresse[3]), .O(n779) );
  NAND_GATE U870 ( .I1(n672), .I2(n132), .O(n773) );
  NAND3_GATE U871 ( .I1(n782), .I2(n783), .I3(n784), .O(n132) );
  NAND_GATE U872 ( .I1(N337), .I2(n676), .O(n784) );
  NAND_GATE U873 ( .I1(\pred_tab[1][BRA_ADR][3] ), .I2(n677), .O(n783) );
  NAND_GATE U874 ( .I1(EX_adresse[3]), .I2(n678), .O(n782) );
  NAND_GATE U875 ( .I1(\pred_tab[1][BRA_ADR][3] ), .I2(n679), .O(n772) );
  NAND_GATE U876 ( .I1(N1247), .I2(n680), .O(n770) );
  NAND_GATE U877 ( .I1(\pred_tab[2][BRA_ADR][3] ), .I2(n681), .O(n769) );
  NAND_GATE U878 ( .I1(\pred_tab[3][BRA_ADR][3] ), .I2(n682), .O(n768) );
  NAND4_GATE U879 ( .I1(n785), .I2(n786), .I3(n787), .I4(n788), .O(
        PR_bra_adr[31]) );
  AND4_GATE U880 ( .I1(n789), .I2(n790), .I3(n791), .I4(n792), .O(n788) );
  NAND_GATE U881 ( .I1(n658), .I2(n390), .O(n792) );
  NAND3_GATE U882 ( .I1(n793), .I2(n794), .I3(n795), .O(n390) );
  NAND_GATE U883 ( .I1(n662), .I2(N365), .O(n795) );
  NAND_GATE U884 ( .I1(\pred_tab[3][BRA_ADR][31] ), .I2(n663), .O(n794) );
  NAND_GATE U885 ( .I1(n664), .I2(EX_adresse[31]), .O(n793) );
  NAND_GATE U886 ( .I1(n665), .I2(n259), .O(n791) );
  NAND3_GATE U887 ( .I1(n796), .I2(n797), .I3(n798), .O(n259) );
  NAND_GATE U888 ( .I1(n669), .I2(N365), .O(n798) );
  NAND_GATE U889 ( .I1(\pred_tab[2][BRA_ADR][31] ), .I2(n670), .O(n797) );
  NAND_GATE U890 ( .I1(n671), .I2(EX_adresse[31]), .O(n796) );
  NAND_GATE U891 ( .I1(n672), .I2(n128), .O(n790) );
  NAND3_GATE U892 ( .I1(n799), .I2(n800), .I3(n801), .O(n128) );
  NAND_GATE U893 ( .I1(N365), .I2(n676), .O(n801) );
  NAND_GATE U894 ( .I1(\pred_tab[1][BRA_ADR][31] ), .I2(n677), .O(n800) );
  NAND_GATE U895 ( .I1(EX_adresse[31]), .I2(n678), .O(n799) );
  NAND_GATE U896 ( .I1(\pred_tab[1][BRA_ADR][31] ), .I2(n679), .O(n789) );
  NAND_GATE U897 ( .I1(N1275), .I2(n680), .O(n787) );
  NAND_GATE U898 ( .I1(\pred_tab[2][BRA_ADR][31] ), .I2(n681), .O(n786) );
  NAND_GATE U899 ( .I1(\pred_tab[3][BRA_ADR][31] ), .I2(n682), .O(n785) );
  NAND4_GATE U900 ( .I1(n802), .I2(n803), .I3(n804), .I4(n805), .O(
        PR_bra_adr[30]) );
  AND4_GATE U901 ( .I1(n806), .I2(n807), .I3(n808), .I4(n809), .O(n805) );
  NAND_GATE U902 ( .I1(n658), .I2(n386), .O(n809) );
  NAND3_GATE U903 ( .I1(n810), .I2(n811), .I3(n812), .O(n386) );
  NAND_GATE U904 ( .I1(n662), .I2(N364), .O(n812) );
  NAND_GATE U905 ( .I1(\pred_tab[3][BRA_ADR][30] ), .I2(n663), .O(n811) );
  NAND_GATE U906 ( .I1(n664), .I2(EX_adresse[30]), .O(n810) );
  NAND_GATE U907 ( .I1(n665), .I2(n255), .O(n808) );
  NAND3_GATE U908 ( .I1(n813), .I2(n814), .I3(n815), .O(n255) );
  NAND_GATE U909 ( .I1(n669), .I2(N364), .O(n815) );
  NAND_GATE U910 ( .I1(\pred_tab[2][BRA_ADR][30] ), .I2(n670), .O(n814) );
  NAND_GATE U911 ( .I1(n671), .I2(EX_adresse[30]), .O(n813) );
  NAND_GATE U912 ( .I1(n672), .I2(n124), .O(n807) );
  NAND3_GATE U913 ( .I1(n816), .I2(n817), .I3(n818), .O(n124) );
  NAND_GATE U914 ( .I1(N364), .I2(n676), .O(n818) );
  NAND_GATE U915 ( .I1(\pred_tab[1][BRA_ADR][30] ), .I2(n677), .O(n817) );
  NAND_GATE U916 ( .I1(EX_adresse[30]), .I2(n678), .O(n816) );
  NAND_GATE U917 ( .I1(\pred_tab[1][BRA_ADR][30] ), .I2(n679), .O(n806) );
  NAND_GATE U918 ( .I1(N1274), .I2(n680), .O(n804) );
  NAND_GATE U919 ( .I1(\pred_tab[2][BRA_ADR][30] ), .I2(n681), .O(n803) );
  NAND_GATE U920 ( .I1(\pred_tab[3][BRA_ADR][30] ), .I2(n682), .O(n802) );
  NAND4_GATE U921 ( .I1(n819), .I2(n820), .I3(n821), .I4(n822), .O(
        PR_bra_adr[2]) );
  AND4_GATE U922 ( .I1(n823), .I2(n824), .I3(n825), .I4(n826), .O(n822) );
  NAND_GATE U923 ( .I1(n658), .I2(n382), .O(n826) );
  NAND3_GATE U924 ( .I1(n827), .I2(n828), .I3(n829), .O(n382) );
  NAND_GATE U925 ( .I1(n662), .I2(N336), .O(n829) );
  NAND_GATE U926 ( .I1(\pred_tab[3][BRA_ADR][2] ), .I2(n663), .O(n828) );
  NAND_GATE U927 ( .I1(n664), .I2(EX_adresse[2]), .O(n827) );
  NAND_GATE U928 ( .I1(n665), .I2(n251), .O(n825) );
  NAND3_GATE U929 ( .I1(n830), .I2(n831), .I3(n832), .O(n251) );
  NAND_GATE U930 ( .I1(n669), .I2(N336), .O(n832) );
  NAND_GATE U931 ( .I1(\pred_tab[2][BRA_ADR][2] ), .I2(n670), .O(n831) );
  NAND_GATE U932 ( .I1(n671), .I2(EX_adresse[2]), .O(n830) );
  NAND_GATE U933 ( .I1(n672), .I2(n120), .O(n824) );
  NAND3_GATE U934 ( .I1(n833), .I2(n834), .I3(n835), .O(n120) );
  NAND_GATE U935 ( .I1(N336), .I2(n676), .O(n835) );
  NAND_GATE U936 ( .I1(\pred_tab[1][BRA_ADR][2] ), .I2(n677), .O(n834) );
  NAND_GATE U937 ( .I1(EX_adresse[2]), .I2(n678), .O(n833) );
  NAND_GATE U938 ( .I1(\pred_tab[1][BRA_ADR][2] ), .I2(n679), .O(n823) );
  NAND_GATE U939 ( .I1(N1246), .I2(n680), .O(n821) );
  NAND_GATE U940 ( .I1(\pred_tab[2][BRA_ADR][2] ), .I2(n681), .O(n820) );
  NAND_GATE U941 ( .I1(\pred_tab[3][BRA_ADR][2] ), .I2(n682), .O(n819) );
  NAND4_GATE U942 ( .I1(n836), .I2(n837), .I3(n838), .I4(n839), .O(
        PR_bra_adr[29]) );
  AND4_GATE U943 ( .I1(n840), .I2(n841), .I3(n842), .I4(n843), .O(n839) );
  NAND_GATE U944 ( .I1(n658), .I2(n378), .O(n843) );
  NAND3_GATE U945 ( .I1(n844), .I2(n845), .I3(n846), .O(n378) );
  NAND_GATE U946 ( .I1(n662), .I2(N363), .O(n846) );
  NAND_GATE U947 ( .I1(\pred_tab[3][BRA_ADR][29] ), .I2(n663), .O(n845) );
  NAND_GATE U948 ( .I1(n664), .I2(EX_adresse[29]), .O(n844) );
  NAND_GATE U949 ( .I1(n665), .I2(n247), .O(n842) );
  NAND3_GATE U950 ( .I1(n847), .I2(n848), .I3(n849), .O(n247) );
  NAND_GATE U951 ( .I1(n669), .I2(N363), .O(n849) );
  NAND_GATE U952 ( .I1(\pred_tab[2][BRA_ADR][29] ), .I2(n670), .O(n848) );
  NAND_GATE U953 ( .I1(n671), .I2(EX_adresse[29]), .O(n847) );
  NAND_GATE U954 ( .I1(n672), .I2(n116), .O(n841) );
  NAND3_GATE U955 ( .I1(n850), .I2(n851), .I3(n852), .O(n116) );
  NAND_GATE U956 ( .I1(N363), .I2(n676), .O(n852) );
  NAND_GATE U957 ( .I1(\pred_tab[1][BRA_ADR][29] ), .I2(n677), .O(n851) );
  NAND_GATE U958 ( .I1(EX_adresse[29]), .I2(n678), .O(n850) );
  NAND_GATE U959 ( .I1(\pred_tab[1][BRA_ADR][29] ), .I2(n679), .O(n840) );
  NAND_GATE U960 ( .I1(N1273), .I2(n680), .O(n838) );
  NAND_GATE U961 ( .I1(\pred_tab[2][BRA_ADR][29] ), .I2(n681), .O(n837) );
  NAND_GATE U962 ( .I1(\pred_tab[3][BRA_ADR][29] ), .I2(n682), .O(n836) );
  NAND4_GATE U963 ( .I1(n853), .I2(n854), .I3(n855), .I4(n856), .O(
        PR_bra_adr[28]) );
  AND4_GATE U964 ( .I1(n857), .I2(n858), .I3(n859), .I4(n860), .O(n856) );
  NAND_GATE U965 ( .I1(n658), .I2(n374), .O(n860) );
  NAND3_GATE U966 ( .I1(n861), .I2(n862), .I3(n863), .O(n374) );
  NAND_GATE U967 ( .I1(n662), .I2(N362), .O(n863) );
  NAND_GATE U968 ( .I1(\pred_tab[3][BRA_ADR][28] ), .I2(n663), .O(n862) );
  NAND_GATE U969 ( .I1(n664), .I2(EX_adresse[28]), .O(n861) );
  NAND_GATE U970 ( .I1(n665), .I2(n243), .O(n859) );
  NAND3_GATE U971 ( .I1(n864), .I2(n865), .I3(n866), .O(n243) );
  NAND_GATE U972 ( .I1(n669), .I2(N362), .O(n866) );
  NAND_GATE U973 ( .I1(\pred_tab[2][BRA_ADR][28] ), .I2(n670), .O(n865) );
  NAND_GATE U974 ( .I1(n671), .I2(EX_adresse[28]), .O(n864) );
  NAND_GATE U975 ( .I1(n672), .I2(n112), .O(n858) );
  NAND3_GATE U976 ( .I1(n867), .I2(n868), .I3(n869), .O(n112) );
  NAND_GATE U977 ( .I1(N362), .I2(n676), .O(n869) );
  NAND_GATE U978 ( .I1(\pred_tab[1][BRA_ADR][28] ), .I2(n677), .O(n868) );
  NAND_GATE U979 ( .I1(EX_adresse[28]), .I2(n678), .O(n867) );
  NAND_GATE U980 ( .I1(\pred_tab[1][BRA_ADR][28] ), .I2(n679), .O(n857) );
  NAND_GATE U981 ( .I1(N1272), .I2(n680), .O(n855) );
  NAND_GATE U982 ( .I1(\pred_tab[2][BRA_ADR][28] ), .I2(n681), .O(n854) );
  NAND_GATE U983 ( .I1(\pred_tab[3][BRA_ADR][28] ), .I2(n682), .O(n853) );
  NAND4_GATE U984 ( .I1(n870), .I2(n871), .I3(n872), .I4(n873), .O(
        PR_bra_adr[27]) );
  AND4_GATE U985 ( .I1(n874), .I2(n875), .I3(n876), .I4(n877), .O(n873) );
  NAND_GATE U986 ( .I1(n658), .I2(n370), .O(n877) );
  NAND3_GATE U987 ( .I1(n878), .I2(n879), .I3(n880), .O(n370) );
  NAND_GATE U988 ( .I1(n662), .I2(N361), .O(n880) );
  NAND_GATE U989 ( .I1(\pred_tab[3][BRA_ADR][27] ), .I2(n663), .O(n879) );
  NAND_GATE U990 ( .I1(n664), .I2(EX_adresse[27]), .O(n878) );
  NAND_GATE U991 ( .I1(n665), .I2(n239), .O(n876) );
  NAND3_GATE U992 ( .I1(n881), .I2(n882), .I3(n883), .O(n239) );
  NAND_GATE U993 ( .I1(n669), .I2(N361), .O(n883) );
  NAND_GATE U994 ( .I1(\pred_tab[2][BRA_ADR][27] ), .I2(n670), .O(n882) );
  NAND_GATE U995 ( .I1(n671), .I2(EX_adresse[27]), .O(n881) );
  NAND_GATE U996 ( .I1(n672), .I2(n108), .O(n875) );
  NAND3_GATE U997 ( .I1(n884), .I2(n885), .I3(n886), .O(n108) );
  NAND_GATE U998 ( .I1(N361), .I2(n676), .O(n886) );
  NAND_GATE U999 ( .I1(\pred_tab[1][BRA_ADR][27] ), .I2(n677), .O(n885) );
  NAND_GATE U1000 ( .I1(EX_adresse[27]), .I2(n678), .O(n884) );
  NAND_GATE U1001 ( .I1(\pred_tab[1][BRA_ADR][27] ), .I2(n679), .O(n874) );
  NAND_GATE U1002 ( .I1(N1271), .I2(n680), .O(n872) );
  NAND_GATE U1003 ( .I1(\pred_tab[2][BRA_ADR][27] ), .I2(n681), .O(n871) );
  NAND_GATE U1004 ( .I1(\pred_tab[3][BRA_ADR][27] ), .I2(n682), .O(n870) );
  NAND4_GATE U1005 ( .I1(n887), .I2(n888), .I3(n889), .I4(n890), .O(
        PR_bra_adr[26]) );
  AND4_GATE U1006 ( .I1(n891), .I2(n892), .I3(n893), .I4(n894), .O(n890) );
  NAND_GATE U1007 ( .I1(n658), .I2(n366), .O(n894) );
  NAND3_GATE U1008 ( .I1(n895), .I2(n896), .I3(n897), .O(n366) );
  NAND_GATE U1009 ( .I1(n662), .I2(N360), .O(n897) );
  NAND_GATE U1010 ( .I1(\pred_tab[3][BRA_ADR][26] ), .I2(n663), .O(n896) );
  NAND_GATE U1011 ( .I1(n664), .I2(EX_adresse[26]), .O(n895) );
  NAND_GATE U1012 ( .I1(n665), .I2(n235), .O(n893) );
  NAND3_GATE U1013 ( .I1(n898), .I2(n899), .I3(n900), .O(n235) );
  NAND_GATE U1014 ( .I1(n669), .I2(N360), .O(n900) );
  NAND_GATE U1015 ( .I1(\pred_tab[2][BRA_ADR][26] ), .I2(n670), .O(n899) );
  NAND_GATE U1016 ( .I1(n671), .I2(EX_adresse[26]), .O(n898) );
  NAND_GATE U1017 ( .I1(n672), .I2(n104), .O(n892) );
  NAND3_GATE U1018 ( .I1(n901), .I2(n902), .I3(n903), .O(n104) );
  NAND_GATE U1019 ( .I1(N360), .I2(n676), .O(n903) );
  NAND_GATE U1020 ( .I1(\pred_tab[1][BRA_ADR][26] ), .I2(n677), .O(n902) );
  NAND_GATE U1021 ( .I1(EX_adresse[26]), .I2(n678), .O(n901) );
  NAND_GATE U1022 ( .I1(\pred_tab[1][BRA_ADR][26] ), .I2(n679), .O(n891) );
  NAND_GATE U1023 ( .I1(N1270), .I2(n680), .O(n889) );
  NAND_GATE U1024 ( .I1(\pred_tab[2][BRA_ADR][26] ), .I2(n681), .O(n888) );
  NAND_GATE U1025 ( .I1(\pred_tab[3][BRA_ADR][26] ), .I2(n682), .O(n887) );
  NAND4_GATE U1026 ( .I1(n904), .I2(n905), .I3(n906), .I4(n907), .O(
        PR_bra_adr[25]) );
  AND4_GATE U1027 ( .I1(n908), .I2(n909), .I3(n910), .I4(n911), .O(n907) );
  NAND_GATE U1028 ( .I1(n658), .I2(n362), .O(n911) );
  NAND3_GATE U1029 ( .I1(n912), .I2(n913), .I3(n914), .O(n362) );
  NAND_GATE U1030 ( .I1(n662), .I2(N359), .O(n914) );
  NAND_GATE U1031 ( .I1(\pred_tab[3][BRA_ADR][25] ), .I2(n663), .O(n913) );
  NAND_GATE U1032 ( .I1(n664), .I2(EX_adresse[25]), .O(n912) );
  NAND_GATE U1033 ( .I1(n665), .I2(n231), .O(n910) );
  NAND3_GATE U1034 ( .I1(n915), .I2(n916), .I3(n917), .O(n231) );
  NAND_GATE U1035 ( .I1(n669), .I2(N359), .O(n917) );
  NAND_GATE U1036 ( .I1(\pred_tab[2][BRA_ADR][25] ), .I2(n670), .O(n916) );
  NAND_GATE U1037 ( .I1(n671), .I2(EX_adresse[25]), .O(n915) );
  NAND_GATE U1038 ( .I1(n672), .I2(n100), .O(n909) );
  NAND3_GATE U1039 ( .I1(n918), .I2(n919), .I3(n920), .O(n100) );
  NAND_GATE U1040 ( .I1(N359), .I2(n676), .O(n920) );
  NAND_GATE U1041 ( .I1(\pred_tab[1][BRA_ADR][25] ), .I2(n677), .O(n919) );
  NAND_GATE U1042 ( .I1(EX_adresse[25]), .I2(n678), .O(n918) );
  NAND_GATE U1043 ( .I1(\pred_tab[1][BRA_ADR][25] ), .I2(n679), .O(n908) );
  NAND_GATE U1044 ( .I1(N1269), .I2(n680), .O(n906) );
  NAND_GATE U1045 ( .I1(\pred_tab[2][BRA_ADR][25] ), .I2(n681), .O(n905) );
  NAND_GATE U1046 ( .I1(\pred_tab[3][BRA_ADR][25] ), .I2(n682), .O(n904) );
  NAND4_GATE U1047 ( .I1(n921), .I2(n922), .I3(n923), .I4(n924), .O(
        PR_bra_adr[24]) );
  AND4_GATE U1048 ( .I1(n925), .I2(n926), .I3(n927), .I4(n928), .O(n924) );
  NAND_GATE U1049 ( .I1(n658), .I2(n358), .O(n928) );
  NAND3_GATE U1050 ( .I1(n929), .I2(n930), .I3(n931), .O(n358) );
  NAND_GATE U1051 ( .I1(n662), .I2(N358), .O(n931) );
  NAND_GATE U1052 ( .I1(\pred_tab[3][BRA_ADR][24] ), .I2(n663), .O(n930) );
  NAND_GATE U1053 ( .I1(n664), .I2(EX_adresse[24]), .O(n929) );
  NAND_GATE U1054 ( .I1(n665), .I2(n227), .O(n927) );
  NAND3_GATE U1055 ( .I1(n932), .I2(n933), .I3(n934), .O(n227) );
  NAND_GATE U1056 ( .I1(n669), .I2(N358), .O(n934) );
  NAND_GATE U1057 ( .I1(\pred_tab[2][BRA_ADR][24] ), .I2(n670), .O(n933) );
  NAND_GATE U1058 ( .I1(n671), .I2(EX_adresse[24]), .O(n932) );
  NAND_GATE U1059 ( .I1(n672), .I2(n96), .O(n926) );
  NAND3_GATE U1060 ( .I1(n935), .I2(n936), .I3(n937), .O(n96) );
  NAND_GATE U1061 ( .I1(N358), .I2(n676), .O(n937) );
  NAND_GATE U1062 ( .I1(\pred_tab[1][BRA_ADR][24] ), .I2(n677), .O(n936) );
  NAND_GATE U1063 ( .I1(EX_adresse[24]), .I2(n678), .O(n935) );
  NAND_GATE U1064 ( .I1(\pred_tab[1][BRA_ADR][24] ), .I2(n679), .O(n925) );
  NAND_GATE U1065 ( .I1(N1268), .I2(n680), .O(n923) );
  NAND_GATE U1066 ( .I1(\pred_tab[2][BRA_ADR][24] ), .I2(n681), .O(n922) );
  NAND_GATE U1067 ( .I1(\pred_tab[3][BRA_ADR][24] ), .I2(n682), .O(n921) );
  NAND4_GATE U1068 ( .I1(n938), .I2(n939), .I3(n940), .I4(n941), .O(
        PR_bra_adr[23]) );
  AND4_GATE U1069 ( .I1(n942), .I2(n943), .I3(n944), .I4(n945), .O(n941) );
  NAND_GATE U1070 ( .I1(n658), .I2(n354), .O(n945) );
  NAND3_GATE U1071 ( .I1(n946), .I2(n947), .I3(n948), .O(n354) );
  NAND_GATE U1072 ( .I1(n662), .I2(N357), .O(n948) );
  NAND_GATE U1073 ( .I1(\pred_tab[3][BRA_ADR][23] ), .I2(n663), .O(n947) );
  NAND_GATE U1074 ( .I1(n664), .I2(EX_adresse[23]), .O(n946) );
  NAND_GATE U1075 ( .I1(n665), .I2(n223), .O(n944) );
  NAND3_GATE U1076 ( .I1(n949), .I2(n950), .I3(n951), .O(n223) );
  NAND_GATE U1077 ( .I1(n669), .I2(N357), .O(n951) );
  NAND_GATE U1078 ( .I1(\pred_tab[2][BRA_ADR][23] ), .I2(n670), .O(n950) );
  NAND_GATE U1079 ( .I1(n671), .I2(EX_adresse[23]), .O(n949) );
  NAND_GATE U1080 ( .I1(n672), .I2(n92), .O(n943) );
  NAND3_GATE U1081 ( .I1(n952), .I2(n953), .I3(n954), .O(n92) );
  NAND_GATE U1082 ( .I1(N357), .I2(n676), .O(n954) );
  NAND_GATE U1083 ( .I1(\pred_tab[1][BRA_ADR][23] ), .I2(n677), .O(n953) );
  NAND_GATE U1084 ( .I1(EX_adresse[23]), .I2(n678), .O(n952) );
  NAND_GATE U1085 ( .I1(\pred_tab[1][BRA_ADR][23] ), .I2(n679), .O(n942) );
  NAND_GATE U1086 ( .I1(N1267), .I2(n680), .O(n940) );
  NAND_GATE U1087 ( .I1(\pred_tab[2][BRA_ADR][23] ), .I2(n681), .O(n939) );
  NAND_GATE U1088 ( .I1(\pred_tab[3][BRA_ADR][23] ), .I2(n682), .O(n938) );
  NAND4_GATE U1089 ( .I1(n955), .I2(n956), .I3(n957), .I4(n958), .O(
        PR_bra_adr[22]) );
  AND4_GATE U1090 ( .I1(n959), .I2(n960), .I3(n961), .I4(n962), .O(n958) );
  NAND_GATE U1091 ( .I1(n658), .I2(n350), .O(n962) );
  NAND3_GATE U1092 ( .I1(n963), .I2(n964), .I3(n965), .O(n350) );
  NAND_GATE U1093 ( .I1(n662), .I2(N356), .O(n965) );
  NAND_GATE U1094 ( .I1(\pred_tab[3][BRA_ADR][22] ), .I2(n663), .O(n964) );
  NAND_GATE U1095 ( .I1(n664), .I2(EX_adresse[22]), .O(n963) );
  NAND_GATE U1096 ( .I1(n665), .I2(n219), .O(n961) );
  NAND3_GATE U1097 ( .I1(n966), .I2(n967), .I3(n968), .O(n219) );
  NAND_GATE U1098 ( .I1(n669), .I2(N356), .O(n968) );
  NAND_GATE U1099 ( .I1(\pred_tab[2][BRA_ADR][22] ), .I2(n670), .O(n967) );
  NAND_GATE U1100 ( .I1(n671), .I2(EX_adresse[22]), .O(n966) );
  NAND_GATE U1101 ( .I1(n672), .I2(n88), .O(n960) );
  NAND3_GATE U1102 ( .I1(n969), .I2(n970), .I3(n971), .O(n88) );
  NAND_GATE U1103 ( .I1(N356), .I2(n676), .O(n971) );
  NAND_GATE U1104 ( .I1(\pred_tab[1][BRA_ADR][22] ), .I2(n677), .O(n970) );
  NAND_GATE U1105 ( .I1(EX_adresse[22]), .I2(n678), .O(n969) );
  NAND_GATE U1106 ( .I1(\pred_tab[1][BRA_ADR][22] ), .I2(n679), .O(n959) );
  NAND_GATE U1107 ( .I1(N1266), .I2(n680), .O(n957) );
  NAND_GATE U1108 ( .I1(\pred_tab[2][BRA_ADR][22] ), .I2(n681), .O(n956) );
  NAND_GATE U1109 ( .I1(\pred_tab[3][BRA_ADR][22] ), .I2(n682), .O(n955) );
  NAND4_GATE U1110 ( .I1(n972), .I2(n973), .I3(n974), .I4(n975), .O(
        PR_bra_adr[21]) );
  AND4_GATE U1111 ( .I1(n976), .I2(n977), .I3(n978), .I4(n979), .O(n975) );
  NAND_GATE U1112 ( .I1(n658), .I2(n346), .O(n979) );
  NAND3_GATE U1113 ( .I1(n980), .I2(n981), .I3(n982), .O(n346) );
  NAND_GATE U1114 ( .I1(n662), .I2(N355), .O(n982) );
  NAND_GATE U1115 ( .I1(\pred_tab[3][BRA_ADR][21] ), .I2(n663), .O(n981) );
  NAND_GATE U1116 ( .I1(n664), .I2(EX_adresse[21]), .O(n980) );
  NAND_GATE U1117 ( .I1(n665), .I2(n215), .O(n978) );
  NAND3_GATE U1118 ( .I1(n983), .I2(n984), .I3(n985), .O(n215) );
  NAND_GATE U1119 ( .I1(n669), .I2(N355), .O(n985) );
  NAND_GATE U1120 ( .I1(\pred_tab[2][BRA_ADR][21] ), .I2(n670), .O(n984) );
  NAND_GATE U1121 ( .I1(n671), .I2(EX_adresse[21]), .O(n983) );
  NAND_GATE U1122 ( .I1(n672), .I2(n84), .O(n977) );
  NAND3_GATE U1123 ( .I1(n986), .I2(n987), .I3(n988), .O(n84) );
  NAND_GATE U1124 ( .I1(N355), .I2(n676), .O(n988) );
  NAND_GATE U1125 ( .I1(\pred_tab[1][BRA_ADR][21] ), .I2(n677), .O(n987) );
  NAND_GATE U1126 ( .I1(EX_adresse[21]), .I2(n678), .O(n986) );
  NAND_GATE U1127 ( .I1(\pred_tab[1][BRA_ADR][21] ), .I2(n679), .O(n976) );
  NAND_GATE U1128 ( .I1(N1265), .I2(n680), .O(n974) );
  NAND_GATE U1129 ( .I1(\pred_tab[2][BRA_ADR][21] ), .I2(n681), .O(n973) );
  NAND_GATE U1130 ( .I1(\pred_tab[3][BRA_ADR][21] ), .I2(n682), .O(n972) );
  NAND4_GATE U1131 ( .I1(n989), .I2(n990), .I3(n991), .I4(n992), .O(
        PR_bra_adr[20]) );
  AND4_GATE U1132 ( .I1(n993), .I2(n994), .I3(n995), .I4(n996), .O(n992) );
  NAND_GATE U1133 ( .I1(n658), .I2(n342), .O(n996) );
  NAND3_GATE U1134 ( .I1(n997), .I2(n998), .I3(n999), .O(n342) );
  NAND_GATE U1135 ( .I1(n662), .I2(N354), .O(n999) );
  NAND_GATE U1136 ( .I1(\pred_tab[3][BRA_ADR][20] ), .I2(n663), .O(n998) );
  NAND_GATE U1137 ( .I1(n664), .I2(EX_adresse[20]), .O(n997) );
  NAND_GATE U1138 ( .I1(n665), .I2(n211), .O(n995) );
  NAND3_GATE U1139 ( .I1(n1000), .I2(n1001), .I3(n1002), .O(n211) );
  NAND_GATE U1140 ( .I1(n669), .I2(N354), .O(n1002) );
  NAND_GATE U1141 ( .I1(\pred_tab[2][BRA_ADR][20] ), .I2(n670), .O(n1001) );
  NAND_GATE U1142 ( .I1(n671), .I2(EX_adresse[20]), .O(n1000) );
  NAND_GATE U1143 ( .I1(n672), .I2(n80), .O(n994) );
  NAND3_GATE U1144 ( .I1(n1003), .I2(n1004), .I3(n1005), .O(n80) );
  NAND_GATE U1145 ( .I1(N354), .I2(n676), .O(n1005) );
  NAND_GATE U1146 ( .I1(\pred_tab[1][BRA_ADR][20] ), .I2(n677), .O(n1004) );
  NAND_GATE U1147 ( .I1(EX_adresse[20]), .I2(n678), .O(n1003) );
  NAND_GATE U1148 ( .I1(\pred_tab[1][BRA_ADR][20] ), .I2(n679), .O(n993) );
  NAND_GATE U1149 ( .I1(N1264), .I2(n680), .O(n991) );
  NAND_GATE U1150 ( .I1(\pred_tab[2][BRA_ADR][20] ), .I2(n681), .O(n990) );
  NAND_GATE U1151 ( .I1(\pred_tab[3][BRA_ADR][20] ), .I2(n682), .O(n989) );
  NAND4_GATE U1152 ( .I1(n1006), .I2(n1007), .I3(n1008), .I4(n1009), .O(
        PR_bra_adr[1]) );
  AND4_GATE U1153 ( .I1(n1010), .I2(n1011), .I3(n1012), .I4(n1013), .O(n1009)
         );
  NAND_GATE U1154 ( .I1(n658), .I2(n338), .O(n1013) );
  NAND3_GATE U1155 ( .I1(n1014), .I2(n1015), .I3(n1016), .O(n338) );
  NAND_GATE U1156 ( .I1(n662), .I2(N335), .O(n1016) );
  NAND_GATE U1157 ( .I1(\pred_tab[3][BRA_ADR][1] ), .I2(n663), .O(n1015) );
  NAND_GATE U1158 ( .I1(n664), .I2(EX_adresse[1]), .O(n1014) );
  NAND_GATE U1159 ( .I1(n665), .I2(n207), .O(n1012) );
  NAND3_GATE U1160 ( .I1(n1017), .I2(n1018), .I3(n1019), .O(n207) );
  NAND_GATE U1161 ( .I1(n669), .I2(N335), .O(n1019) );
  NAND_GATE U1162 ( .I1(\pred_tab[2][BRA_ADR][1] ), .I2(n670), .O(n1018) );
  NAND_GATE U1163 ( .I1(n671), .I2(EX_adresse[1]), .O(n1017) );
  NAND_GATE U1164 ( .I1(n672), .I2(n76), .O(n1011) );
  NAND3_GATE U1165 ( .I1(n1020), .I2(n1021), .I3(n1022), .O(n76) );
  NAND_GATE U1166 ( .I1(N335), .I2(n676), .O(n1022) );
  NAND_GATE U1167 ( .I1(\pred_tab[1][BRA_ADR][1] ), .I2(n677), .O(n1021) );
  NAND_GATE U1168 ( .I1(EX_adresse[1]), .I2(n678), .O(n1020) );
  NAND_GATE U1169 ( .I1(\pred_tab[1][BRA_ADR][1] ), .I2(n679), .O(n1010) );
  NAND_GATE U1170 ( .I1(N1245), .I2(n680), .O(n1008) );
  NAND_GATE U1171 ( .I1(\pred_tab[2][BRA_ADR][1] ), .I2(n681), .O(n1007) );
  NAND_GATE U1172 ( .I1(\pred_tab[3][BRA_ADR][1] ), .I2(n682), .O(n1006) );
  NAND4_GATE U1173 ( .I1(n1023), .I2(n1024), .I3(n1025), .I4(n1026), .O(
        PR_bra_adr[19]) );
  AND4_GATE U1174 ( .I1(n1027), .I2(n1028), .I3(n1029), .I4(n1030), .O(n1026)
         );
  NAND_GATE U1175 ( .I1(n658), .I2(n334), .O(n1030) );
  NAND3_GATE U1176 ( .I1(n1031), .I2(n1032), .I3(n1033), .O(n334) );
  NAND_GATE U1177 ( .I1(n662), .I2(N353), .O(n1033) );
  NAND_GATE U1178 ( .I1(\pred_tab[3][BRA_ADR][19] ), .I2(n663), .O(n1032) );
  NAND_GATE U1179 ( .I1(n664), .I2(EX_adresse[19]), .O(n1031) );
  NAND_GATE U1180 ( .I1(n665), .I2(n203), .O(n1029) );
  NAND3_GATE U1181 ( .I1(n1034), .I2(n1035), .I3(n1036), .O(n203) );
  NAND_GATE U1182 ( .I1(n669), .I2(N353), .O(n1036) );
  NAND_GATE U1183 ( .I1(\pred_tab[2][BRA_ADR][19] ), .I2(n670), .O(n1035) );
  NAND_GATE U1184 ( .I1(n671), .I2(EX_adresse[19]), .O(n1034) );
  NAND_GATE U1185 ( .I1(n672), .I2(n72), .O(n1028) );
  NAND3_GATE U1186 ( .I1(n1037), .I2(n1038), .I3(n1039), .O(n72) );
  NAND_GATE U1187 ( .I1(N353), .I2(n676), .O(n1039) );
  NAND_GATE U1188 ( .I1(\pred_tab[1][BRA_ADR][19] ), .I2(n677), .O(n1038) );
  NAND_GATE U1189 ( .I1(EX_adresse[19]), .I2(n678), .O(n1037) );
  NAND_GATE U1190 ( .I1(\pred_tab[1][BRA_ADR][19] ), .I2(n679), .O(n1027) );
  NAND_GATE U1191 ( .I1(N1263), .I2(n680), .O(n1025) );
  NAND_GATE U1192 ( .I1(\pred_tab[2][BRA_ADR][19] ), .I2(n681), .O(n1024) );
  NAND_GATE U1193 ( .I1(\pred_tab[3][BRA_ADR][19] ), .I2(n682), .O(n1023) );
  NAND4_GATE U1194 ( .I1(n1040), .I2(n1041), .I3(n1042), .I4(n1043), .O(
        PR_bra_adr[18]) );
  AND4_GATE U1195 ( .I1(n1044), .I2(n1045), .I3(n1046), .I4(n1047), .O(n1043)
         );
  NAND_GATE U1196 ( .I1(n658), .I2(n330), .O(n1047) );
  NAND3_GATE U1197 ( .I1(n1048), .I2(n1049), .I3(n1050), .O(n330) );
  NAND_GATE U1198 ( .I1(n662), .I2(N352), .O(n1050) );
  NAND_GATE U1199 ( .I1(\pred_tab[3][BRA_ADR][18] ), .I2(n663), .O(n1049) );
  NAND_GATE U1200 ( .I1(n664), .I2(EX_adresse[18]), .O(n1048) );
  NAND_GATE U1201 ( .I1(n665), .I2(n199), .O(n1046) );
  NAND3_GATE U1202 ( .I1(n1051), .I2(n1052), .I3(n1053), .O(n199) );
  NAND_GATE U1203 ( .I1(n669), .I2(N352), .O(n1053) );
  NAND_GATE U1204 ( .I1(\pred_tab[2][BRA_ADR][18] ), .I2(n670), .O(n1052) );
  NAND_GATE U1205 ( .I1(n671), .I2(EX_adresse[18]), .O(n1051) );
  NAND_GATE U1206 ( .I1(n672), .I2(n68), .O(n1045) );
  NAND3_GATE U1207 ( .I1(n1054), .I2(n1055), .I3(n1056), .O(n68) );
  NAND_GATE U1208 ( .I1(N352), .I2(n676), .O(n1056) );
  NAND_GATE U1209 ( .I1(\pred_tab[1][BRA_ADR][18] ), .I2(n677), .O(n1055) );
  NAND_GATE U1210 ( .I1(EX_adresse[18]), .I2(n678), .O(n1054) );
  NAND_GATE U1211 ( .I1(\pred_tab[1][BRA_ADR][18] ), .I2(n679), .O(n1044) );
  NAND_GATE U1212 ( .I1(N1262), .I2(n680), .O(n1042) );
  NAND_GATE U1213 ( .I1(\pred_tab[2][BRA_ADR][18] ), .I2(n681), .O(n1041) );
  NAND_GATE U1214 ( .I1(\pred_tab[3][BRA_ADR][18] ), .I2(n682), .O(n1040) );
  NAND4_GATE U1215 ( .I1(n1057), .I2(n1058), .I3(n1059), .I4(n1060), .O(
        PR_bra_adr[17]) );
  AND4_GATE U1216 ( .I1(n1061), .I2(n1062), .I3(n1063), .I4(n1064), .O(n1060)
         );
  NAND_GATE U1217 ( .I1(n658), .I2(n326), .O(n1064) );
  NAND3_GATE U1218 ( .I1(n1065), .I2(n1066), .I3(n1067), .O(n326) );
  NAND_GATE U1219 ( .I1(n662), .I2(N351), .O(n1067) );
  NAND_GATE U1220 ( .I1(\pred_tab[3][BRA_ADR][17] ), .I2(n663), .O(n1066) );
  NAND_GATE U1221 ( .I1(n664), .I2(EX_adresse[17]), .O(n1065) );
  NAND_GATE U1222 ( .I1(n665), .I2(n195), .O(n1063) );
  NAND3_GATE U1223 ( .I1(n1068), .I2(n1069), .I3(n1070), .O(n195) );
  NAND_GATE U1224 ( .I1(n669), .I2(N351), .O(n1070) );
  NAND_GATE U1225 ( .I1(\pred_tab[2][BRA_ADR][17] ), .I2(n670), .O(n1069) );
  NAND_GATE U1226 ( .I1(n671), .I2(EX_adresse[17]), .O(n1068) );
  NAND_GATE U1227 ( .I1(n672), .I2(n64), .O(n1062) );
  NAND3_GATE U1228 ( .I1(n1071), .I2(n1072), .I3(n1073), .O(n64) );
  NAND_GATE U1229 ( .I1(N351), .I2(n676), .O(n1073) );
  NAND_GATE U1230 ( .I1(\pred_tab[1][BRA_ADR][17] ), .I2(n677), .O(n1072) );
  NAND_GATE U1231 ( .I1(EX_adresse[17]), .I2(n678), .O(n1071) );
  NAND_GATE U1232 ( .I1(\pred_tab[1][BRA_ADR][17] ), .I2(n679), .O(n1061) );
  NAND_GATE U1233 ( .I1(N1261), .I2(n680), .O(n1059) );
  NAND_GATE U1234 ( .I1(\pred_tab[2][BRA_ADR][17] ), .I2(n681), .O(n1058) );
  NAND_GATE U1235 ( .I1(\pred_tab[3][BRA_ADR][17] ), .I2(n682), .O(n1057) );
  NAND4_GATE U1236 ( .I1(n1074), .I2(n1075), .I3(n1076), .I4(n1077), .O(
        PR_bra_adr[16]) );
  AND4_GATE U1237 ( .I1(n1078), .I2(n1079), .I3(n1080), .I4(n1081), .O(n1077)
         );
  NAND_GATE U1238 ( .I1(n658), .I2(n322), .O(n1081) );
  NAND3_GATE U1239 ( .I1(n1082), .I2(n1083), .I3(n1084), .O(n322) );
  NAND_GATE U1240 ( .I1(n662), .I2(N350), .O(n1084) );
  NAND_GATE U1241 ( .I1(\pred_tab[3][BRA_ADR][16] ), .I2(n663), .O(n1083) );
  NAND_GATE U1242 ( .I1(n664), .I2(EX_adresse[16]), .O(n1082) );
  NAND_GATE U1243 ( .I1(n665), .I2(n191), .O(n1080) );
  NAND3_GATE U1244 ( .I1(n1085), .I2(n1086), .I3(n1087), .O(n191) );
  NAND_GATE U1245 ( .I1(n669), .I2(N350), .O(n1087) );
  NAND_GATE U1246 ( .I1(\pred_tab[2][BRA_ADR][16] ), .I2(n670), .O(n1086) );
  NAND_GATE U1247 ( .I1(n671), .I2(EX_adresse[16]), .O(n1085) );
  NAND_GATE U1248 ( .I1(n672), .I2(n60), .O(n1079) );
  NAND3_GATE U1249 ( .I1(n1088), .I2(n1089), .I3(n1090), .O(n60) );
  NAND_GATE U1250 ( .I1(N350), .I2(n676), .O(n1090) );
  NAND_GATE U1251 ( .I1(\pred_tab[1][BRA_ADR][16] ), .I2(n677), .O(n1089) );
  NAND_GATE U1252 ( .I1(EX_adresse[16]), .I2(n678), .O(n1088) );
  NAND_GATE U1253 ( .I1(\pred_tab[1][BRA_ADR][16] ), .I2(n679), .O(n1078) );
  NAND_GATE U1254 ( .I1(N1260), .I2(n680), .O(n1076) );
  NAND_GATE U1255 ( .I1(\pred_tab[2][BRA_ADR][16] ), .I2(n681), .O(n1075) );
  NAND_GATE U1256 ( .I1(\pred_tab[3][BRA_ADR][16] ), .I2(n682), .O(n1074) );
  NAND4_GATE U1257 ( .I1(n1091), .I2(n1092), .I3(n1093), .I4(n1094), .O(
        PR_bra_adr[15]) );
  AND4_GATE U1258 ( .I1(n1095), .I2(n1096), .I3(n1097), .I4(n1098), .O(n1094)
         );
  NAND_GATE U1259 ( .I1(n658), .I2(n318), .O(n1098) );
  NAND3_GATE U1260 ( .I1(n1099), .I2(n1100), .I3(n1101), .O(n318) );
  NAND_GATE U1261 ( .I1(n662), .I2(N349), .O(n1101) );
  NAND_GATE U1262 ( .I1(\pred_tab[3][BRA_ADR][15] ), .I2(n663), .O(n1100) );
  NAND_GATE U1263 ( .I1(n664), .I2(EX_adresse[15]), .O(n1099) );
  NAND_GATE U1264 ( .I1(n665), .I2(n187), .O(n1097) );
  NAND3_GATE U1265 ( .I1(n1102), .I2(n1103), .I3(n1104), .O(n187) );
  NAND_GATE U1266 ( .I1(n669), .I2(N349), .O(n1104) );
  NAND_GATE U1267 ( .I1(\pred_tab[2][BRA_ADR][15] ), .I2(n670), .O(n1103) );
  NAND_GATE U1268 ( .I1(n671), .I2(EX_adresse[15]), .O(n1102) );
  NAND_GATE U1269 ( .I1(n672), .I2(n56), .O(n1096) );
  NAND3_GATE U1270 ( .I1(n1105), .I2(n1106), .I3(n1107), .O(n56) );
  NAND_GATE U1271 ( .I1(N349), .I2(n676), .O(n1107) );
  NAND_GATE U1272 ( .I1(\pred_tab[1][BRA_ADR][15] ), .I2(n677), .O(n1106) );
  NAND_GATE U1273 ( .I1(EX_adresse[15]), .I2(n678), .O(n1105) );
  NAND_GATE U1274 ( .I1(\pred_tab[1][BRA_ADR][15] ), .I2(n679), .O(n1095) );
  NAND_GATE U1275 ( .I1(N1259), .I2(n680), .O(n1093) );
  NAND_GATE U1276 ( .I1(\pred_tab[2][BRA_ADR][15] ), .I2(n681), .O(n1092) );
  NAND_GATE U1277 ( .I1(\pred_tab[3][BRA_ADR][15] ), .I2(n682), .O(n1091) );
  NAND4_GATE U1278 ( .I1(n1108), .I2(n1109), .I3(n1110), .I4(n1111), .O(
        PR_bra_adr[14]) );
  AND4_GATE U1279 ( .I1(n1112), .I2(n1113), .I3(n1114), .I4(n1115), .O(n1111)
         );
  NAND_GATE U1280 ( .I1(n658), .I2(n314), .O(n1115) );
  NAND3_GATE U1281 ( .I1(n1116), .I2(n1117), .I3(n1118), .O(n314) );
  NAND_GATE U1282 ( .I1(n662), .I2(N348), .O(n1118) );
  NAND_GATE U1283 ( .I1(\pred_tab[3][BRA_ADR][14] ), .I2(n663), .O(n1117) );
  NAND_GATE U1284 ( .I1(n664), .I2(EX_adresse[14]), .O(n1116) );
  NAND_GATE U1285 ( .I1(n665), .I2(n183), .O(n1114) );
  NAND3_GATE U1286 ( .I1(n1119), .I2(n1120), .I3(n1121), .O(n183) );
  NAND_GATE U1287 ( .I1(n669), .I2(N348), .O(n1121) );
  NAND_GATE U1288 ( .I1(\pred_tab[2][BRA_ADR][14] ), .I2(n670), .O(n1120) );
  NAND_GATE U1289 ( .I1(n671), .I2(EX_adresse[14]), .O(n1119) );
  NAND_GATE U1290 ( .I1(n672), .I2(n52), .O(n1113) );
  NAND3_GATE U1291 ( .I1(n1122), .I2(n1123), .I3(n1124), .O(n52) );
  NAND_GATE U1292 ( .I1(N348), .I2(n676), .O(n1124) );
  NAND_GATE U1293 ( .I1(\pred_tab[1][BRA_ADR][14] ), .I2(n677), .O(n1123) );
  NAND_GATE U1294 ( .I1(EX_adresse[14]), .I2(n678), .O(n1122) );
  NAND_GATE U1295 ( .I1(\pred_tab[1][BRA_ADR][14] ), .I2(n679), .O(n1112) );
  NAND_GATE U1296 ( .I1(N1258), .I2(n680), .O(n1110) );
  NAND_GATE U1297 ( .I1(\pred_tab[2][BRA_ADR][14] ), .I2(n681), .O(n1109) );
  NAND_GATE U1298 ( .I1(\pred_tab[3][BRA_ADR][14] ), .I2(n682), .O(n1108) );
  NAND4_GATE U1299 ( .I1(n1125), .I2(n1126), .I3(n1127), .I4(n1128), .O(
        PR_bra_adr[13]) );
  AND4_GATE U1300 ( .I1(n1129), .I2(n1130), .I3(n1131), .I4(n1132), .O(n1128)
         );
  NAND_GATE U1301 ( .I1(n658), .I2(n310), .O(n1132) );
  NAND3_GATE U1302 ( .I1(n1133), .I2(n1134), .I3(n1135), .O(n310) );
  NAND_GATE U1303 ( .I1(n662), .I2(N347), .O(n1135) );
  NAND_GATE U1304 ( .I1(\pred_tab[3][BRA_ADR][13] ), .I2(n663), .O(n1134) );
  NAND_GATE U1305 ( .I1(n664), .I2(EX_adresse[13]), .O(n1133) );
  NAND_GATE U1306 ( .I1(n665), .I2(n179), .O(n1131) );
  NAND3_GATE U1307 ( .I1(n1136), .I2(n1137), .I3(n1138), .O(n179) );
  NAND_GATE U1308 ( .I1(n669), .I2(N347), .O(n1138) );
  NAND_GATE U1309 ( .I1(\pred_tab[2][BRA_ADR][13] ), .I2(n670), .O(n1137) );
  NAND_GATE U1310 ( .I1(n671), .I2(EX_adresse[13]), .O(n1136) );
  NAND_GATE U1311 ( .I1(n672), .I2(n48), .O(n1130) );
  NAND3_GATE U1312 ( .I1(n1139), .I2(n1140), .I3(n1141), .O(n48) );
  NAND_GATE U1313 ( .I1(N347), .I2(n676), .O(n1141) );
  NAND_GATE U1314 ( .I1(\pred_tab[1][BRA_ADR][13] ), .I2(n677), .O(n1140) );
  NAND_GATE U1315 ( .I1(EX_adresse[13]), .I2(n678), .O(n1139) );
  NAND_GATE U1316 ( .I1(\pred_tab[1][BRA_ADR][13] ), .I2(n679), .O(n1129) );
  NAND_GATE U1317 ( .I1(N1257), .I2(n680), .O(n1127) );
  NAND_GATE U1318 ( .I1(\pred_tab[2][BRA_ADR][13] ), .I2(n681), .O(n1126) );
  NAND_GATE U1319 ( .I1(\pred_tab[3][BRA_ADR][13] ), .I2(n682), .O(n1125) );
  NAND4_GATE U1320 ( .I1(n1142), .I2(n1143), .I3(n1144), .I4(n1145), .O(
        PR_bra_adr[12]) );
  AND4_GATE U1321 ( .I1(n1146), .I2(n1147), .I3(n1148), .I4(n1149), .O(n1145)
         );
  NAND_GATE U1322 ( .I1(n658), .I2(n306), .O(n1149) );
  NAND3_GATE U1323 ( .I1(n1150), .I2(n1151), .I3(n1152), .O(n306) );
  NAND_GATE U1324 ( .I1(n662), .I2(N346), .O(n1152) );
  NAND_GATE U1325 ( .I1(\pred_tab[3][BRA_ADR][12] ), .I2(n663), .O(n1151) );
  NAND_GATE U1326 ( .I1(n664), .I2(EX_adresse[12]), .O(n1150) );
  NAND_GATE U1327 ( .I1(n665), .I2(n175), .O(n1148) );
  NAND3_GATE U1328 ( .I1(n1153), .I2(n1154), .I3(n1155), .O(n175) );
  NAND_GATE U1329 ( .I1(n669), .I2(N346), .O(n1155) );
  NAND_GATE U1330 ( .I1(\pred_tab[2][BRA_ADR][12] ), .I2(n670), .O(n1154) );
  NAND_GATE U1331 ( .I1(n671), .I2(EX_adresse[12]), .O(n1153) );
  NAND_GATE U1332 ( .I1(n672), .I2(n44), .O(n1147) );
  NAND3_GATE U1333 ( .I1(n1156), .I2(n1157), .I3(n1158), .O(n44) );
  NAND_GATE U1334 ( .I1(N346), .I2(n676), .O(n1158) );
  NAND_GATE U1335 ( .I1(\pred_tab[1][BRA_ADR][12] ), .I2(n677), .O(n1157) );
  NAND_GATE U1336 ( .I1(EX_adresse[12]), .I2(n678), .O(n1156) );
  NAND_GATE U1337 ( .I1(\pred_tab[1][BRA_ADR][12] ), .I2(n679), .O(n1146) );
  NAND_GATE U1338 ( .I1(N1256), .I2(n680), .O(n1144) );
  NAND_GATE U1339 ( .I1(\pred_tab[2][BRA_ADR][12] ), .I2(n681), .O(n1143) );
  NAND_GATE U1340 ( .I1(\pred_tab[3][BRA_ADR][12] ), .I2(n682), .O(n1142) );
  NAND4_GATE U1341 ( .I1(n1159), .I2(n1160), .I3(n1161), .I4(n1162), .O(
        PR_bra_adr[11]) );
  AND4_GATE U1342 ( .I1(n1163), .I2(n1164), .I3(n1165), .I4(n1166), .O(n1162)
         );
  NAND_GATE U1343 ( .I1(n658), .I2(n302), .O(n1166) );
  NAND3_GATE U1344 ( .I1(n1167), .I2(n1168), .I3(n1169), .O(n302) );
  NAND_GATE U1345 ( .I1(n662), .I2(N345), .O(n1169) );
  NAND_GATE U1346 ( .I1(\pred_tab[3][BRA_ADR][11] ), .I2(n663), .O(n1168) );
  NAND_GATE U1347 ( .I1(n664), .I2(EX_adresse[11]), .O(n1167) );
  NAND_GATE U1348 ( .I1(n665), .I2(n171), .O(n1165) );
  NAND3_GATE U1349 ( .I1(n1170), .I2(n1171), .I3(n1172), .O(n171) );
  NAND_GATE U1350 ( .I1(n669), .I2(N345), .O(n1172) );
  NAND_GATE U1351 ( .I1(\pred_tab[2][BRA_ADR][11] ), .I2(n670), .O(n1171) );
  NAND_GATE U1352 ( .I1(n671), .I2(EX_adresse[11]), .O(n1170) );
  NAND_GATE U1353 ( .I1(n672), .I2(n40), .O(n1164) );
  NAND3_GATE U1354 ( .I1(n1173), .I2(n1174), .I3(n1175), .O(n40) );
  NAND_GATE U1355 ( .I1(N345), .I2(n676), .O(n1175) );
  NAND_GATE U1356 ( .I1(\pred_tab[1][BRA_ADR][11] ), .I2(n677), .O(n1174) );
  NAND_GATE U1357 ( .I1(EX_adresse[11]), .I2(n678), .O(n1173) );
  NAND_GATE U1358 ( .I1(\pred_tab[1][BRA_ADR][11] ), .I2(n679), .O(n1163) );
  NAND_GATE U1359 ( .I1(N1255), .I2(n680), .O(n1161) );
  NAND_GATE U1360 ( .I1(\pred_tab[2][BRA_ADR][11] ), .I2(n681), .O(n1160) );
  NAND_GATE U1361 ( .I1(\pred_tab[3][BRA_ADR][11] ), .I2(n682), .O(n1159) );
  NAND4_GATE U1362 ( .I1(n1176), .I2(n1177), .I3(n1178), .I4(n1179), .O(
        PR_bra_adr[10]) );
  AND4_GATE U1363 ( .I1(n1180), .I2(n1181), .I3(n1182), .I4(n1183), .O(n1179)
         );
  NAND_GATE U1364 ( .I1(n658), .I2(n298), .O(n1183) );
  NAND3_GATE U1365 ( .I1(n1184), .I2(n1185), .I3(n1186), .O(n298) );
  NAND_GATE U1366 ( .I1(n662), .I2(N344), .O(n1186) );
  NAND_GATE U1367 ( .I1(\pred_tab[3][BRA_ADR][10] ), .I2(n663), .O(n1185) );
  NAND_GATE U1368 ( .I1(n664), .I2(EX_adresse[10]), .O(n1184) );
  NAND_GATE U1369 ( .I1(n665), .I2(n167), .O(n1182) );
  NAND3_GATE U1370 ( .I1(n1187), .I2(n1188), .I3(n1189), .O(n167) );
  NAND_GATE U1371 ( .I1(n669), .I2(N344), .O(n1189) );
  NAND_GATE U1372 ( .I1(\pred_tab[2][BRA_ADR][10] ), .I2(n670), .O(n1188) );
  NAND_GATE U1373 ( .I1(n671), .I2(EX_adresse[10]), .O(n1187) );
  NAND_GATE U1374 ( .I1(n672), .I2(n35), .O(n1181) );
  NAND3_GATE U1375 ( .I1(n1190), .I2(n1191), .I3(n1192), .O(n35) );
  NAND_GATE U1376 ( .I1(N344), .I2(n676), .O(n1192) );
  NAND_GATE U1377 ( .I1(\pred_tab[1][BRA_ADR][10] ), .I2(n677), .O(n1191) );
  NAND_GATE U1378 ( .I1(EX_adresse[10]), .I2(n678), .O(n1190) );
  NAND_GATE U1379 ( .I1(\pred_tab[1][BRA_ADR][10] ), .I2(n679), .O(n1180) );
  NAND_GATE U1380 ( .I1(N1254), .I2(n680), .O(n1178) );
  NAND_GATE U1381 ( .I1(\pred_tab[2][BRA_ADR][10] ), .I2(n681), .O(n1177) );
  NAND_GATE U1382 ( .I1(\pred_tab[3][BRA_ADR][10] ), .I2(n682), .O(n1176) );
  NAND4_GATE U1383 ( .I1(n1193), .I2(n1194), .I3(n1195), .I4(n1196), .O(
        PR_bra_adr[0]) );
  AND4_GATE U1384 ( .I1(n1197), .I2(n1198), .I3(n1199), .I4(n1200), .O(n1196)
         );
  NAND_GATE U1385 ( .I1(n658), .I2(n293), .O(n1200) );
  NAND3_GATE U1386 ( .I1(n1201), .I2(n1202), .I3(n1203), .O(n293) );
  NAND_GATE U1387 ( .I1(n662), .I2(N334), .O(n1203) );
  AND_GATE U1388 ( .I1(n1204), .I2(n440), .O(n662) );
  NAND_GATE U1389 ( .I1(\pred_tab[3][BRA_ADR][0] ), .I2(n663), .O(n1202) );
  NAND_GATE U1390 ( .I1(n1205), .I2(n440), .O(n663) );
  NAND_GATE U1391 ( .I1(n664), .I2(EX_adresse[0]), .O(n1201) );
  AND_GATE U1392 ( .I1(n440), .I2(n1206), .O(n664) );
  AND_GATE U1393 ( .I1(n1207), .I2(n441), .O(n658) );
  NAND_GATE U1394 ( .I1(n665), .I2(n162), .O(n1199) );
  NAND3_GATE U1395 ( .I1(n1208), .I2(n1209), .I3(n1210), .O(n162) );
  NAND_GATE U1396 ( .I1(N334), .I2(n669), .O(n1210) );
  AND_GATE U1397 ( .I1(n425), .I2(n1204), .O(n669) );
  NAND_GATE U1398 ( .I1(\pred_tab[2][BRA_ADR][0] ), .I2(n670), .O(n1209) );
  NAND_GATE U1399 ( .I1(n425), .I2(n1205), .O(n670) );
  NAND_GATE U1400 ( .I1(EX_adresse[0]), .I2(n671), .O(n1208) );
  AND_GATE U1401 ( .I1(n425), .I2(n1206), .O(n671) );
  AND_GATE U1402 ( .I1(n1211), .I2(n1212), .O(n425) );
  AND_GATE U1403 ( .I1(n1213), .I2(n447), .O(n665) );
  NAND_GATE U1405 ( .I1(n672), .I2(n422), .O(n1198) );
  NAND3_GATE U1406 ( .I1(n1214), .I2(n1215), .I3(n1216), .O(n422) );
  NAND_GATE U1407 ( .I1(N334), .I2(n676), .O(n1216) );
  AND_GATE U1408 ( .I1(n1204), .I2(n433), .O(n676) );
  NOR_GATE U1409 ( .I1(n1217), .I2(EX_bra_confirm), .O(n1204) );
  NAND_GATE U1410 ( .I1(\pred_tab[1][BRA_ADR][0] ), .I2(n677), .O(n1215) );
  NAND_GATE U1411 ( .I1(n1205), .I2(n433), .O(n677) );
  NAND_GATE U1412 ( .I1(EX_adresse[0]), .I2(n678), .O(n1214) );
  AND_GATE U1413 ( .I1(n433), .I2(n1206), .O(n678) );
  NAND_GATE U1414 ( .I1(n1218), .I2(n1219), .O(n1206) );
  NAND_GATE U1415 ( .I1(n1223), .I2(EX_bra_confirm), .O(n1219) );
  NAND_GATE U1416 ( .I1(N599), .I2(n1217), .O(n1218) );
  NOR_GATE U1417 ( .I1(n1212), .I2(n1211), .O(n433) );
  AND_GATE U1418 ( .I1(n1221), .I2(n577), .O(n672) );
  NAND_GATE U1420 ( .I1(\pred_tab[1][BRA_ADR][0] ), .I2(n679), .O(n1197) );
  AND_GATE U1421 ( .I1(n1222), .I2(n1229), .O(n679) );
  NAND_GATE U1422 ( .I1(N1244), .I2(n680), .O(n1195) );
  NAND3_GATE U1423 ( .I1(n1224), .I2(n1225), .I3(n1226), .O(n680) );
  NAND_GATE U1424 ( .I1(n1221), .I2(n29), .O(n1226) );
  AND3_GATE U1425 ( .I1(\next_out[0] ), .I2(n1238), .I3(n646), .O(n29) );
  NOR_GATE U1427 ( .I1(n1228), .I2(n1212), .O(n1221) );
  NAND_GATE U1428 ( .I1(n1207), .I2(n642), .O(n1225) );
  OR_GATE U1430 ( .I1(n647), .I2(N1582), .O(n441) );
  AND_GATE U1431 ( .I1(PR_clear), .I2(n440), .O(n1207) );
  NAND_GATE U1432 ( .I1(n1213), .I2(n28), .O(n1224) );
  AND3_GATE U1433 ( .I1(\next_out[1] ), .I2(n512), .I3(n646), .O(n28) );
  NAND4_GATE U1435 ( .I1(DI_bra), .I2(n1230), .I3(n1231), .I4(n1232), .O(n647)
         );
  NAND_GATE U1436 ( .I1(\pred_tab[1][IS_AFFECTED] ), .I2(N70), .O(n1232) );
  NAND_GATE U1437 ( .I1(\pred_tab[2][IS_AFFECTED] ), .I2(N79), .O(n1231) );
  NAND_GATE U1438 ( .I1(\pred_tab[3][IS_AFFECTED] ), .I2(N96), .O(n1230) );
  AND_GATE U1440 ( .I1(PR_clear), .I2(n1211), .O(n1213) );
  NAND_GATE U1442 ( .I1(\pred_tab[2][BRA_ADR][0] ), .I2(n681), .O(n1194) );
  AND_GATE U1443 ( .I1(n1222), .I2(n1233), .O(n681) );
  NAND_GATE U1444 ( .I1(\pred_tab[3][BRA_ADR][0] ), .I2(n682), .O(n1193) );
  AND3_GATE U1445 ( .I1(n1234), .I2(n1235), .I3(n1222), .O(n682) );
  AND_GATE U1446 ( .I1(N1579), .I2(n1228), .O(n1222) );
  NAND_GATE U1447 ( .I1(n1205), .I2(EX_uncleared), .O(n1228) );
  AND_GATE U1448 ( .I1(n1236), .I2(n1237), .O(n1205) );
  NAND_GATE U1449 ( .I1(n1211), .I2(n1227), .O(n1237) );
  OR_GATE U1450 ( .I1(n1223), .I2(N599), .O(n1236) );
  NAND_GATE U1452 ( .I1(n1239), .I2(n1240), .O(n1217) );
  NAND_GATE U1453 ( .I1(EX_bra_confirm), .I2(n1241), .O(n1240) );
  OR_GATE U1454 ( .I1(n1241), .I2(EX_bra_confirm), .O(n1239) );
  NAND3_GATE U1455 ( .I1(n1242), .I2(n1243), .I3(n1244), .O(n1241) );
  NAND_GATE U1456 ( .I1(\pred_tab[2][LAST_BRA] ), .I2(n1211), .O(n1244) );
  NAND_GATE U1457 ( .I1(\pred_tab[3][LAST_BRA] ), .I2(n440), .O(n1243) );
  NAND_GATE U1458 ( .I1(\pred_tab[1][LAST_BRA] ), .I2(n1227), .O(n1242) );
  NAND3_GATE U1459 ( .I1(n1245), .I2(n1246), .I3(n1247), .O(N598) );
  NAND_GATE U1460 ( .I1(\pred_tab[2][BRA_ADR][0] ), .I2(n1211), .O(n1247) );
  NAND_GATE U1461 ( .I1(\pred_tab[3][BRA_ADR][0] ), .I2(n440), .O(n1246) );
  NAND_GATE U1462 ( .I1(\pred_tab[1][BRA_ADR][0] ), .I2(n1227), .O(n1245) );
  NAND3_GATE U1463 ( .I1(n1248), .I2(n1249), .I3(n1250), .O(N597) );
  NAND_GATE U1464 ( .I1(\pred_tab[2][BRA_ADR][1] ), .I2(n1211), .O(n1250) );
  NAND_GATE U1465 ( .I1(\pred_tab[3][BRA_ADR][1] ), .I2(n440), .O(n1249) );
  NAND_GATE U1466 ( .I1(\pred_tab[1][BRA_ADR][1] ), .I2(n1227), .O(n1248) );
  NAND3_GATE U1467 ( .I1(n1251), .I2(n1252), .I3(n1253), .O(N596) );
  NAND_GATE U1468 ( .I1(\pred_tab[2][BRA_ADR][2] ), .I2(n1211), .O(n1253) );
  NAND_GATE U1469 ( .I1(\pred_tab[3][BRA_ADR][2] ), .I2(n440), .O(n1252) );
  NAND_GATE U1470 ( .I1(\pred_tab[1][BRA_ADR][2] ), .I2(n1227), .O(n1251) );
  NAND3_GATE U1471 ( .I1(n1254), .I2(n1255), .I3(n1256), .O(N595) );
  NAND_GATE U1472 ( .I1(\pred_tab[2][BRA_ADR][3] ), .I2(n1211), .O(n1256) );
  NAND_GATE U1473 ( .I1(\pred_tab[3][BRA_ADR][3] ), .I2(n440), .O(n1255) );
  NAND_GATE U1474 ( .I1(\pred_tab[1][BRA_ADR][3] ), .I2(n1227), .O(n1254) );
  NAND3_GATE U1475 ( .I1(n1257), .I2(n1258), .I3(n1259), .O(N594) );
  NAND_GATE U1476 ( .I1(\pred_tab[2][BRA_ADR][4] ), .I2(n1211), .O(n1259) );
  NAND_GATE U1477 ( .I1(\pred_tab[3][BRA_ADR][4] ), .I2(n440), .O(n1258) );
  NAND_GATE U1478 ( .I1(\pred_tab[1][BRA_ADR][4] ), .I2(n1227), .O(n1257) );
  NAND3_GATE U1479 ( .I1(n1260), .I2(n1261), .I3(n1262), .O(N593) );
  NAND_GATE U1480 ( .I1(\pred_tab[2][BRA_ADR][5] ), .I2(n1211), .O(n1262) );
  NAND_GATE U1481 ( .I1(\pred_tab[3][BRA_ADR][5] ), .I2(n440), .O(n1261) );
  NAND_GATE U1482 ( .I1(\pred_tab[1][BRA_ADR][5] ), .I2(n1227), .O(n1260) );
  NAND3_GATE U1483 ( .I1(n1263), .I2(n1264), .I3(n1265), .O(N592) );
  NAND_GATE U1484 ( .I1(\pred_tab[2][BRA_ADR][6] ), .I2(n1211), .O(n1265) );
  NAND_GATE U1485 ( .I1(\pred_tab[3][BRA_ADR][6] ), .I2(n440), .O(n1264) );
  NAND_GATE U1486 ( .I1(\pred_tab[1][BRA_ADR][6] ), .I2(n1227), .O(n1263) );
  NAND3_GATE U1487 ( .I1(n1266), .I2(n1267), .I3(n1268), .O(N591) );
  NAND_GATE U1488 ( .I1(\pred_tab[2][BRA_ADR][7] ), .I2(n1211), .O(n1268) );
  NAND_GATE U1489 ( .I1(\pred_tab[3][BRA_ADR][7] ), .I2(n440), .O(n1267) );
  NAND_GATE U1490 ( .I1(\pred_tab[1][BRA_ADR][7] ), .I2(n1227), .O(n1266) );
  NAND3_GATE U1491 ( .I1(n1269), .I2(n1270), .I3(n1271), .O(N590) );
  NAND_GATE U1492 ( .I1(\pred_tab[2][BRA_ADR][8] ), .I2(n1211), .O(n1271) );
  NAND_GATE U1493 ( .I1(\pred_tab[3][BRA_ADR][8] ), .I2(n440), .O(n1270) );
  NAND_GATE U1494 ( .I1(\pred_tab[1][BRA_ADR][8] ), .I2(n1227), .O(n1269) );
  NAND3_GATE U1495 ( .I1(n1272), .I2(n1273), .I3(n1274), .O(N589) );
  NAND_GATE U1496 ( .I1(\pred_tab[2][BRA_ADR][9] ), .I2(n1211), .O(n1274) );
  NAND_GATE U1497 ( .I1(\pred_tab[3][BRA_ADR][9] ), .I2(n440), .O(n1273) );
  NAND_GATE U1498 ( .I1(\pred_tab[1][BRA_ADR][9] ), .I2(n1227), .O(n1272) );
  NAND3_GATE U1499 ( .I1(n1275), .I2(n1276), .I3(n1277), .O(N588) );
  NAND_GATE U1500 ( .I1(\pred_tab[2][BRA_ADR][10] ), .I2(n1211), .O(n1277) );
  NAND_GATE U1501 ( .I1(\pred_tab[3][BRA_ADR][10] ), .I2(n440), .O(n1276) );
  NAND_GATE U1502 ( .I1(\pred_tab[1][BRA_ADR][10] ), .I2(n1227), .O(n1275) );
  NAND3_GATE U1503 ( .I1(n1278), .I2(n1279), .I3(n1280), .O(N587) );
  NAND_GATE U1504 ( .I1(\pred_tab[2][BRA_ADR][11] ), .I2(n1211), .O(n1280) );
  NAND_GATE U1505 ( .I1(\pred_tab[3][BRA_ADR][11] ), .I2(n440), .O(n1279) );
  NAND_GATE U1506 ( .I1(\pred_tab[1][BRA_ADR][11] ), .I2(n1227), .O(n1278) );
  NAND3_GATE U1507 ( .I1(n1281), .I2(n1282), .I3(n1283), .O(N586) );
  NAND_GATE U1508 ( .I1(\pred_tab[2][BRA_ADR][12] ), .I2(n1211), .O(n1283) );
  NAND_GATE U1509 ( .I1(\pred_tab[3][BRA_ADR][12] ), .I2(n440), .O(n1282) );
  NAND_GATE U1510 ( .I1(\pred_tab[1][BRA_ADR][12] ), .I2(n1227), .O(n1281) );
  NAND3_GATE U1511 ( .I1(n1284), .I2(n1285), .I3(n1286), .O(N585) );
  NAND_GATE U1512 ( .I1(\pred_tab[2][BRA_ADR][13] ), .I2(n1211), .O(n1286) );
  NAND_GATE U1513 ( .I1(\pred_tab[3][BRA_ADR][13] ), .I2(n440), .O(n1285) );
  NAND_GATE U1514 ( .I1(\pred_tab[1][BRA_ADR][13] ), .I2(n1227), .O(n1284) );
  NAND3_GATE U1515 ( .I1(n1287), .I2(n1288), .I3(n1289), .O(N584) );
  NAND_GATE U1516 ( .I1(\pred_tab[2][BRA_ADR][14] ), .I2(n1211), .O(n1289) );
  NAND_GATE U1517 ( .I1(\pred_tab[3][BRA_ADR][14] ), .I2(n440), .O(n1288) );
  NAND_GATE U1518 ( .I1(\pred_tab[1][BRA_ADR][14] ), .I2(n1227), .O(n1287) );
  NAND3_GATE U1519 ( .I1(n1290), .I2(n1291), .I3(n1292), .O(N583) );
  NAND_GATE U1520 ( .I1(\pred_tab[2][BRA_ADR][15] ), .I2(n1211), .O(n1292) );
  NAND_GATE U1521 ( .I1(\pred_tab[3][BRA_ADR][15] ), .I2(n440), .O(n1291) );
  NAND_GATE U1522 ( .I1(\pred_tab[1][BRA_ADR][15] ), .I2(n1227), .O(n1290) );
  NAND3_GATE U1523 ( .I1(n1293), .I2(n1294), .I3(n1295), .O(N582) );
  NAND_GATE U1524 ( .I1(\pred_tab[2][BRA_ADR][16] ), .I2(n1211), .O(n1295) );
  NAND_GATE U1525 ( .I1(\pred_tab[3][BRA_ADR][16] ), .I2(n440), .O(n1294) );
  NAND_GATE U1526 ( .I1(\pred_tab[1][BRA_ADR][16] ), .I2(n1227), .O(n1293) );
  NAND3_GATE U1527 ( .I1(n1296), .I2(n1297), .I3(n1298), .O(N581) );
  NAND_GATE U1528 ( .I1(\pred_tab[2][BRA_ADR][17] ), .I2(n1211), .O(n1298) );
  NAND_GATE U1529 ( .I1(\pred_tab[3][BRA_ADR][17] ), .I2(n440), .O(n1297) );
  NAND_GATE U1530 ( .I1(\pred_tab[1][BRA_ADR][17] ), .I2(n1227), .O(n1296) );
  NAND3_GATE U1531 ( .I1(n1299), .I2(n1300), .I3(n1301), .O(N580) );
  NAND_GATE U1532 ( .I1(\pred_tab[2][BRA_ADR][18] ), .I2(n1211), .O(n1301) );
  NAND_GATE U1533 ( .I1(\pred_tab[3][BRA_ADR][18] ), .I2(n440), .O(n1300) );
  NAND_GATE U1534 ( .I1(\pred_tab[1][BRA_ADR][18] ), .I2(n1227), .O(n1299) );
  NAND3_GATE U1535 ( .I1(n1302), .I2(n1303), .I3(n1304), .O(N579) );
  NAND_GATE U1536 ( .I1(\pred_tab[2][BRA_ADR][19] ), .I2(n1211), .O(n1304) );
  NAND_GATE U1537 ( .I1(\pred_tab[3][BRA_ADR][19] ), .I2(n440), .O(n1303) );
  NAND_GATE U1538 ( .I1(\pred_tab[1][BRA_ADR][19] ), .I2(n1227), .O(n1302) );
  NAND3_GATE U1539 ( .I1(n1305), .I2(n1306), .I3(n1307), .O(N578) );
  NAND_GATE U1540 ( .I1(\pred_tab[2][BRA_ADR][20] ), .I2(n1211), .O(n1307) );
  NAND_GATE U1541 ( .I1(\pred_tab[3][BRA_ADR][20] ), .I2(n440), .O(n1306) );
  NAND_GATE U1542 ( .I1(\pred_tab[1][BRA_ADR][20] ), .I2(n1227), .O(n1305) );
  NAND3_GATE U1543 ( .I1(n1308), .I2(n1309), .I3(n1310), .O(N577) );
  NAND_GATE U1544 ( .I1(\pred_tab[2][BRA_ADR][21] ), .I2(n1211), .O(n1310) );
  NAND_GATE U1545 ( .I1(\pred_tab[3][BRA_ADR][21] ), .I2(n440), .O(n1309) );
  NAND_GATE U1546 ( .I1(\pred_tab[1][BRA_ADR][21] ), .I2(n1227), .O(n1308) );
  NAND3_GATE U1547 ( .I1(n1311), .I2(n1312), .I3(n1313), .O(N576) );
  NAND_GATE U1548 ( .I1(\pred_tab[2][BRA_ADR][22] ), .I2(n1211), .O(n1313) );
  NAND_GATE U1549 ( .I1(\pred_tab[3][BRA_ADR][22] ), .I2(n440), .O(n1312) );
  NAND_GATE U1550 ( .I1(\pred_tab[1][BRA_ADR][22] ), .I2(n1227), .O(n1311) );
  NAND3_GATE U1551 ( .I1(n1314), .I2(n1315), .I3(n1316), .O(N575) );
  NAND_GATE U1552 ( .I1(\pred_tab[2][BRA_ADR][23] ), .I2(n1211), .O(n1316) );
  NAND_GATE U1553 ( .I1(\pred_tab[3][BRA_ADR][23] ), .I2(n440), .O(n1315) );
  NAND_GATE U1554 ( .I1(\pred_tab[1][BRA_ADR][23] ), .I2(n1227), .O(n1314) );
  NAND3_GATE U1555 ( .I1(n1317), .I2(n1318), .I3(n1319), .O(N574) );
  NAND_GATE U1556 ( .I1(\pred_tab[2][BRA_ADR][24] ), .I2(n1211), .O(n1319) );
  NAND_GATE U1557 ( .I1(\pred_tab[3][BRA_ADR][24] ), .I2(n440), .O(n1318) );
  NAND_GATE U1558 ( .I1(\pred_tab[1][BRA_ADR][24] ), .I2(n1227), .O(n1317) );
  NAND3_GATE U1559 ( .I1(n1320), .I2(n1321), .I3(n1322), .O(N573) );
  NAND_GATE U1560 ( .I1(\pred_tab[2][BRA_ADR][25] ), .I2(n1211), .O(n1322) );
  NAND_GATE U1561 ( .I1(\pred_tab[3][BRA_ADR][25] ), .I2(n440), .O(n1321) );
  NAND_GATE U1562 ( .I1(\pred_tab[1][BRA_ADR][25] ), .I2(n1227), .O(n1320) );
  NAND3_GATE U1563 ( .I1(n1323), .I2(n1324), .I3(n1325), .O(N572) );
  NAND_GATE U1564 ( .I1(\pred_tab[2][BRA_ADR][26] ), .I2(n1211), .O(n1325) );
  NAND_GATE U1565 ( .I1(\pred_tab[3][BRA_ADR][26] ), .I2(n440), .O(n1324) );
  NAND_GATE U1566 ( .I1(\pred_tab[1][BRA_ADR][26] ), .I2(n1227), .O(n1323) );
  NAND3_GATE U1567 ( .I1(n1326), .I2(n1327), .I3(n1328), .O(N571) );
  NAND_GATE U1568 ( .I1(\pred_tab[2][BRA_ADR][27] ), .I2(n1211), .O(n1328) );
  NAND_GATE U1569 ( .I1(\pred_tab[3][BRA_ADR][27] ), .I2(n440), .O(n1327) );
  NAND_GATE U1570 ( .I1(\pred_tab[1][BRA_ADR][27] ), .I2(n1227), .O(n1326) );
  NAND3_GATE U1571 ( .I1(n1329), .I2(n1330), .I3(n1331), .O(N570) );
  NAND_GATE U1572 ( .I1(\pred_tab[2][BRA_ADR][28] ), .I2(n1211), .O(n1331) );
  NAND_GATE U1573 ( .I1(\pred_tab[3][BRA_ADR][28] ), .I2(n440), .O(n1330) );
  NAND_GATE U1574 ( .I1(\pred_tab[1][BRA_ADR][28] ), .I2(n1227), .O(n1329) );
  NAND3_GATE U1575 ( .I1(n1332), .I2(n1333), .I3(n1334), .O(N569) );
  NAND_GATE U1576 ( .I1(\pred_tab[2][BRA_ADR][29] ), .I2(n1211), .O(n1334) );
  NAND_GATE U1577 ( .I1(\pred_tab[3][BRA_ADR][29] ), .I2(n440), .O(n1333) );
  NAND_GATE U1578 ( .I1(\pred_tab[1][BRA_ADR][29] ), .I2(n1227), .O(n1332) );
  NAND3_GATE U1579 ( .I1(n1335), .I2(n1336), .I3(n1337), .O(N568) );
  NAND_GATE U1580 ( .I1(\pred_tab[2][BRA_ADR][30] ), .I2(n1211), .O(n1337) );
  NAND_GATE U1581 ( .I1(\pred_tab[3][BRA_ADR][30] ), .I2(n440), .O(n1336) );
  NAND_GATE U1582 ( .I1(\pred_tab[1][BRA_ADR][30] ), .I2(n1227), .O(n1335) );
  NAND3_GATE U1583 ( .I1(n1338), .I2(n1339), .I3(n1340), .O(N567) );
  NAND_GATE U1584 ( .I1(\pred_tab[2][BRA_ADR][31] ), .I2(n1211), .O(n1340) );
  NAND_GATE U1585 ( .I1(\pred_tab[3][BRA_ADR][31] ), .I2(n440), .O(n1339) );
  NAND_GATE U1586 ( .I1(\pred_tab[1][BRA_ADR][31] ), .I2(n1227), .O(n1338) );
  NAND3_GATE U1587 ( .I1(n1341), .I2(n1342), .I3(n1343), .O(N333) );
  NAND_GATE U1588 ( .I1(\pred_tab[2][CODE_ADR][0] ), .I2(n1211), .O(n1343) );
  NAND_GATE U1589 ( .I1(\pred_tab[3][CODE_ADR][0] ), .I2(n440), .O(n1342) );
  NAND_GATE U1590 ( .I1(\pred_tab[1][CODE_ADR][0] ), .I2(n1227), .O(n1341) );
  NAND3_GATE U1591 ( .I1(n1344), .I2(n1345), .I3(n1346), .O(N332) );
  NAND_GATE U1592 ( .I1(\pred_tab[2][CODE_ADR][1] ), .I2(n1211), .O(n1346) );
  NAND_GATE U1593 ( .I1(\pred_tab[3][CODE_ADR][1] ), .I2(n440), .O(n1345) );
  NAND_GATE U1594 ( .I1(\pred_tab[1][CODE_ADR][1] ), .I2(n1227), .O(n1344) );
  NAND3_GATE U1595 ( .I1(n1347), .I2(n1348), .I3(n1349), .O(N331) );
  NAND_GATE U1596 ( .I1(\pred_tab[2][CODE_ADR][2] ), .I2(n1211), .O(n1349) );
  NAND_GATE U1597 ( .I1(\pred_tab[3][CODE_ADR][2] ), .I2(n440), .O(n1348) );
  NAND_GATE U1598 ( .I1(\pred_tab[1][CODE_ADR][2] ), .I2(n1227), .O(n1347) );
  NAND3_GATE U1599 ( .I1(n1350), .I2(n1351), .I3(n1352), .O(N330) );
  NAND_GATE U1600 ( .I1(\pred_tab[2][CODE_ADR][3] ), .I2(n1211), .O(n1352) );
  NAND_GATE U1601 ( .I1(\pred_tab[3][CODE_ADR][3] ), .I2(n440), .O(n1351) );
  NAND_GATE U1602 ( .I1(\pred_tab[1][CODE_ADR][3] ), .I2(n1227), .O(n1350) );
  NAND3_GATE U1603 ( .I1(n1353), .I2(n1354), .I3(n1355), .O(N329) );
  NAND_GATE U1604 ( .I1(\pred_tab[2][CODE_ADR][4] ), .I2(n1211), .O(n1355) );
  NAND_GATE U1605 ( .I1(\pred_tab[3][CODE_ADR][4] ), .I2(n440), .O(n1354) );
  NAND_GATE U1606 ( .I1(\pred_tab[1][CODE_ADR][4] ), .I2(n1227), .O(n1353) );
  NAND3_GATE U1607 ( .I1(n1356), .I2(n1357), .I3(n1358), .O(N328) );
  NAND_GATE U1608 ( .I1(\pred_tab[2][CODE_ADR][5] ), .I2(n1211), .O(n1358) );
  NAND_GATE U1609 ( .I1(\pred_tab[3][CODE_ADR][5] ), .I2(n440), .O(n1357) );
  NAND_GATE U1610 ( .I1(\pred_tab[1][CODE_ADR][5] ), .I2(n1227), .O(n1356) );
  NAND3_GATE U1611 ( .I1(n1359), .I2(n1360), .I3(n1361), .O(N327) );
  NAND_GATE U1612 ( .I1(\pred_tab[2][CODE_ADR][6] ), .I2(n1211), .O(n1361) );
  NAND_GATE U1613 ( .I1(\pred_tab[3][CODE_ADR][6] ), .I2(n440), .O(n1360) );
  NAND_GATE U1614 ( .I1(\pred_tab[1][CODE_ADR][6] ), .I2(n1227), .O(n1359) );
  NAND3_GATE U1615 ( .I1(n1362), .I2(n1363), .I3(n1364), .O(N326) );
  NAND_GATE U1616 ( .I1(\pred_tab[2][CODE_ADR][7] ), .I2(n1211), .O(n1364) );
  NAND_GATE U1617 ( .I1(\pred_tab[3][CODE_ADR][7] ), .I2(n440), .O(n1363) );
  NAND_GATE U1618 ( .I1(\pred_tab[1][CODE_ADR][7] ), .I2(n1227), .O(n1362) );
  NAND3_GATE U1619 ( .I1(n1365), .I2(n1366), .I3(n1367), .O(N325) );
  NAND_GATE U1620 ( .I1(\pred_tab[2][CODE_ADR][8] ), .I2(n1211), .O(n1367) );
  NAND_GATE U1621 ( .I1(\pred_tab[3][CODE_ADR][8] ), .I2(n440), .O(n1366) );
  NAND_GATE U1622 ( .I1(\pred_tab[1][CODE_ADR][8] ), .I2(n1227), .O(n1365) );
  NAND3_GATE U1623 ( .I1(n1368), .I2(n1369), .I3(n1370), .O(N324) );
  NAND_GATE U1624 ( .I1(\pred_tab[2][CODE_ADR][9] ), .I2(n1211), .O(n1370) );
  NAND_GATE U1625 ( .I1(\pred_tab[3][CODE_ADR][9] ), .I2(n440), .O(n1369) );
  NAND_GATE U1626 ( .I1(\pred_tab[1][CODE_ADR][9] ), .I2(n1227), .O(n1368) );
  NAND3_GATE U1627 ( .I1(n1371), .I2(n1372), .I3(n1373), .O(N323) );
  NAND_GATE U1628 ( .I1(\pred_tab[2][CODE_ADR][10] ), .I2(n1211), .O(n1373) );
  NAND_GATE U1629 ( .I1(\pred_tab[3][CODE_ADR][10] ), .I2(n440), .O(n1372) );
  NAND_GATE U1630 ( .I1(\pred_tab[1][CODE_ADR][10] ), .I2(n1227), .O(n1371) );
  NAND3_GATE U1631 ( .I1(n1374), .I2(n1375), .I3(n1376), .O(N322) );
  NAND_GATE U1632 ( .I1(\pred_tab[2][CODE_ADR][11] ), .I2(n1211), .O(n1376) );
  NAND_GATE U1633 ( .I1(\pred_tab[3][CODE_ADR][11] ), .I2(n440), .O(n1375) );
  NAND_GATE U1634 ( .I1(\pred_tab[1][CODE_ADR][11] ), .I2(n1227), .O(n1374) );
  NAND3_GATE U1635 ( .I1(n1377), .I2(n1378), .I3(n1379), .O(N321) );
  NAND_GATE U1636 ( .I1(\pred_tab[2][CODE_ADR][12] ), .I2(n1211), .O(n1379) );
  NAND_GATE U1637 ( .I1(\pred_tab[3][CODE_ADR][12] ), .I2(n440), .O(n1378) );
  NAND_GATE U1638 ( .I1(\pred_tab[1][CODE_ADR][12] ), .I2(n1227), .O(n1377) );
  NAND3_GATE U1639 ( .I1(n1380), .I2(n1381), .I3(n1382), .O(N320) );
  NAND_GATE U1640 ( .I1(\pred_tab[2][CODE_ADR][13] ), .I2(n1211), .O(n1382) );
  NAND_GATE U1641 ( .I1(\pred_tab[3][CODE_ADR][13] ), .I2(n440), .O(n1381) );
  NAND_GATE U1642 ( .I1(\pred_tab[1][CODE_ADR][13] ), .I2(n1227), .O(n1380) );
  NAND3_GATE U1643 ( .I1(n1383), .I2(n1384), .I3(n1385), .O(N319) );
  NAND_GATE U1644 ( .I1(\pred_tab[2][CODE_ADR][14] ), .I2(n1211), .O(n1385) );
  NAND_GATE U1645 ( .I1(\pred_tab[3][CODE_ADR][14] ), .I2(n440), .O(n1384) );
  NAND_GATE U1646 ( .I1(\pred_tab[1][CODE_ADR][14] ), .I2(n1227), .O(n1383) );
  NAND3_GATE U1647 ( .I1(n1386), .I2(n1387), .I3(n1388), .O(N318) );
  NAND_GATE U1648 ( .I1(\pred_tab[2][CODE_ADR][15] ), .I2(n1211), .O(n1388) );
  NAND_GATE U1649 ( .I1(\pred_tab[3][CODE_ADR][15] ), .I2(n440), .O(n1387) );
  NAND_GATE U1650 ( .I1(\pred_tab[1][CODE_ADR][15] ), .I2(n1227), .O(n1386) );
  NAND3_GATE U1651 ( .I1(n1389), .I2(n1390), .I3(n1391), .O(N317) );
  NAND_GATE U1652 ( .I1(\pred_tab[2][CODE_ADR][16] ), .I2(n1211), .O(n1391) );
  NAND_GATE U1653 ( .I1(\pred_tab[3][CODE_ADR][16] ), .I2(n440), .O(n1390) );
  NAND_GATE U1654 ( .I1(\pred_tab[1][CODE_ADR][16] ), .I2(n1227), .O(n1389) );
  NAND3_GATE U1655 ( .I1(n1392), .I2(n1393), .I3(n1394), .O(N316) );
  NAND_GATE U1656 ( .I1(\pred_tab[2][CODE_ADR][17] ), .I2(n1211), .O(n1394) );
  NAND_GATE U1657 ( .I1(\pred_tab[3][CODE_ADR][17] ), .I2(n440), .O(n1393) );
  NAND_GATE U1658 ( .I1(\pred_tab[1][CODE_ADR][17] ), .I2(n1227), .O(n1392) );
  NAND3_GATE U1659 ( .I1(n1395), .I2(n1396), .I3(n1397), .O(N315) );
  NAND_GATE U1660 ( .I1(\pred_tab[2][CODE_ADR][18] ), .I2(n1211), .O(n1397) );
  NAND_GATE U1661 ( .I1(\pred_tab[3][CODE_ADR][18] ), .I2(n440), .O(n1396) );
  NAND_GATE U1662 ( .I1(\pred_tab[1][CODE_ADR][18] ), .I2(n1227), .O(n1395) );
  NAND3_GATE U1663 ( .I1(n1398), .I2(n1399), .I3(n1400), .O(N314) );
  NAND_GATE U1664 ( .I1(\pred_tab[2][CODE_ADR][19] ), .I2(n1211), .O(n1400) );
  NAND_GATE U1665 ( .I1(\pred_tab[3][CODE_ADR][19] ), .I2(n440), .O(n1399) );
  NAND_GATE U1666 ( .I1(\pred_tab[1][CODE_ADR][19] ), .I2(n1227), .O(n1398) );
  NAND3_GATE U1667 ( .I1(n1401), .I2(n1402), .I3(n1403), .O(N313) );
  NAND_GATE U1668 ( .I1(\pred_tab[2][CODE_ADR][20] ), .I2(n1211), .O(n1403) );
  NAND_GATE U1669 ( .I1(\pred_tab[3][CODE_ADR][20] ), .I2(n440), .O(n1402) );
  NAND_GATE U1670 ( .I1(\pred_tab[1][CODE_ADR][20] ), .I2(n1227), .O(n1401) );
  NAND3_GATE U1671 ( .I1(n1404), .I2(n1405), .I3(n1406), .O(N312) );
  NAND_GATE U1672 ( .I1(\pred_tab[2][CODE_ADR][21] ), .I2(n1211), .O(n1406) );
  NAND_GATE U1673 ( .I1(\pred_tab[3][CODE_ADR][21] ), .I2(n440), .O(n1405) );
  NAND_GATE U1674 ( .I1(\pred_tab[1][CODE_ADR][21] ), .I2(n1227), .O(n1404) );
  NAND3_GATE U1675 ( .I1(n1407), .I2(n1408), .I3(n1409), .O(N311) );
  NAND_GATE U1676 ( .I1(\pred_tab[2][CODE_ADR][22] ), .I2(n1211), .O(n1409) );
  NAND_GATE U1677 ( .I1(\pred_tab[3][CODE_ADR][22] ), .I2(n440), .O(n1408) );
  NAND_GATE U1678 ( .I1(\pred_tab[1][CODE_ADR][22] ), .I2(n1227), .O(n1407) );
  NAND3_GATE U1679 ( .I1(n1410), .I2(n1411), .I3(n1412), .O(N310) );
  NAND_GATE U1680 ( .I1(\pred_tab[2][CODE_ADR][23] ), .I2(n1211), .O(n1412) );
  NAND_GATE U1681 ( .I1(\pred_tab[3][CODE_ADR][23] ), .I2(n440), .O(n1411) );
  NAND_GATE U1682 ( .I1(\pred_tab[1][CODE_ADR][23] ), .I2(n1227), .O(n1410) );
  NAND3_GATE U1683 ( .I1(n1413), .I2(n1414), .I3(n1415), .O(N309) );
  NAND_GATE U1684 ( .I1(\pred_tab[2][CODE_ADR][24] ), .I2(n1211), .O(n1415) );
  NAND_GATE U1685 ( .I1(\pred_tab[3][CODE_ADR][24] ), .I2(n440), .O(n1414) );
  NAND_GATE U1686 ( .I1(\pred_tab[1][CODE_ADR][24] ), .I2(n1227), .O(n1413) );
  NAND3_GATE U1687 ( .I1(n1416), .I2(n1417), .I3(n1418), .O(N308) );
  NAND_GATE U1688 ( .I1(\pred_tab[2][CODE_ADR][25] ), .I2(n1211), .O(n1418) );
  NAND_GATE U1689 ( .I1(\pred_tab[3][CODE_ADR][25] ), .I2(n440), .O(n1417) );
  NAND_GATE U1690 ( .I1(\pred_tab[1][CODE_ADR][25] ), .I2(n1227), .O(n1416) );
  NAND3_GATE U1691 ( .I1(n1419), .I2(n1420), .I3(n1421), .O(N307) );
  NAND_GATE U1692 ( .I1(\pred_tab[2][CODE_ADR][26] ), .I2(n1211), .O(n1421) );
  NAND_GATE U1693 ( .I1(\pred_tab[3][CODE_ADR][26] ), .I2(n440), .O(n1420) );
  NAND_GATE U1694 ( .I1(\pred_tab[1][CODE_ADR][26] ), .I2(n1227), .O(n1419) );
  NAND3_GATE U1695 ( .I1(n1422), .I2(n1423), .I3(n1424), .O(N306) );
  NAND_GATE U1696 ( .I1(\pred_tab[2][CODE_ADR][27] ), .I2(n1211), .O(n1424) );
  NAND_GATE U1697 ( .I1(\pred_tab[3][CODE_ADR][27] ), .I2(n440), .O(n1423) );
  NAND_GATE U1698 ( .I1(\pred_tab[1][CODE_ADR][27] ), .I2(n1227), .O(n1422) );
  NAND3_GATE U1699 ( .I1(n1425), .I2(n1426), .I3(n1427), .O(N305) );
  NAND_GATE U1700 ( .I1(\pred_tab[2][CODE_ADR][28] ), .I2(n1211), .O(n1427) );
  NAND_GATE U1701 ( .I1(\pred_tab[3][CODE_ADR][28] ), .I2(n440), .O(n1426) );
  NAND_GATE U1702 ( .I1(\pred_tab[1][CODE_ADR][28] ), .I2(n1227), .O(n1425) );
  NAND3_GATE U1703 ( .I1(n1428), .I2(n1429), .I3(n1430), .O(N304) );
  NAND_GATE U1704 ( .I1(\pred_tab[2][CODE_ADR][29] ), .I2(n1211), .O(n1430) );
  NAND_GATE U1705 ( .I1(\pred_tab[3][CODE_ADR][29] ), .I2(n440), .O(n1429) );
  NAND_GATE U1706 ( .I1(\pred_tab[1][CODE_ADR][29] ), .I2(n1227), .O(n1428) );
  NAND3_GATE U1707 ( .I1(n1431), .I2(n1432), .I3(n1433), .O(N303) );
  NAND_GATE U1708 ( .I1(\pred_tab[2][CODE_ADR][30] ), .I2(n1211), .O(n1433) );
  NAND_GATE U1709 ( .I1(\pred_tab[3][CODE_ADR][30] ), .I2(n440), .O(n1432) );
  NAND_GATE U1710 ( .I1(\pred_tab[1][CODE_ADR][30] ), .I2(n1227), .O(n1431) );
  NAND3_GATE U1711 ( .I1(n1434), .I2(n1435), .I3(n1436), .O(N302) );
  NAND_GATE U1712 ( .I1(\pred_tab[2][CODE_ADR][31] ), .I2(n1211), .O(n1436) );
  NAND_GATE U1713 ( .I1(\pred_tab[3][CODE_ADR][31] ), .I2(n440), .O(n1435) );
  NOR_GATE U1714 ( .I1(n1227), .I2(n1211), .O(n440) );
  AND_GATE U1715 ( .I1(n1437), .I2(n1438), .O(n1211) );
  NAND3_GATE U1716 ( .I1(\pred_tab[1][IS_AFFECTED] ), .I2(n1439), .I3(N71), 
        .O(n1438) );
  NAND_GATE U1717 ( .I1(\pred_tab[1][CODE_ADR][31] ), .I2(n1227), .O(n1434) );
  NAND_GATE U1719 ( .I1(n1439), .I2(n1437), .O(n1212) );
  NAND_GATE U1720 ( .I1(N100), .I2(\pred_tab[3][IS_AFFECTED] ), .O(n1437) );
  NAND_GATE U1721 ( .I1(N82), .I2(\pred_tab[2][IS_AFFECTED] ), .O(n1439) );
  NAND_GATE U1722 ( .I1(\next_out[1] ), .I2(\next_out[0] ), .O(N1582) );
  NAND_GATE U1723 ( .I1(n1229), .I2(n1233), .O(N1579) );
  NAND_GATE U1725 ( .I1(n1440), .I2(n1441), .O(n1234) );
  NAND3_GATE U1726 ( .I1(\pred_tab[1][IS_AFFECTED] ), .I2(n1442), .I3(N69), 
        .O(n1441) );
  NAND_GATE U1728 ( .I1(n1442), .I2(n1440), .O(n1235) );
  NAND_GATE U1729 ( .I1(N92), .I2(\pred_tab[3][IS_AFFECTED] ), .O(n1440) );
  NAND_GATE U1730 ( .I1(N76), .I2(\pred_tab[2][IS_AFFECTED] ), .O(n1442) );
  predict_nb_record3_1_DW01_add_0 add_195 ( .A(DI_adr), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N1275, N1274, N1273, 
        N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, 
        N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, 
        N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244}) );
  predict_nb_record3_1_DW01_cmp6_0 ne_172 ( .A({N567, N568, N569, N570, N571, 
        N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, 
        N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, 
        N596, N597, N598}), .B(EX_adresse), .TC(1'b0), .NE(N599) );
  predict_nb_record3_1_DW01_add_1 add_167 ( .A({N302, N303, N304, N305, N306, 
        N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, 
        N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, 
        N331, N332, N333}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, 
        N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, 
        N343, N342, N341, N340, N339, N338, N337, N336, N335, N334}) );
  predict_nb_record3_1_DW01_cmp6_1 eq_145_I3 ( .A(EX_adr), .B({
        \pred_tab[3][CODE_ADR][31] , \pred_tab[3][CODE_ADR][30] , 
        \pred_tab[3][CODE_ADR][29] , \pred_tab[3][CODE_ADR][28] , 
        \pred_tab[3][CODE_ADR][27] , \pred_tab[3][CODE_ADR][26] , 
        \pred_tab[3][CODE_ADR][25] , \pred_tab[3][CODE_ADR][24] , 
        \pred_tab[3][CODE_ADR][23] , \pred_tab[3][CODE_ADR][22] , 
        \pred_tab[3][CODE_ADR][21] , \pred_tab[3][CODE_ADR][20] , 
        \pred_tab[3][CODE_ADR][19] , \pred_tab[3][CODE_ADR][18] , 
        \pred_tab[3][CODE_ADR][17] , \pred_tab[3][CODE_ADR][16] , 
        \pred_tab[3][CODE_ADR][15] , \pred_tab[3][CODE_ADR][14] , 
        \pred_tab[3][CODE_ADR][13] , \pred_tab[3][CODE_ADR][12] , 
        \pred_tab[3][CODE_ADR][11] , \pred_tab[3][CODE_ADR][10] , 
        \pred_tab[3][CODE_ADR][9] , \pred_tab[3][CODE_ADR][8] , 
        \pred_tab[3][CODE_ADR][7] , \pred_tab[3][CODE_ADR][6] , 
        \pred_tab[3][CODE_ADR][5] , \pred_tab[3][CODE_ADR][4] , 
        \pred_tab[3][CODE_ADR][3] , \pred_tab[3][CODE_ADR][2] , 
        \pred_tab[3][CODE_ADR][1] , \pred_tab[3][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N100) );
  predict_nb_record3_1_DW01_cmp6_2 eq_142_I3 ( .A(DI_adr), .B({
        \pred_tab[3][CODE_ADR][31] , \pred_tab[3][CODE_ADR][30] , 
        \pred_tab[3][CODE_ADR][29] , \pred_tab[3][CODE_ADR][28] , 
        \pred_tab[3][CODE_ADR][27] , \pred_tab[3][CODE_ADR][26] , 
        \pred_tab[3][CODE_ADR][25] , \pred_tab[3][CODE_ADR][24] , 
        \pred_tab[3][CODE_ADR][23] , \pred_tab[3][CODE_ADR][22] , 
        \pred_tab[3][CODE_ADR][21] , \pred_tab[3][CODE_ADR][20] , 
        \pred_tab[3][CODE_ADR][19] , \pred_tab[3][CODE_ADR][18] , 
        \pred_tab[3][CODE_ADR][17] , \pred_tab[3][CODE_ADR][16] , 
        \pred_tab[3][CODE_ADR][15] , \pred_tab[3][CODE_ADR][14] , 
        \pred_tab[3][CODE_ADR][13] , \pred_tab[3][CODE_ADR][12] , 
        \pred_tab[3][CODE_ADR][11] , \pred_tab[3][CODE_ADR][10] , 
        \pred_tab[3][CODE_ADR][9] , \pred_tab[3][CODE_ADR][8] , 
        \pred_tab[3][CODE_ADR][7] , \pred_tab[3][CODE_ADR][6] , 
        \pred_tab[3][CODE_ADR][5] , \pred_tab[3][CODE_ADR][4] , 
        \pred_tab[3][CODE_ADR][3] , \pred_tab[3][CODE_ADR][2] , 
        \pred_tab[3][CODE_ADR][1] , \pred_tab[3][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N96) );
  predict_nb_record3_1_DW01_cmp6_3 eq_139_I3 ( .A(PF_pc), .B({
        \pred_tab[3][CODE_ADR][31] , \pred_tab[3][CODE_ADR][30] , 
        \pred_tab[3][CODE_ADR][29] , \pred_tab[3][CODE_ADR][28] , 
        \pred_tab[3][CODE_ADR][27] , \pred_tab[3][CODE_ADR][26] , 
        \pred_tab[3][CODE_ADR][25] , \pred_tab[3][CODE_ADR][24] , 
        \pred_tab[3][CODE_ADR][23] , \pred_tab[3][CODE_ADR][22] , 
        \pred_tab[3][CODE_ADR][21] , \pred_tab[3][CODE_ADR][20] , 
        \pred_tab[3][CODE_ADR][19] , \pred_tab[3][CODE_ADR][18] , 
        \pred_tab[3][CODE_ADR][17] , \pred_tab[3][CODE_ADR][16] , 
        \pred_tab[3][CODE_ADR][15] , \pred_tab[3][CODE_ADR][14] , 
        \pred_tab[3][CODE_ADR][13] , \pred_tab[3][CODE_ADR][12] , 
        \pred_tab[3][CODE_ADR][11] , \pred_tab[3][CODE_ADR][10] , 
        \pred_tab[3][CODE_ADR][9] , \pred_tab[3][CODE_ADR][8] , 
        \pred_tab[3][CODE_ADR][7] , \pred_tab[3][CODE_ADR][6] , 
        \pred_tab[3][CODE_ADR][5] , \pred_tab[3][CODE_ADR][4] , 
        \pred_tab[3][CODE_ADR][3] , \pred_tab[3][CODE_ADR][2] , 
        \pred_tab[3][CODE_ADR][1] , \pred_tab[3][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N92) );
  predict_nb_record3_1_DW01_cmp6_4 eq_145_I2 ( .A(EX_adr), .B({
        \pred_tab[2][CODE_ADR][31] , \pred_tab[2][CODE_ADR][30] , 
        \pred_tab[2][CODE_ADR][29] , \pred_tab[2][CODE_ADR][28] , 
        \pred_tab[2][CODE_ADR][27] , \pred_tab[2][CODE_ADR][26] , 
        \pred_tab[2][CODE_ADR][25] , \pred_tab[2][CODE_ADR][24] , 
        \pred_tab[2][CODE_ADR][23] , \pred_tab[2][CODE_ADR][22] , 
        \pred_tab[2][CODE_ADR][21] , \pred_tab[2][CODE_ADR][20] , 
        \pred_tab[2][CODE_ADR][19] , \pred_tab[2][CODE_ADR][18] , 
        \pred_tab[2][CODE_ADR][17] , \pred_tab[2][CODE_ADR][16] , 
        \pred_tab[2][CODE_ADR][15] , \pred_tab[2][CODE_ADR][14] , 
        \pred_tab[2][CODE_ADR][13] , \pred_tab[2][CODE_ADR][12] , 
        \pred_tab[2][CODE_ADR][11] , \pred_tab[2][CODE_ADR][10] , 
        \pred_tab[2][CODE_ADR][9] , \pred_tab[2][CODE_ADR][8] , 
        \pred_tab[2][CODE_ADR][7] , \pred_tab[2][CODE_ADR][6] , 
        \pred_tab[2][CODE_ADR][5] , \pred_tab[2][CODE_ADR][4] , 
        \pred_tab[2][CODE_ADR][3] , \pred_tab[2][CODE_ADR][2] , 
        \pred_tab[2][CODE_ADR][1] , \pred_tab[2][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N82) );
  predict_nb_record3_1_DW01_cmp6_5 eq_142_I2 ( .A(DI_adr), .B({
        \pred_tab[2][CODE_ADR][31] , \pred_tab[2][CODE_ADR][30] , 
        \pred_tab[2][CODE_ADR][29] , \pred_tab[2][CODE_ADR][28] , 
        \pred_tab[2][CODE_ADR][27] , \pred_tab[2][CODE_ADR][26] , 
        \pred_tab[2][CODE_ADR][25] , \pred_tab[2][CODE_ADR][24] , 
        \pred_tab[2][CODE_ADR][23] , \pred_tab[2][CODE_ADR][22] , 
        \pred_tab[2][CODE_ADR][21] , \pred_tab[2][CODE_ADR][20] , 
        \pred_tab[2][CODE_ADR][19] , \pred_tab[2][CODE_ADR][18] , 
        \pred_tab[2][CODE_ADR][17] , \pred_tab[2][CODE_ADR][16] , 
        \pred_tab[2][CODE_ADR][15] , \pred_tab[2][CODE_ADR][14] , 
        \pred_tab[2][CODE_ADR][13] , \pred_tab[2][CODE_ADR][12] , 
        \pred_tab[2][CODE_ADR][11] , \pred_tab[2][CODE_ADR][10] , 
        \pred_tab[2][CODE_ADR][9] , \pred_tab[2][CODE_ADR][8] , 
        \pred_tab[2][CODE_ADR][7] , \pred_tab[2][CODE_ADR][6] , 
        \pred_tab[2][CODE_ADR][5] , \pred_tab[2][CODE_ADR][4] , 
        \pred_tab[2][CODE_ADR][3] , \pred_tab[2][CODE_ADR][2] , 
        \pred_tab[2][CODE_ADR][1] , \pred_tab[2][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N79) );
  predict_nb_record3_1_DW01_cmp6_6 eq_139_I2 ( .A(PF_pc), .B({
        \pred_tab[2][CODE_ADR][31] , \pred_tab[2][CODE_ADR][30] , 
        \pred_tab[2][CODE_ADR][29] , \pred_tab[2][CODE_ADR][28] , 
        \pred_tab[2][CODE_ADR][27] , \pred_tab[2][CODE_ADR][26] , 
        \pred_tab[2][CODE_ADR][25] , \pred_tab[2][CODE_ADR][24] , 
        \pred_tab[2][CODE_ADR][23] , \pred_tab[2][CODE_ADR][22] , 
        \pred_tab[2][CODE_ADR][21] , \pred_tab[2][CODE_ADR][20] , 
        \pred_tab[2][CODE_ADR][19] , \pred_tab[2][CODE_ADR][18] , 
        \pred_tab[2][CODE_ADR][17] , \pred_tab[2][CODE_ADR][16] , 
        \pred_tab[2][CODE_ADR][15] , \pred_tab[2][CODE_ADR][14] , 
        \pred_tab[2][CODE_ADR][13] , \pred_tab[2][CODE_ADR][12] , 
        \pred_tab[2][CODE_ADR][11] , \pred_tab[2][CODE_ADR][10] , 
        \pred_tab[2][CODE_ADR][9] , \pred_tab[2][CODE_ADR][8] , 
        \pred_tab[2][CODE_ADR][7] , \pred_tab[2][CODE_ADR][6] , 
        \pred_tab[2][CODE_ADR][5] , \pred_tab[2][CODE_ADR][4] , 
        \pred_tab[2][CODE_ADR][3] , \pred_tab[2][CODE_ADR][2] , 
        \pred_tab[2][CODE_ADR][1] , \pred_tab[2][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N76) );
  predict_nb_record3_1_DW01_cmp6_7 eq_145 ( .A(EX_adr), .B({
        \pred_tab[1][CODE_ADR][31] , \pred_tab[1][CODE_ADR][30] , 
        \pred_tab[1][CODE_ADR][29] , \pred_tab[1][CODE_ADR][28] , 
        \pred_tab[1][CODE_ADR][27] , \pred_tab[1][CODE_ADR][26] , 
        \pred_tab[1][CODE_ADR][25] , \pred_tab[1][CODE_ADR][24] , 
        \pred_tab[1][CODE_ADR][23] , \pred_tab[1][CODE_ADR][22] , 
        \pred_tab[1][CODE_ADR][21] , \pred_tab[1][CODE_ADR][20] , 
        \pred_tab[1][CODE_ADR][19] , \pred_tab[1][CODE_ADR][18] , 
        \pred_tab[1][CODE_ADR][17] , \pred_tab[1][CODE_ADR][16] , 
        \pred_tab[1][CODE_ADR][15] , \pred_tab[1][CODE_ADR][14] , 
        \pred_tab[1][CODE_ADR][13] , \pred_tab[1][CODE_ADR][12] , 
        \pred_tab[1][CODE_ADR][11] , \pred_tab[1][CODE_ADR][10] , 
        \pred_tab[1][CODE_ADR][9] , \pred_tab[1][CODE_ADR][8] , 
        \pred_tab[1][CODE_ADR][7] , \pred_tab[1][CODE_ADR][6] , 
        \pred_tab[1][CODE_ADR][5] , \pred_tab[1][CODE_ADR][4] , 
        \pred_tab[1][CODE_ADR][3] , \pred_tab[1][CODE_ADR][2] , 
        \pred_tab[1][CODE_ADR][1] , \pred_tab[1][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N71) );
  predict_nb_record3_1_DW01_cmp6_8 eq_142 ( .A(DI_adr), .B({
        \pred_tab[1][CODE_ADR][31] , \pred_tab[1][CODE_ADR][30] , 
        \pred_tab[1][CODE_ADR][29] , \pred_tab[1][CODE_ADR][28] , 
        \pred_tab[1][CODE_ADR][27] , \pred_tab[1][CODE_ADR][26] , 
        \pred_tab[1][CODE_ADR][25] , \pred_tab[1][CODE_ADR][24] , 
        \pred_tab[1][CODE_ADR][23] , \pred_tab[1][CODE_ADR][22] , 
        \pred_tab[1][CODE_ADR][21] , \pred_tab[1][CODE_ADR][20] , 
        \pred_tab[1][CODE_ADR][19] , \pred_tab[1][CODE_ADR][18] , 
        \pred_tab[1][CODE_ADR][17] , \pred_tab[1][CODE_ADR][16] , 
        \pred_tab[1][CODE_ADR][15] , \pred_tab[1][CODE_ADR][14] , 
        \pred_tab[1][CODE_ADR][13] , \pred_tab[1][CODE_ADR][12] , 
        \pred_tab[1][CODE_ADR][11] , \pred_tab[1][CODE_ADR][10] , 
        \pred_tab[1][CODE_ADR][9] , \pred_tab[1][CODE_ADR][8] , 
        \pred_tab[1][CODE_ADR][7] , \pred_tab[1][CODE_ADR][6] , 
        \pred_tab[1][CODE_ADR][5] , \pred_tab[1][CODE_ADR][4] , 
        \pred_tab[1][CODE_ADR][3] , \pred_tab[1][CODE_ADR][2] , 
        \pred_tab[1][CODE_ADR][1] , \pred_tab[1][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N70) );
  predict_nb_record3_1_DW01_cmp6_9 eq_139 ( .A(PF_pc), .B({
        \pred_tab[1][CODE_ADR][31] , \pred_tab[1][CODE_ADR][30] , 
        \pred_tab[1][CODE_ADR][29] , \pred_tab[1][CODE_ADR][28] , 
        \pred_tab[1][CODE_ADR][27] , \pred_tab[1][CODE_ADR][26] , 
        \pred_tab[1][CODE_ADR][25] , \pred_tab[1][CODE_ADR][24] , 
        \pred_tab[1][CODE_ADR][23] , \pred_tab[1][CODE_ADR][22] , 
        \pred_tab[1][CODE_ADR][21] , \pred_tab[1][CODE_ADR][20] , 
        \pred_tab[1][CODE_ADR][19] , \pred_tab[1][CODE_ADR][18] , 
        \pred_tab[1][CODE_ADR][17] , \pred_tab[1][CODE_ADR][16] , 
        \pred_tab[1][CODE_ADR][15] , \pred_tab[1][CODE_ADR][14] , 
        \pred_tab[1][CODE_ADR][13] , \pred_tab[1][CODE_ADR][12] , 
        \pred_tab[1][CODE_ADR][11] , \pred_tab[1][CODE_ADR][10] , 
        \pred_tab[1][CODE_ADR][9] , \pred_tab[1][CODE_ADR][8] , 
        \pred_tab[1][CODE_ADR][7] , \pred_tab[1][CODE_ADR][6] , 
        \pred_tab[1][CODE_ADR][5] , \pred_tab[1][CODE_ADR][4] , 
        \pred_tab[1][CODE_ADR][3] , \pred_tab[1][CODE_ADR][2] , 
        \pred_tab[1][CODE_ADR][1] , \pred_tab[1][CODE_ADR][0] }), .TC(1'b0), 
        .EQ(N69) );
  NAND_GATE U523 ( .I1(\next_out[0] ), .I2(N1582), .O(n13) );
  INV_GATE U621 ( .I1(n18), .O(n14) );
  INV_GATE U719 ( .I1(n18), .O(n15) );
  INV_GATE U721 ( .I1(n18), .O(n16) );
  INV_GATE U730 ( .I1(n18), .O(n17) );
  INV_GATE U1404 ( .I1(n294), .O(n18) );
  INV_GATE U1419 ( .I1(n23), .O(n19) );
  INV_GATE U1426 ( .I1(n23), .O(n20) );
  INV_GATE U1429 ( .I1(n23), .O(n21) );
  INV_GATE U1434 ( .I1(n23), .O(n22) );
  INV_GATE U1439 ( .I1(n163), .O(n23) );
  INV_GATE U1441 ( .I1(n427), .O(n24) );
  INV_GATE U1451 ( .I1(n427), .O(n25) );
  INV_GATE U1718 ( .I1(n427), .O(n26) );
  INV_GATE U1724 ( .I1(n427), .O(n27) );
  INV_GATE U1727 ( .I1(n36), .O(n427) );
  INV_GATE U1731 ( .I1(reset), .O(n434) );
  INV_GATE U1732 ( .I1(n28), .O(n447) );
  INV_GATE U1733 ( .I1(\next_out[0] ), .O(n512) );
  INV_GATE U1734 ( .I1(n29), .O(n577) );
  INV_GATE U1735 ( .I1(n441), .O(n642) );
  INV_GATE U1736 ( .I1(n647), .O(n646) );
  INV_GATE U1737 ( .I1(n1228), .O(PR_clear) );
  INV_GATE U1738 ( .I1(n1217), .O(n1223) );
  INV_GATE U1739 ( .I1(n1212), .O(n1227) );
  INV_GATE U1740 ( .I1(n1235), .O(n1229) );
  INV_GATE U1741 ( .I1(n1234), .O(n1233) );
  INV_GATE U1742 ( .I1(\next_out[1] ), .O(n1238) );
  AND_GATE U1743 ( .I1(N1582), .I2(\next_out[1] ), .O(N1614) );
endmodule


module bus_ctrl ( clock, reset, interrupt, adr_from_ei, instr_to_ei, 
        req_from_mem, r_w_from_mem, adr_from_mem, data_from_mem, data_to_mem, 
        req_to_ram, adr_to_ram, r_w_to_ram, ack_from_ram, data_inout_ram, 
        stop_all );
  input [31:0] adr_from_ei;
  output [31:0] instr_to_ei;
  input [31:0] adr_from_mem;
  input [31:0] data_from_mem;
  output [31:0] data_to_mem;
  output [31:0] adr_to_ram;
  inout [31:0] data_inout_ram;
  input clock, reset, interrupt, req_from_mem, r_w_from_mem, ack_from_ram;
  output req_to_ram, r_w_to_ram, stop_all;
  wire   cs, N46, req_allowed, n65, n67, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n1, n2,
         n3, n4, n5, n6;
  wire   [31:0] ei_buffer;
  tri   [31:0] data_inout_ram;

  FLIP_FLOP_D cs_reg ( .D(N46), .CK(clock), .Q(cs) );
  FLIP_FLOP_D \ei_buffer_reg[0]  ( .D(n237), .CK(clock), .Q(ei_buffer[0]) );
  FLIP_FLOP_D \ei_buffer_reg[10]  ( .D(n227), .CK(clock), .Q(ei_buffer[10]) );
  FLIP_FLOP_D \ei_buffer_reg[11]  ( .D(n226), .CK(clock), .Q(ei_buffer[11]) );
  FLIP_FLOP_D \ei_buffer_reg[12]  ( .D(n225), .CK(clock), .Q(ei_buffer[12]) );
  FLIP_FLOP_D \ei_buffer_reg[13]  ( .D(n224), .CK(clock), .Q(ei_buffer[13]) );
  FLIP_FLOP_D \ei_buffer_reg[14]  ( .D(n223), .CK(clock), .Q(ei_buffer[14]) );
  FLIP_FLOP_D \ei_buffer_reg[15]  ( .D(n222), .CK(clock), .Q(ei_buffer[15]) );
  FLIP_FLOP_D \ei_buffer_reg[16]  ( .D(n221), .CK(clock), .Q(ei_buffer[16]) );
  FLIP_FLOP_D \ei_buffer_reg[17]  ( .D(n220), .CK(clock), .Q(ei_buffer[17]) );
  FLIP_FLOP_D \ei_buffer_reg[18]  ( .D(n219), .CK(clock), .Q(ei_buffer[18]) );
  FLIP_FLOP_D \ei_buffer_reg[19]  ( .D(n218), .CK(clock), .Q(ei_buffer[19]) );
  FLIP_FLOP_D \ei_buffer_reg[1]  ( .D(n236), .CK(clock), .Q(ei_buffer[1]) );
  FLIP_FLOP_D \ei_buffer_reg[20]  ( .D(n217), .CK(clock), .Q(ei_buffer[20]) );
  FLIP_FLOP_D \ei_buffer_reg[21]  ( .D(n216), .CK(clock), .Q(ei_buffer[21]) );
  FLIP_FLOP_D \ei_buffer_reg[22]  ( .D(n215), .CK(clock), .Q(ei_buffer[22]) );
  FLIP_FLOP_D \ei_buffer_reg[23]  ( .D(n214), .CK(clock), .Q(ei_buffer[23]) );
  FLIP_FLOP_D \ei_buffer_reg[24]  ( .D(n213), .CK(clock), .Q(ei_buffer[24]) );
  FLIP_FLOP_D \ei_buffer_reg[25]  ( .D(n212), .CK(clock), .Q(ei_buffer[25]) );
  FLIP_FLOP_D \ei_buffer_reg[26]  ( .D(n211), .CK(clock), .Q(ei_buffer[26]) );
  FLIP_FLOP_D \ei_buffer_reg[27]  ( .D(n210), .CK(clock), .Q(ei_buffer[27]) );
  FLIP_FLOP_D \ei_buffer_reg[28]  ( .D(n209), .CK(clock), .Q(ei_buffer[28]) );
  FLIP_FLOP_D \ei_buffer_reg[29]  ( .D(n208), .CK(clock), .Q(ei_buffer[29]) );
  FLIP_FLOP_D \ei_buffer_reg[2]  ( .D(n235), .CK(clock), .Q(ei_buffer[2]) );
  FLIP_FLOP_D \ei_buffer_reg[30]  ( .D(n207), .CK(clock), .Q(ei_buffer[30]) );
  FLIP_FLOP_D \ei_buffer_reg[31]  ( .D(n206), .CK(clock), .Q(ei_buffer[31]) );
  FLIP_FLOP_D \ei_buffer_reg[3]  ( .D(n234), .CK(clock), .Q(ei_buffer[3]) );
  FLIP_FLOP_D \ei_buffer_reg[4]  ( .D(n233), .CK(clock), .Q(ei_buffer[4]) );
  FLIP_FLOP_D \ei_buffer_reg[5]  ( .D(n232), .CK(clock), .Q(ei_buffer[5]) );
  FLIP_FLOP_D \ei_buffer_reg[6]  ( .D(n231), .CK(clock), .Q(ei_buffer[6]) );
  FLIP_FLOP_D \ei_buffer_reg[7]  ( .D(n230), .CK(clock), .Q(ei_buffer[7]) );
  FLIP_FLOP_D \ei_buffer_reg[8]  ( .D(n229), .CK(clock), .Q(ei_buffer[8]) );
  FLIP_FLOP_D \ei_buffer_reg[9]  ( .D(n228), .CK(clock), .Q(ei_buffer[9]) );
  FLIP_FLOP_D_RESET req_allowed_reg ( .D(n205), .CK(clock), .RESET(
        ack_from_ram), .Q(req_allowed) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[0]  ( .I1(data_from_mem[0]), .E(n4), 
        .O(data_inout_ram[0]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[1]  ( .I1(data_from_mem[1]), .E(n4), 
        .O(data_inout_ram[1]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[2]  ( .I1(data_from_mem[2]), .E(n4), 
        .O(data_inout_ram[2]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[3]  ( .I1(data_from_mem[3]), .E(n4), 
        .O(data_inout_ram[3]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[4]  ( .I1(data_from_mem[4]), .E(n4), 
        .O(data_inout_ram[4]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[5]  ( .I1(data_from_mem[5]), .E(n4), 
        .O(data_inout_ram[5]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[6]  ( .I1(data_from_mem[6]), .E(n4), 
        .O(data_inout_ram[6]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[7]  ( .I1(data_from_mem[7]), .E(n4), 
        .O(data_inout_ram[7]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[8]  ( .I1(data_from_mem[8]), .E(n4), 
        .O(data_inout_ram[8]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[9]  ( .I1(data_from_mem[9]), .E(n4), 
        .O(data_inout_ram[9]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[10]  ( .I1(data_from_mem[10]), .E(
        n4), .O(data_inout_ram[10]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[11]  ( .I1(data_from_mem[11]), .E(
        n4), .O(data_inout_ram[11]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[12]  ( .I1(data_from_mem[12]), .E(
        n4), .O(data_inout_ram[12]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[13]  ( .I1(data_from_mem[13]), .E(
        n4), .O(data_inout_ram[13]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[14]  ( .I1(data_from_mem[14]), .E(
        n4), .O(data_inout_ram[14]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[15]  ( .I1(data_from_mem[15]), .E(
        n4), .O(data_inout_ram[15]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[16]  ( .I1(data_from_mem[16]), .E(
        n4), .O(data_inout_ram[16]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[17]  ( .I1(data_from_mem[17]), .E(
        n4), .O(data_inout_ram[17]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[18]  ( .I1(data_from_mem[18]), .E(
        n4), .O(data_inout_ram[18]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[19]  ( .I1(data_from_mem[19]), .E(
        n4), .O(data_inout_ram[19]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[20]  ( .I1(data_from_mem[20]), .E(
        n4), .O(data_inout_ram[20]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[21]  ( .I1(data_from_mem[21]), .E(
        n4), .O(data_inout_ram[21]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[22]  ( .I1(data_from_mem[22]), .E(
        n4), .O(data_inout_ram[22]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[23]  ( .I1(data_from_mem[23]), .E(
        n4), .O(data_inout_ram[23]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[24]  ( .I1(data_from_mem[24]), .E(
        n4), .O(data_inout_ram[24]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[25]  ( .I1(data_from_mem[25]), .E(
        n4), .O(data_inout_ram[25]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[26]  ( .I1(data_from_mem[26]), .E(
        n4), .O(data_inout_ram[26]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[27]  ( .I1(data_from_mem[27]), .E(
        n4), .O(data_inout_ram[27]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[28]  ( .I1(data_from_mem[28]), .E(
        n4), .O(data_inout_ram[28]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[29]  ( .I1(data_from_mem[29]), .E(
        n4), .O(data_inout_ram[29]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[30]  ( .I1(data_from_mem[30]), .E(
        n4), .O(data_inout_ram[30]) );
  THREE_STATE_BUF_GATE \data_inout_ram_tri[31]  ( .I1(data_from_mem[31]), .E(
        n4), .O(data_inout_ram[31]) );
  AND_GATE U3 ( .I1(n65), .I2(n5), .O(stop_all) );
  NAND_GATE U4 ( .I1(ack_from_ram), .I2(n67), .O(n65) );
  NAND_GATE U5 ( .I1(req_from_mem), .I2(n2), .O(n67) );
  OR_GATE U6 ( .I1(n6), .I2(req_allowed), .O(req_to_ram) );
  OR_GATE U7 ( .I1(ack_from_ram), .I2(req_allowed), .O(n205) );
  AND_GATE U8 ( .I1(instr_to_ei[31]), .I2(n3), .O(n206) );
  AND_GATE U9 ( .I1(instr_to_ei[30]), .I2(n3), .O(n207) );
  AND_GATE U10 ( .I1(instr_to_ei[29]), .I2(n3), .O(n208) );
  AND_GATE U11 ( .I1(instr_to_ei[28]), .I2(n3), .O(n209) );
  AND_GATE U12 ( .I1(instr_to_ei[27]), .I2(n3), .O(n210) );
  AND_GATE U13 ( .I1(instr_to_ei[26]), .I2(n3), .O(n211) );
  AND_GATE U14 ( .I1(instr_to_ei[25]), .I2(n3), .O(n212) );
  AND_GATE U15 ( .I1(instr_to_ei[24]), .I2(n3), .O(n213) );
  AND_GATE U16 ( .I1(instr_to_ei[23]), .I2(n3), .O(n214) );
  AND_GATE U17 ( .I1(instr_to_ei[22]), .I2(n3), .O(n215) );
  AND_GATE U18 ( .I1(instr_to_ei[21]), .I2(n3), .O(n216) );
  AND_GATE U19 ( .I1(instr_to_ei[20]), .I2(n3), .O(n217) );
  AND_GATE U20 ( .I1(instr_to_ei[19]), .I2(n3), .O(n218) );
  AND_GATE U21 ( .I1(instr_to_ei[18]), .I2(n3), .O(n219) );
  AND_GATE U22 ( .I1(instr_to_ei[17]), .I2(n3), .O(n220) );
  AND_GATE U23 ( .I1(instr_to_ei[16]), .I2(n3), .O(n221) );
  AND_GATE U24 ( .I1(instr_to_ei[15]), .I2(n3), .O(n222) );
  AND_GATE U25 ( .I1(instr_to_ei[14]), .I2(n3), .O(n223) );
  AND_GATE U26 ( .I1(instr_to_ei[13]), .I2(n3), .O(n224) );
  AND_GATE U27 ( .I1(instr_to_ei[12]), .I2(n3), .O(n225) );
  AND_GATE U28 ( .I1(instr_to_ei[11]), .I2(n3), .O(n226) );
  AND_GATE U29 ( .I1(instr_to_ei[10]), .I2(n3), .O(n227) );
  AND_GATE U30 ( .I1(instr_to_ei[9]), .I2(n3), .O(n228) );
  AND_GATE U31 ( .I1(instr_to_ei[8]), .I2(n3), .O(n229) );
  AND_GATE U32 ( .I1(instr_to_ei[7]), .I2(n3), .O(n230) );
  AND_GATE U33 ( .I1(instr_to_ei[6]), .I2(n3), .O(n231) );
  AND_GATE U34 ( .I1(instr_to_ei[5]), .I2(n3), .O(n232) );
  AND_GATE U35 ( .I1(instr_to_ei[4]), .I2(n3), .O(n233) );
  AND_GATE U36 ( .I1(instr_to_ei[3]), .I2(n3), .O(n234) );
  AND_GATE U37 ( .I1(instr_to_ei[2]), .I2(n3), .O(n235) );
  AND_GATE U38 ( .I1(instr_to_ei[1]), .I2(n3), .O(n236) );
  AND_GATE U39 ( .I1(instr_to_ei[0]), .I2(n3), .O(n237) );
  NAND_GATE U40 ( .I1(n71), .I2(n72), .O(instr_to_ei[9]) );
  NAND_GATE U41 ( .I1(data_to_mem[9]), .I2(n2), .O(n72) );
  NAND_GATE U42 ( .I1(ei_buffer[9]), .I2(cs), .O(n71) );
  NAND_GATE U43 ( .I1(n73), .I2(n74), .O(instr_to_ei[8]) );
  NAND_GATE U44 ( .I1(data_to_mem[8]), .I2(n2), .O(n74) );
  NAND_GATE U45 ( .I1(ei_buffer[8]), .I2(cs), .O(n73) );
  NAND_GATE U46 ( .I1(n75), .I2(n76), .O(instr_to_ei[7]) );
  NAND_GATE U47 ( .I1(data_to_mem[7]), .I2(n2), .O(n76) );
  NAND_GATE U48 ( .I1(ei_buffer[7]), .I2(cs), .O(n75) );
  NAND_GATE U49 ( .I1(n77), .I2(n78), .O(instr_to_ei[6]) );
  NAND_GATE U50 ( .I1(data_to_mem[6]), .I2(n2), .O(n78) );
  NAND_GATE U51 ( .I1(ei_buffer[6]), .I2(cs), .O(n77) );
  NAND_GATE U52 ( .I1(n79), .I2(n80), .O(instr_to_ei[5]) );
  NAND_GATE U53 ( .I1(data_to_mem[5]), .I2(n2), .O(n80) );
  NAND_GATE U54 ( .I1(ei_buffer[5]), .I2(cs), .O(n79) );
  NAND_GATE U55 ( .I1(n81), .I2(n82), .O(instr_to_ei[4]) );
  NAND_GATE U56 ( .I1(data_to_mem[4]), .I2(n2), .O(n82) );
  NAND_GATE U57 ( .I1(ei_buffer[4]), .I2(cs), .O(n81) );
  NAND_GATE U58 ( .I1(n83), .I2(n84), .O(instr_to_ei[3]) );
  NAND_GATE U59 ( .I1(data_to_mem[3]), .I2(n2), .O(n84) );
  NAND_GATE U60 ( .I1(ei_buffer[3]), .I2(cs), .O(n83) );
  NAND_GATE U61 ( .I1(n85), .I2(n86), .O(instr_to_ei[31]) );
  NAND_GATE U62 ( .I1(data_to_mem[31]), .I2(n2), .O(n86) );
  NAND_GATE U63 ( .I1(ei_buffer[31]), .I2(cs), .O(n85) );
  NAND_GATE U64 ( .I1(n87), .I2(n88), .O(instr_to_ei[30]) );
  NAND_GATE U65 ( .I1(data_to_mem[30]), .I2(n2), .O(n88) );
  NAND_GATE U66 ( .I1(ei_buffer[30]), .I2(cs), .O(n87) );
  NAND_GATE U67 ( .I1(n89), .I2(n90), .O(instr_to_ei[2]) );
  NAND_GATE U68 ( .I1(data_to_mem[2]), .I2(n2), .O(n90) );
  NAND_GATE U69 ( .I1(ei_buffer[2]), .I2(cs), .O(n89) );
  NAND_GATE U70 ( .I1(n91), .I2(n92), .O(instr_to_ei[29]) );
  NAND_GATE U71 ( .I1(data_to_mem[29]), .I2(n2), .O(n92) );
  NAND_GATE U72 ( .I1(ei_buffer[29]), .I2(cs), .O(n91) );
  NAND_GATE U73 ( .I1(n93), .I2(n94), .O(instr_to_ei[28]) );
  NAND_GATE U74 ( .I1(data_to_mem[28]), .I2(n2), .O(n94) );
  NAND_GATE U75 ( .I1(ei_buffer[28]), .I2(cs), .O(n93) );
  NAND_GATE U76 ( .I1(n95), .I2(n96), .O(instr_to_ei[27]) );
  NAND_GATE U77 ( .I1(data_to_mem[27]), .I2(n2), .O(n96) );
  NAND_GATE U78 ( .I1(ei_buffer[27]), .I2(cs), .O(n95) );
  NAND_GATE U79 ( .I1(n97), .I2(n98), .O(instr_to_ei[26]) );
  NAND_GATE U80 ( .I1(data_to_mem[26]), .I2(n2), .O(n98) );
  NAND_GATE U81 ( .I1(ei_buffer[26]), .I2(cs), .O(n97) );
  NAND_GATE U82 ( .I1(n99), .I2(n100), .O(instr_to_ei[25]) );
  NAND_GATE U83 ( .I1(data_to_mem[25]), .I2(n2), .O(n100) );
  NAND_GATE U84 ( .I1(ei_buffer[25]), .I2(cs), .O(n99) );
  NAND_GATE U85 ( .I1(n101), .I2(n102), .O(instr_to_ei[24]) );
  NAND_GATE U86 ( .I1(data_to_mem[24]), .I2(n2), .O(n102) );
  NAND_GATE U87 ( .I1(ei_buffer[24]), .I2(cs), .O(n101) );
  NAND_GATE U88 ( .I1(n103), .I2(n104), .O(instr_to_ei[23]) );
  NAND_GATE U89 ( .I1(data_to_mem[23]), .I2(n2), .O(n104) );
  NAND_GATE U90 ( .I1(ei_buffer[23]), .I2(cs), .O(n103) );
  NAND_GATE U91 ( .I1(n105), .I2(n106), .O(instr_to_ei[22]) );
  NAND_GATE U92 ( .I1(data_to_mem[22]), .I2(n2), .O(n106) );
  NAND_GATE U93 ( .I1(ei_buffer[22]), .I2(cs), .O(n105) );
  NAND_GATE U94 ( .I1(n107), .I2(n108), .O(instr_to_ei[21]) );
  NAND_GATE U95 ( .I1(data_to_mem[21]), .I2(n2), .O(n108) );
  NAND_GATE U96 ( .I1(ei_buffer[21]), .I2(cs), .O(n107) );
  NAND_GATE U97 ( .I1(n109), .I2(n110), .O(instr_to_ei[20]) );
  NAND_GATE U98 ( .I1(data_to_mem[20]), .I2(n2), .O(n110) );
  NAND_GATE U99 ( .I1(ei_buffer[20]), .I2(cs), .O(n109) );
  NAND_GATE U100 ( .I1(n111), .I2(n112), .O(instr_to_ei[1]) );
  NAND_GATE U101 ( .I1(data_to_mem[1]), .I2(n2), .O(n112) );
  NAND_GATE U102 ( .I1(ei_buffer[1]), .I2(cs), .O(n111) );
  NAND_GATE U103 ( .I1(n113), .I2(n114), .O(instr_to_ei[19]) );
  NAND_GATE U104 ( .I1(data_to_mem[19]), .I2(n2), .O(n114) );
  NAND_GATE U105 ( .I1(ei_buffer[19]), .I2(cs), .O(n113) );
  NAND_GATE U106 ( .I1(n115), .I2(n116), .O(instr_to_ei[18]) );
  NAND_GATE U107 ( .I1(data_to_mem[18]), .I2(n2), .O(n116) );
  NAND_GATE U108 ( .I1(ei_buffer[18]), .I2(cs), .O(n115) );
  NAND_GATE U109 ( .I1(n117), .I2(n118), .O(instr_to_ei[17]) );
  NAND_GATE U110 ( .I1(data_to_mem[17]), .I2(n2), .O(n118) );
  NAND_GATE U111 ( .I1(ei_buffer[17]), .I2(cs), .O(n117) );
  NAND_GATE U112 ( .I1(n119), .I2(n120), .O(instr_to_ei[16]) );
  NAND_GATE U113 ( .I1(data_to_mem[16]), .I2(n2), .O(n120) );
  NAND_GATE U114 ( .I1(ei_buffer[16]), .I2(cs), .O(n119) );
  NAND_GATE U115 ( .I1(n121), .I2(n122), .O(instr_to_ei[15]) );
  NAND_GATE U116 ( .I1(data_to_mem[15]), .I2(n2), .O(n122) );
  NAND_GATE U117 ( .I1(ei_buffer[15]), .I2(cs), .O(n121) );
  NAND_GATE U118 ( .I1(n123), .I2(n124), .O(instr_to_ei[14]) );
  NAND_GATE U119 ( .I1(data_to_mem[14]), .I2(n2), .O(n124) );
  NAND_GATE U120 ( .I1(ei_buffer[14]), .I2(cs), .O(n123) );
  NAND_GATE U121 ( .I1(n125), .I2(n126), .O(instr_to_ei[13]) );
  NAND_GATE U122 ( .I1(data_to_mem[13]), .I2(n2), .O(n126) );
  NAND_GATE U123 ( .I1(ei_buffer[13]), .I2(cs), .O(n125) );
  NAND_GATE U124 ( .I1(n127), .I2(n128), .O(instr_to_ei[12]) );
  NAND_GATE U125 ( .I1(data_to_mem[12]), .I2(n2), .O(n128) );
  NAND_GATE U126 ( .I1(ei_buffer[12]), .I2(cs), .O(n127) );
  NAND_GATE U127 ( .I1(n129), .I2(n130), .O(instr_to_ei[11]) );
  NAND_GATE U128 ( .I1(data_to_mem[11]), .I2(n2), .O(n130) );
  NAND_GATE U129 ( .I1(ei_buffer[11]), .I2(cs), .O(n129) );
  NAND_GATE U130 ( .I1(n131), .I2(n132), .O(instr_to_ei[10]) );
  NAND_GATE U131 ( .I1(data_to_mem[10]), .I2(n2), .O(n132) );
  NAND_GATE U132 ( .I1(ei_buffer[10]), .I2(cs), .O(n131) );
  NAND_GATE U133 ( .I1(n133), .I2(n134), .O(instr_to_ei[0]) );
  NAND_GATE U134 ( .I1(data_to_mem[0]), .I2(n2), .O(n134) );
  NAND_GATE U135 ( .I1(ei_buffer[0]), .I2(cs), .O(n133) );
  AND_GATE U136 ( .I1(data_inout_ram[9]), .I2(n4), .O(data_to_mem[9]) );
  AND_GATE U137 ( .I1(data_inout_ram[8]), .I2(n4), .O(data_to_mem[8]) );
  AND_GATE U138 ( .I1(data_inout_ram[7]), .I2(n4), .O(data_to_mem[7]) );
  AND_GATE U139 ( .I1(data_inout_ram[6]), .I2(n4), .O(data_to_mem[6]) );
  AND_GATE U140 ( .I1(data_inout_ram[5]), .I2(n4), .O(data_to_mem[5]) );
  AND_GATE U141 ( .I1(data_inout_ram[4]), .I2(n4), .O(data_to_mem[4]) );
  AND_GATE U142 ( .I1(data_inout_ram[3]), .I2(n4), .O(data_to_mem[3]) );
  AND_GATE U143 ( .I1(data_inout_ram[31]), .I2(n4), .O(data_to_mem[31]) );
  AND_GATE U144 ( .I1(data_inout_ram[30]), .I2(n4), .O(data_to_mem[30]) );
  AND_GATE U145 ( .I1(data_inout_ram[2]), .I2(n4), .O(data_to_mem[2]) );
  AND_GATE U146 ( .I1(data_inout_ram[29]), .I2(n4), .O(data_to_mem[29]) );
  AND_GATE U147 ( .I1(data_inout_ram[28]), .I2(n4), .O(data_to_mem[28]) );
  AND_GATE U148 ( .I1(data_inout_ram[27]), .I2(n4), .O(data_to_mem[27]) );
  AND_GATE U149 ( .I1(data_inout_ram[26]), .I2(n4), .O(data_to_mem[26]) );
  AND_GATE U150 ( .I1(data_inout_ram[25]), .I2(n4), .O(data_to_mem[25]) );
  AND_GATE U151 ( .I1(data_inout_ram[24]), .I2(n4), .O(data_to_mem[24]) );
  AND_GATE U152 ( .I1(data_inout_ram[23]), .I2(n4), .O(data_to_mem[23]) );
  AND_GATE U153 ( .I1(data_inout_ram[22]), .I2(n4), .O(data_to_mem[22]) );
  AND_GATE U154 ( .I1(data_inout_ram[21]), .I2(n4), .O(data_to_mem[21]) );
  AND_GATE U155 ( .I1(data_inout_ram[20]), .I2(n4), .O(data_to_mem[20]) );
  AND_GATE U156 ( .I1(data_inout_ram[1]), .I2(n4), .O(data_to_mem[1]) );
  AND_GATE U157 ( .I1(data_inout_ram[19]), .I2(n4), .O(data_to_mem[19]) );
  AND_GATE U158 ( .I1(data_inout_ram[18]), .I2(n4), .O(data_to_mem[18]) );
  AND_GATE U159 ( .I1(data_inout_ram[17]), .I2(n4), .O(data_to_mem[17]) );
  AND_GATE U160 ( .I1(data_inout_ram[16]), .I2(n4), .O(data_to_mem[16]) );
  AND_GATE U161 ( .I1(data_inout_ram[15]), .I2(n4), .O(data_to_mem[15]) );
  AND_GATE U162 ( .I1(data_inout_ram[14]), .I2(n4), .O(data_to_mem[14]) );
  AND_GATE U163 ( .I1(data_inout_ram[13]), .I2(n4), .O(data_to_mem[13]) );
  AND_GATE U164 ( .I1(data_inout_ram[12]), .I2(n4), .O(data_to_mem[12]) );
  AND_GATE U165 ( .I1(data_inout_ram[11]), .I2(n4), .O(data_to_mem[11]) );
  AND_GATE U166 ( .I1(data_inout_ram[10]), .I2(n4), .O(data_to_mem[10]) );
  AND_GATE U167 ( .I1(data_inout_ram[0]), .I2(n4), .O(data_to_mem[0]) );
  AND_GATE U169 ( .I1(r_w_from_mem), .I2(n135), .O(r_w_to_ram) );
  NAND_GATE U170 ( .I1(n136), .I2(n137), .O(adr_to_ram[9]) );
  NAND_GATE U171 ( .I1(adr_from_ei[9]), .I2(n1), .O(n137) );
  NAND_GATE U172 ( .I1(adr_from_mem[9]), .I2(n135), .O(n136) );
  NAND_GATE U173 ( .I1(n139), .I2(n140), .O(adr_to_ram[8]) );
  NAND_GATE U174 ( .I1(adr_from_ei[8]), .I2(n1), .O(n140) );
  NAND_GATE U175 ( .I1(adr_from_mem[8]), .I2(n135), .O(n139) );
  NAND_GATE U176 ( .I1(n141), .I2(n142), .O(adr_to_ram[7]) );
  NAND_GATE U177 ( .I1(adr_from_ei[7]), .I2(n1), .O(n142) );
  NAND_GATE U178 ( .I1(adr_from_mem[7]), .I2(n135), .O(n141) );
  NAND_GATE U179 ( .I1(n143), .I2(n144), .O(adr_to_ram[6]) );
  NAND_GATE U180 ( .I1(adr_from_ei[6]), .I2(n1), .O(n144) );
  NAND_GATE U181 ( .I1(adr_from_mem[6]), .I2(n135), .O(n143) );
  NAND_GATE U182 ( .I1(n145), .I2(n146), .O(adr_to_ram[5]) );
  NAND_GATE U183 ( .I1(adr_from_ei[5]), .I2(n1), .O(n146) );
  NAND_GATE U184 ( .I1(adr_from_mem[5]), .I2(n135), .O(n145) );
  NAND_GATE U185 ( .I1(n147), .I2(n148), .O(adr_to_ram[4]) );
  NAND_GATE U186 ( .I1(adr_from_ei[4]), .I2(n1), .O(n148) );
  NAND_GATE U187 ( .I1(adr_from_mem[4]), .I2(n135), .O(n147) );
  NAND_GATE U188 ( .I1(n149), .I2(n150), .O(adr_to_ram[3]) );
  NAND_GATE U189 ( .I1(adr_from_ei[3]), .I2(n1), .O(n150) );
  NAND_GATE U190 ( .I1(adr_from_mem[3]), .I2(n135), .O(n149) );
  NAND_GATE U191 ( .I1(n151), .I2(n152), .O(adr_to_ram[31]) );
  NAND_GATE U192 ( .I1(adr_from_ei[31]), .I2(n1), .O(n152) );
  NAND_GATE U193 ( .I1(adr_from_mem[31]), .I2(n135), .O(n151) );
  NAND_GATE U194 ( .I1(n153), .I2(n154), .O(adr_to_ram[30]) );
  NAND_GATE U195 ( .I1(adr_from_ei[30]), .I2(n1), .O(n154) );
  NAND_GATE U196 ( .I1(adr_from_mem[30]), .I2(n135), .O(n153) );
  NAND_GATE U197 ( .I1(n155), .I2(n156), .O(adr_to_ram[2]) );
  NAND_GATE U198 ( .I1(adr_from_ei[2]), .I2(n1), .O(n156) );
  NAND_GATE U199 ( .I1(adr_from_mem[2]), .I2(n135), .O(n155) );
  NAND_GATE U200 ( .I1(n157), .I2(n158), .O(adr_to_ram[29]) );
  NAND_GATE U201 ( .I1(adr_from_ei[29]), .I2(n1), .O(n158) );
  NAND_GATE U202 ( .I1(adr_from_mem[29]), .I2(n135), .O(n157) );
  NAND_GATE U203 ( .I1(n159), .I2(n160), .O(adr_to_ram[28]) );
  NAND_GATE U204 ( .I1(adr_from_ei[28]), .I2(n1), .O(n160) );
  NAND_GATE U205 ( .I1(adr_from_mem[28]), .I2(n135), .O(n159) );
  NAND_GATE U206 ( .I1(n161), .I2(n162), .O(adr_to_ram[27]) );
  NAND_GATE U207 ( .I1(adr_from_ei[27]), .I2(n1), .O(n162) );
  NAND_GATE U208 ( .I1(adr_from_mem[27]), .I2(n135), .O(n161) );
  NAND_GATE U209 ( .I1(n163), .I2(n164), .O(adr_to_ram[26]) );
  NAND_GATE U210 ( .I1(adr_from_ei[26]), .I2(n1), .O(n164) );
  NAND_GATE U211 ( .I1(adr_from_mem[26]), .I2(n135), .O(n163) );
  NAND_GATE U212 ( .I1(n165), .I2(n166), .O(adr_to_ram[25]) );
  NAND_GATE U213 ( .I1(adr_from_ei[25]), .I2(n1), .O(n166) );
  NAND_GATE U214 ( .I1(adr_from_mem[25]), .I2(n135), .O(n165) );
  NAND_GATE U215 ( .I1(n167), .I2(n168), .O(adr_to_ram[24]) );
  NAND_GATE U216 ( .I1(adr_from_ei[24]), .I2(n1), .O(n168) );
  NAND_GATE U217 ( .I1(adr_from_mem[24]), .I2(n135), .O(n167) );
  NAND_GATE U218 ( .I1(n169), .I2(n170), .O(adr_to_ram[23]) );
  NAND_GATE U219 ( .I1(adr_from_ei[23]), .I2(n1), .O(n170) );
  NAND_GATE U220 ( .I1(adr_from_mem[23]), .I2(n135), .O(n169) );
  NAND_GATE U221 ( .I1(n171), .I2(n172), .O(adr_to_ram[22]) );
  NAND_GATE U222 ( .I1(adr_from_ei[22]), .I2(n1), .O(n172) );
  NAND_GATE U223 ( .I1(adr_from_mem[22]), .I2(n135), .O(n171) );
  NAND_GATE U224 ( .I1(n173), .I2(n174), .O(adr_to_ram[21]) );
  NAND_GATE U225 ( .I1(adr_from_ei[21]), .I2(n1), .O(n174) );
  NAND_GATE U226 ( .I1(adr_from_mem[21]), .I2(n135), .O(n173) );
  NAND_GATE U227 ( .I1(n175), .I2(n176), .O(adr_to_ram[20]) );
  NAND_GATE U228 ( .I1(adr_from_ei[20]), .I2(n1), .O(n176) );
  NAND_GATE U229 ( .I1(adr_from_mem[20]), .I2(n135), .O(n175) );
  NAND_GATE U230 ( .I1(n177), .I2(n178), .O(adr_to_ram[1]) );
  NAND_GATE U231 ( .I1(adr_from_ei[1]), .I2(n1), .O(n178) );
  NAND_GATE U232 ( .I1(adr_from_mem[1]), .I2(n135), .O(n177) );
  NAND_GATE U233 ( .I1(n179), .I2(n180), .O(adr_to_ram[19]) );
  NAND_GATE U234 ( .I1(adr_from_ei[19]), .I2(n1), .O(n180) );
  NAND_GATE U235 ( .I1(adr_from_mem[19]), .I2(n135), .O(n179) );
  NAND_GATE U236 ( .I1(n181), .I2(n182), .O(adr_to_ram[18]) );
  NAND_GATE U237 ( .I1(adr_from_ei[18]), .I2(n1), .O(n182) );
  NAND_GATE U238 ( .I1(adr_from_mem[18]), .I2(n135), .O(n181) );
  NAND_GATE U239 ( .I1(n183), .I2(n184), .O(adr_to_ram[17]) );
  NAND_GATE U240 ( .I1(adr_from_ei[17]), .I2(n1), .O(n184) );
  NAND_GATE U241 ( .I1(adr_from_mem[17]), .I2(n135), .O(n183) );
  NAND_GATE U242 ( .I1(n185), .I2(n186), .O(adr_to_ram[16]) );
  NAND_GATE U243 ( .I1(adr_from_ei[16]), .I2(n1), .O(n186) );
  NAND_GATE U244 ( .I1(adr_from_mem[16]), .I2(n135), .O(n185) );
  NAND_GATE U245 ( .I1(n187), .I2(n188), .O(adr_to_ram[15]) );
  NAND_GATE U246 ( .I1(adr_from_ei[15]), .I2(n1), .O(n188) );
  NAND_GATE U247 ( .I1(adr_from_mem[15]), .I2(n135), .O(n187) );
  NAND_GATE U248 ( .I1(n189), .I2(n190), .O(adr_to_ram[14]) );
  NAND_GATE U249 ( .I1(adr_from_ei[14]), .I2(n1), .O(n190) );
  NAND_GATE U250 ( .I1(adr_from_mem[14]), .I2(n135), .O(n189) );
  NAND_GATE U251 ( .I1(n191), .I2(n192), .O(adr_to_ram[13]) );
  NAND_GATE U252 ( .I1(adr_from_ei[13]), .I2(n1), .O(n192) );
  NAND_GATE U253 ( .I1(adr_from_mem[13]), .I2(n135), .O(n191) );
  NAND_GATE U254 ( .I1(n193), .I2(n194), .O(adr_to_ram[12]) );
  NAND_GATE U255 ( .I1(adr_from_ei[12]), .I2(n1), .O(n194) );
  NAND_GATE U256 ( .I1(adr_from_mem[12]), .I2(n135), .O(n193) );
  NAND_GATE U257 ( .I1(n195), .I2(n196), .O(adr_to_ram[11]) );
  NAND_GATE U258 ( .I1(adr_from_ei[11]), .I2(n1), .O(n196) );
  NAND_GATE U259 ( .I1(adr_from_mem[11]), .I2(n135), .O(n195) );
  NAND_GATE U260 ( .I1(n197), .I2(n198), .O(adr_to_ram[10]) );
  NAND_GATE U261 ( .I1(adr_from_ei[10]), .I2(n1), .O(n198) );
  NAND_GATE U262 ( .I1(adr_from_mem[10]), .I2(n135), .O(n197) );
  NAND_GATE U263 ( .I1(n199), .I2(n200), .O(adr_to_ram[0]) );
  NAND_GATE U264 ( .I1(adr_from_ei[0]), .I2(n1), .O(n200) );
  NAND_GATE U266 ( .I1(adr_from_mem[0]), .I2(n135), .O(n199) );
  AND_GATE U267 ( .I1(n201), .I2(n3), .O(N46) );
  NAND_GATE U269 ( .I1(n202), .I2(n203), .O(n201) );
  NAND4_GATE U270 ( .I1(ack_from_ram), .I2(req_from_mem), .I3(n2), .I4(n5), 
        .O(n203) );
  NAND_GATE U272 ( .I1(n135), .I2(n6), .O(n202) );
  NOR_GATE U274 ( .I1(n2), .I2(interrupt), .O(n135) );
  INV_GATE U168 ( .I1(n135), .O(n1) );
  INV_GATE U265 ( .I1(cs), .O(n2) );
  INV_GATE U268 ( .I1(reset), .O(n3) );
  INV_GATE U271 ( .I1(r_w_to_ram), .O(n4) );
  INV_GATE U273 ( .I1(interrupt), .O(n5) );
  INV_GATE U275 ( .I1(ack_from_ram), .O(n6) );
endmodule


module syscop ( clock, reset, MEM_adr, MEM_exc_cause, MEM_it_ok, it_mat, 
        interrupt, vecteur_it, write_data, write_adr, write_SCP, read_adr1, 
        read_adr2, read_data1, read_data2 );
  input [31:0] MEM_adr;
  input [31:0] MEM_exc_cause;
  output [31:0] vecteur_it;
  input [31:0] write_data;
  input [4:0] write_adr;
  input [4:0] read_adr1;
  input [4:0] read_adr2;
  output [31:0] read_data1;
  output [31:0] read_data2;
  input clock, reset, MEM_it_ok, it_mat, write_SCP;
  output interrupt;
  wire   \scp_reg[12][31] , \scp_reg[12][30] , \scp_reg[12][29] ,
         \scp_reg[12][28] , \scp_reg[12][27] , \scp_reg[12][26] ,
         \scp_reg[12][25] , \scp_reg[12][24] , \scp_reg[12][23] ,
         \scp_reg[12][22] , \scp_reg[12][21] , \scp_reg[12][20] ,
         \scp_reg[12][19] , \scp_reg[12][18] , \scp_reg[12][17] ,
         \scp_reg[12][16] , \scp_reg[12][15] , \scp_reg[12][14] ,
         \scp_reg[12][13] , \scp_reg[12][12] , \scp_reg[12][11] ,
         \scp_reg[12][10] , \scp_reg[12][9] , \scp_reg[12][8] ,
         \scp_reg[12][7] , \scp_reg[12][6] , \scp_reg[12][5] ,
         \scp_reg[12][4] , \scp_reg[12][3] , \scp_reg[12][2] ,
         \scp_reg[12][1] , \scp_reg[12][0] , \scp_reg[13][31] ,
         \scp_reg[13][30] , \scp_reg[13][29] , \scp_reg[13][28] ,
         \scp_reg[13][27] , \scp_reg[13][26] , \scp_reg[13][25] ,
         \scp_reg[13][24] , \scp_reg[13][23] , \scp_reg[13][22] ,
         \scp_reg[13][21] , \scp_reg[13][20] , \scp_reg[13][19] ,
         \scp_reg[13][18] , \scp_reg[13][17] , \scp_reg[13][16] ,
         \scp_reg[13][15] , \scp_reg[13][14] , \scp_reg[13][13] ,
         \scp_reg[13][12] , \scp_reg[13][11] , \scp_reg[13][10] ,
         \scp_reg[13][9] , \scp_reg[13][8] , \scp_reg[13][7] ,
         \scp_reg[13][6] , \scp_reg[13][5] , \scp_reg[13][4] ,
         \scp_reg[13][3] , \scp_reg[13][2] , \scp_reg[13][1] ,
         \scp_reg[13][0] , \scp_reg[14][31] , \scp_reg[14][30] ,
         \scp_reg[14][29] , \scp_reg[14][28] , \scp_reg[14][27] ,
         \scp_reg[14][26] , \scp_reg[14][25] , \scp_reg[14][24] ,
         \scp_reg[14][23] , \scp_reg[14][22] , \scp_reg[14][21] ,
         \scp_reg[14][20] , \scp_reg[14][19] , \scp_reg[14][18] ,
         \scp_reg[14][17] , \scp_reg[14][16] , \scp_reg[14][15] ,
         \scp_reg[14][14] , \scp_reg[14][13] , \scp_reg[14][12] ,
         \scp_reg[14][11] , \scp_reg[14][10] , \scp_reg[14][9] ,
         \scp_reg[14][8] , \scp_reg[14][7] , \scp_reg[14][6] ,
         \scp_reg[14][5] , \scp_reg[14][4] , \scp_reg[14][3] ,
         \scp_reg[14][2] , \scp_reg[14][1] , \scp_reg[14][0] ,
         \scp_reg[15][31] , \scp_reg[15][30] , \scp_reg[15][29] ,
         \scp_reg[15][28] , \scp_reg[15][27] , \scp_reg[15][26] ,
         \scp_reg[15][25] , \scp_reg[15][24] , \scp_reg[15][23] ,
         \scp_reg[15][22] , \scp_reg[15][21] , \scp_reg[15][20] ,
         \scp_reg[15][19] , \scp_reg[15][18] , \scp_reg[15][17] ,
         \scp_reg[15][16] , \scp_reg[15][15] , \scp_reg[15][14] ,
         \scp_reg[15][13] , \scp_reg[15][12] , \scp_reg[15][11] ,
         \scp_reg[15][10] , \scp_reg[15][9] , \scp_reg[15][8] ,
         \scp_reg[15][7] , \scp_reg[15][6] , \scp_reg[15][5] ,
         \scp_reg[15][4] , \scp_reg[15][3] , \scp_reg[15][2] ,
         \scp_reg[15][1] , \scp_reg[15][0] , N30, N72, \pre_reg[12][0] ,
         \pre_reg[13][31] , \pre_reg[13][30] , \pre_reg[13][29] ,
         \pre_reg[13][28] , \pre_reg[13][27] , \pre_reg[13][26] ,
         \pre_reg[13][25] , \pre_reg[13][24] , \pre_reg[13][23] ,
         \pre_reg[13][22] , \pre_reg[13][21] , \pre_reg[13][20] ,
         \pre_reg[13][19] , \pre_reg[13][18] , \pre_reg[13][17] ,
         \pre_reg[13][16] , \pre_reg[13][15] , \pre_reg[13][14] ,
         \pre_reg[13][13] , \pre_reg[13][12] , \pre_reg[13][11] ,
         \pre_reg[13][10] , \pre_reg[13][9] , \pre_reg[13][8] ,
         \pre_reg[13][7] , \pre_reg[13][6] , \pre_reg[13][5] ,
         \pre_reg[13][4] , \pre_reg[13][3] , \pre_reg[13][2] ,
         \pre_reg[13][1] , \pre_reg[13][0] , \pre_reg[14][31] ,
         \pre_reg[14][30] , \pre_reg[14][29] , \pre_reg[14][28] ,
         \pre_reg[14][27] , \pre_reg[14][26] , \pre_reg[14][25] ,
         \pre_reg[14][24] , \pre_reg[14][23] , \pre_reg[14][22] ,
         \pre_reg[14][21] , \pre_reg[14][20] , \pre_reg[14][19] ,
         \pre_reg[14][18] , \pre_reg[14][17] , \pre_reg[14][16] ,
         \pre_reg[14][15] , \pre_reg[14][14] , \pre_reg[14][13] ,
         \pre_reg[14][12] , \pre_reg[14][11] , \pre_reg[14][10] ,
         \pre_reg[14][9] , \pre_reg[14][8] , \pre_reg[14][7] ,
         \pre_reg[14][6] , \pre_reg[14][5] , \pre_reg[14][4] ,
         \pre_reg[14][3] , \pre_reg[14][2] , \pre_reg[14][1] ,
         \pre_reg[14][0] , save_msk, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719;
  assign N30 = read_adr1[4];
  assign N72 = read_adr2[4];

  FLIP_FLOP_D \scp_reg_reg[12][31]  ( .D(n763), .CK(clock), .Q(
        \scp_reg[12][31] ) );
  FLIP_FLOP_D \scp_reg_reg[12][30]  ( .D(n764), .CK(clock), .Q(
        \scp_reg[12][30] ) );
  FLIP_FLOP_D \scp_reg_reg[12][29]  ( .D(n765), .CK(clock), .Q(
        \scp_reg[12][29] ) );
  FLIP_FLOP_D \scp_reg_reg[12][28]  ( .D(n766), .CK(clock), .Q(
        \scp_reg[12][28] ) );
  FLIP_FLOP_D \scp_reg_reg[12][27]  ( .D(n767), .CK(clock), .Q(
        \scp_reg[12][27] ) );
  FLIP_FLOP_D \scp_reg_reg[12][26]  ( .D(n768), .CK(clock), .Q(
        \scp_reg[12][26] ) );
  FLIP_FLOP_D \scp_reg_reg[12][25]  ( .D(n769), .CK(clock), .Q(
        \scp_reg[12][25] ) );
  FLIP_FLOP_D \scp_reg_reg[12][24]  ( .D(n770), .CK(clock), .Q(
        \scp_reg[12][24] ) );
  FLIP_FLOP_D \scp_reg_reg[12][23]  ( .D(n771), .CK(clock), .Q(
        \scp_reg[12][23] ) );
  FLIP_FLOP_D \scp_reg_reg[12][22]  ( .D(n772), .CK(clock), .Q(
        \scp_reg[12][22] ) );
  FLIP_FLOP_D \scp_reg_reg[12][21]  ( .D(n773), .CK(clock), .Q(
        \scp_reg[12][21] ) );
  FLIP_FLOP_D \scp_reg_reg[12][20]  ( .D(n774), .CK(clock), .Q(
        \scp_reg[12][20] ) );
  FLIP_FLOP_D \scp_reg_reg[12][19]  ( .D(n775), .CK(clock), .Q(
        \scp_reg[12][19] ) );
  FLIP_FLOP_D \scp_reg_reg[12][18]  ( .D(n776), .CK(clock), .Q(
        \scp_reg[12][18] ) );
  FLIP_FLOP_D \scp_reg_reg[12][17]  ( .D(n777), .CK(clock), .Q(
        \scp_reg[12][17] ) );
  FLIP_FLOP_D \scp_reg_reg[12][16]  ( .D(n778), .CK(clock), .Q(
        \scp_reg[12][16] ) );
  FLIP_FLOP_D \scp_reg_reg[12][15]  ( .D(n779), .CK(clock), .Q(
        \scp_reg[12][15] ) );
  FLIP_FLOP_D \scp_reg_reg[12][14]  ( .D(n780), .CK(clock), .Q(
        \scp_reg[12][14] ) );
  FLIP_FLOP_D \scp_reg_reg[12][13]  ( .D(n781), .CK(clock), .Q(
        \scp_reg[12][13] ) );
  FLIP_FLOP_D \scp_reg_reg[12][12]  ( .D(n782), .CK(clock), .Q(
        \scp_reg[12][12] ) );
  FLIP_FLOP_D \scp_reg_reg[12][11]  ( .D(n783), .CK(clock), .Q(
        \scp_reg[12][11] ) );
  FLIP_FLOP_D \scp_reg_reg[12][10]  ( .D(n784), .CK(clock), .Q(
        \scp_reg[12][10] ) );
  FLIP_FLOP_D \scp_reg_reg[12][9]  ( .D(n785), .CK(clock), .Q(\scp_reg[12][9] ) );
  FLIP_FLOP_D \scp_reg_reg[12][8]  ( .D(n786), .CK(clock), .Q(\scp_reg[12][8] ) );
  FLIP_FLOP_D \scp_reg_reg[12][7]  ( .D(n787), .CK(clock), .Q(\scp_reg[12][7] ) );
  FLIP_FLOP_D \scp_reg_reg[12][6]  ( .D(n788), .CK(clock), .Q(\scp_reg[12][6] ) );
  FLIP_FLOP_D \scp_reg_reg[12][5]  ( .D(n789), .CK(clock), .Q(\scp_reg[12][5] ) );
  FLIP_FLOP_D \scp_reg_reg[12][4]  ( .D(n790), .CK(clock), .Q(\scp_reg[12][4] ) );
  FLIP_FLOP_D \scp_reg_reg[12][3]  ( .D(n791), .CK(clock), .Q(\scp_reg[12][3] ) );
  FLIP_FLOP_D \scp_reg_reg[12][2]  ( .D(n792), .CK(clock), .Q(\scp_reg[12][2] ) );
  FLIP_FLOP_D \scp_reg_reg[12][1]  ( .D(n793), .CK(clock), .Q(\scp_reg[12][1] ) );
  FLIP_FLOP_D \scp_reg_reg[12][0]  ( .D(\pre_reg[12][0] ), .CK(clock), .Q(
        \scp_reg[12][0] ) );
  FLIP_FLOP_D save_msk_reg ( .D(n794), .CK(clock), .Q(save_msk) );
  FLIP_FLOP_D \scp_reg_reg[13][31]  ( .D(\pre_reg[13][31] ), .CK(clock), .Q(
        \scp_reg[13][31] ) );
  FLIP_FLOP_D \scp_reg_reg[13][30]  ( .D(\pre_reg[13][30] ), .CK(clock), .Q(
        \scp_reg[13][30] ) );
  FLIP_FLOP_D \scp_reg_reg[13][29]  ( .D(\pre_reg[13][29] ), .CK(clock), .Q(
        \scp_reg[13][29] ) );
  FLIP_FLOP_D \scp_reg_reg[13][28]  ( .D(\pre_reg[13][28] ), .CK(clock), .Q(
        \scp_reg[13][28] ) );
  FLIP_FLOP_D \scp_reg_reg[13][27]  ( .D(\pre_reg[13][27] ), .CK(clock), .Q(
        \scp_reg[13][27] ) );
  FLIP_FLOP_D \scp_reg_reg[13][26]  ( .D(\pre_reg[13][26] ), .CK(clock), .Q(
        \scp_reg[13][26] ) );
  FLIP_FLOP_D \scp_reg_reg[13][25]  ( .D(\pre_reg[13][25] ), .CK(clock), .Q(
        \scp_reg[13][25] ) );
  FLIP_FLOP_D \scp_reg_reg[13][24]  ( .D(\pre_reg[13][24] ), .CK(clock), .Q(
        \scp_reg[13][24] ) );
  FLIP_FLOP_D \scp_reg_reg[13][23]  ( .D(\pre_reg[13][23] ), .CK(clock), .Q(
        \scp_reg[13][23] ) );
  FLIP_FLOP_D \scp_reg_reg[13][22]  ( .D(\pre_reg[13][22] ), .CK(clock), .Q(
        \scp_reg[13][22] ) );
  FLIP_FLOP_D \scp_reg_reg[13][21]  ( .D(\pre_reg[13][21] ), .CK(clock), .Q(
        \scp_reg[13][21] ) );
  FLIP_FLOP_D \scp_reg_reg[13][20]  ( .D(\pre_reg[13][20] ), .CK(clock), .Q(
        \scp_reg[13][20] ) );
  FLIP_FLOP_D \scp_reg_reg[13][19]  ( .D(\pre_reg[13][19] ), .CK(clock), .Q(
        \scp_reg[13][19] ) );
  FLIP_FLOP_D \scp_reg_reg[13][18]  ( .D(\pre_reg[13][18] ), .CK(clock), .Q(
        \scp_reg[13][18] ) );
  FLIP_FLOP_D \scp_reg_reg[13][17]  ( .D(\pre_reg[13][17] ), .CK(clock), .Q(
        \scp_reg[13][17] ) );
  FLIP_FLOP_D \scp_reg_reg[13][16]  ( .D(\pre_reg[13][16] ), .CK(clock), .Q(
        \scp_reg[13][16] ) );
  FLIP_FLOP_D \scp_reg_reg[13][15]  ( .D(\pre_reg[13][15] ), .CK(clock), .Q(
        \scp_reg[13][15] ) );
  FLIP_FLOP_D \scp_reg_reg[13][14]  ( .D(\pre_reg[13][14] ), .CK(clock), .Q(
        \scp_reg[13][14] ) );
  FLIP_FLOP_D \scp_reg_reg[13][13]  ( .D(\pre_reg[13][13] ), .CK(clock), .Q(
        \scp_reg[13][13] ) );
  FLIP_FLOP_D \scp_reg_reg[13][12]  ( .D(\pre_reg[13][12] ), .CK(clock), .Q(
        \scp_reg[13][12] ) );
  FLIP_FLOP_D \scp_reg_reg[13][11]  ( .D(\pre_reg[13][11] ), .CK(clock), .Q(
        \scp_reg[13][11] ) );
  FLIP_FLOP_D \scp_reg_reg[13][10]  ( .D(\pre_reg[13][10] ), .CK(clock), .Q(
        \scp_reg[13][10] ) );
  FLIP_FLOP_D \scp_reg_reg[13][9]  ( .D(\pre_reg[13][9] ), .CK(clock), .Q(
        \scp_reg[13][9] ) );
  FLIP_FLOP_D \scp_reg_reg[13][8]  ( .D(\pre_reg[13][8] ), .CK(clock), .Q(
        \scp_reg[13][8] ) );
  FLIP_FLOP_D \scp_reg_reg[13][7]  ( .D(\pre_reg[13][7] ), .CK(clock), .Q(
        \scp_reg[13][7] ) );
  FLIP_FLOP_D \scp_reg_reg[13][6]  ( .D(\pre_reg[13][6] ), .CK(clock), .Q(
        \scp_reg[13][6] ) );
  FLIP_FLOP_D \scp_reg_reg[13][5]  ( .D(\pre_reg[13][5] ), .CK(clock), .Q(
        \scp_reg[13][5] ) );
  FLIP_FLOP_D \scp_reg_reg[13][4]  ( .D(\pre_reg[13][4] ), .CK(clock), .Q(
        \scp_reg[13][4] ) );
  FLIP_FLOP_D \scp_reg_reg[13][3]  ( .D(\pre_reg[13][3] ), .CK(clock), .Q(
        \scp_reg[13][3] ) );
  FLIP_FLOP_D \scp_reg_reg[13][2]  ( .D(\pre_reg[13][2] ), .CK(clock), .Q(
        \scp_reg[13][2] ) );
  FLIP_FLOP_D \scp_reg_reg[13][1]  ( .D(\pre_reg[13][1] ), .CK(clock), .Q(
        \scp_reg[13][1] ) );
  FLIP_FLOP_D \scp_reg_reg[13][0]  ( .D(\pre_reg[13][0] ), .CK(clock), .Q(
        \scp_reg[13][0] ) );
  FLIP_FLOP_D \scp_reg_reg[14][31]  ( .D(\pre_reg[14][31] ), .CK(clock), .Q(
        \scp_reg[14][31] ) );
  FLIP_FLOP_D \scp_reg_reg[14][30]  ( .D(\pre_reg[14][30] ), .CK(clock), .Q(
        \scp_reg[14][30] ) );
  FLIP_FLOP_D \scp_reg_reg[14][29]  ( .D(\pre_reg[14][29] ), .CK(clock), .Q(
        \scp_reg[14][29] ) );
  FLIP_FLOP_D \scp_reg_reg[14][28]  ( .D(\pre_reg[14][28] ), .CK(clock), .Q(
        \scp_reg[14][28] ) );
  FLIP_FLOP_D \scp_reg_reg[14][27]  ( .D(\pre_reg[14][27] ), .CK(clock), .Q(
        \scp_reg[14][27] ) );
  FLIP_FLOP_D \scp_reg_reg[14][26]  ( .D(\pre_reg[14][26] ), .CK(clock), .Q(
        \scp_reg[14][26] ) );
  FLIP_FLOP_D \scp_reg_reg[14][25]  ( .D(\pre_reg[14][25] ), .CK(clock), .Q(
        \scp_reg[14][25] ) );
  FLIP_FLOP_D \scp_reg_reg[14][24]  ( .D(\pre_reg[14][24] ), .CK(clock), .Q(
        \scp_reg[14][24] ) );
  FLIP_FLOP_D \scp_reg_reg[14][23]  ( .D(\pre_reg[14][23] ), .CK(clock), .Q(
        \scp_reg[14][23] ) );
  FLIP_FLOP_D \scp_reg_reg[14][22]  ( .D(\pre_reg[14][22] ), .CK(clock), .Q(
        \scp_reg[14][22] ) );
  FLIP_FLOP_D \scp_reg_reg[14][21]  ( .D(\pre_reg[14][21] ), .CK(clock), .Q(
        \scp_reg[14][21] ) );
  FLIP_FLOP_D \scp_reg_reg[14][20]  ( .D(\pre_reg[14][20] ), .CK(clock), .Q(
        \scp_reg[14][20] ) );
  FLIP_FLOP_D \scp_reg_reg[14][19]  ( .D(\pre_reg[14][19] ), .CK(clock), .Q(
        \scp_reg[14][19] ) );
  FLIP_FLOP_D \scp_reg_reg[14][18]  ( .D(\pre_reg[14][18] ), .CK(clock), .Q(
        \scp_reg[14][18] ) );
  FLIP_FLOP_D \scp_reg_reg[14][17]  ( .D(\pre_reg[14][17] ), .CK(clock), .Q(
        \scp_reg[14][17] ) );
  FLIP_FLOP_D \scp_reg_reg[14][16]  ( .D(\pre_reg[14][16] ), .CK(clock), .Q(
        \scp_reg[14][16] ) );
  FLIP_FLOP_D \scp_reg_reg[14][15]  ( .D(\pre_reg[14][15] ), .CK(clock), .Q(
        \scp_reg[14][15] ) );
  FLIP_FLOP_D \scp_reg_reg[14][14]  ( .D(\pre_reg[14][14] ), .CK(clock), .Q(
        \scp_reg[14][14] ) );
  FLIP_FLOP_D \scp_reg_reg[14][13]  ( .D(\pre_reg[14][13] ), .CK(clock), .Q(
        \scp_reg[14][13] ) );
  FLIP_FLOP_D \scp_reg_reg[14][12]  ( .D(\pre_reg[14][12] ), .CK(clock), .Q(
        \scp_reg[14][12] ) );
  FLIP_FLOP_D \scp_reg_reg[14][11]  ( .D(\pre_reg[14][11] ), .CK(clock), .Q(
        \scp_reg[14][11] ) );
  FLIP_FLOP_D \scp_reg_reg[14][10]  ( .D(\pre_reg[14][10] ), .CK(clock), .Q(
        \scp_reg[14][10] ) );
  FLIP_FLOP_D \scp_reg_reg[14][9]  ( .D(\pre_reg[14][9] ), .CK(clock), .Q(
        \scp_reg[14][9] ) );
  FLIP_FLOP_D \scp_reg_reg[14][8]  ( .D(\pre_reg[14][8] ), .CK(clock), .Q(
        \scp_reg[14][8] ) );
  FLIP_FLOP_D \scp_reg_reg[14][7]  ( .D(\pre_reg[14][7] ), .CK(clock), .Q(
        \scp_reg[14][7] ) );
  FLIP_FLOP_D \scp_reg_reg[14][6]  ( .D(\pre_reg[14][6] ), .CK(clock), .Q(
        \scp_reg[14][6] ) );
  FLIP_FLOP_D \scp_reg_reg[14][5]  ( .D(\pre_reg[14][5] ), .CK(clock), .Q(
        \scp_reg[14][5] ) );
  FLIP_FLOP_D \scp_reg_reg[14][4]  ( .D(\pre_reg[14][4] ), .CK(clock), .Q(
        \scp_reg[14][4] ) );
  FLIP_FLOP_D \scp_reg_reg[14][3]  ( .D(\pre_reg[14][3] ), .CK(clock), .Q(
        \scp_reg[14][3] ) );
  FLIP_FLOP_D \scp_reg_reg[14][2]  ( .D(\pre_reg[14][2] ), .CK(clock), .Q(
        \scp_reg[14][2] ) );
  FLIP_FLOP_D \scp_reg_reg[14][1]  ( .D(\pre_reg[14][1] ), .CK(clock), .Q(
        \scp_reg[14][1] ) );
  FLIP_FLOP_D \scp_reg_reg[14][0]  ( .D(\pre_reg[14][0] ), .CK(clock), .Q(
        \scp_reg[14][0] ) );
  FLIP_FLOP_D \scp_reg_reg[15][31]  ( .D(n762), .CK(clock), .Q(
        \scp_reg[15][31] ) );
  FLIP_FLOP_D \scp_reg_reg[15][30]  ( .D(n761), .CK(clock), .Q(
        \scp_reg[15][30] ) );
  FLIP_FLOP_D \scp_reg_reg[15][29]  ( .D(n760), .CK(clock), .Q(
        \scp_reg[15][29] ) );
  FLIP_FLOP_D \scp_reg_reg[15][28]  ( .D(n759), .CK(clock), .Q(
        \scp_reg[15][28] ) );
  FLIP_FLOP_D \scp_reg_reg[15][27]  ( .D(n758), .CK(clock), .Q(
        \scp_reg[15][27] ) );
  FLIP_FLOP_D \scp_reg_reg[15][26]  ( .D(n757), .CK(clock), .Q(
        \scp_reg[15][26] ) );
  FLIP_FLOP_D \scp_reg_reg[15][25]  ( .D(n756), .CK(clock), .Q(
        \scp_reg[15][25] ) );
  FLIP_FLOP_D \scp_reg_reg[15][24]  ( .D(n755), .CK(clock), .Q(
        \scp_reg[15][24] ) );
  FLIP_FLOP_D \scp_reg_reg[15][23]  ( .D(n754), .CK(clock), .Q(
        \scp_reg[15][23] ) );
  FLIP_FLOP_D \scp_reg_reg[15][22]  ( .D(n753), .CK(clock), .Q(
        \scp_reg[15][22] ) );
  FLIP_FLOP_D \scp_reg_reg[15][21]  ( .D(n752), .CK(clock), .Q(
        \scp_reg[15][21] ) );
  FLIP_FLOP_D \scp_reg_reg[15][20]  ( .D(n751), .CK(clock), .Q(
        \scp_reg[15][20] ) );
  FLIP_FLOP_D \scp_reg_reg[15][19]  ( .D(n750), .CK(clock), .Q(
        \scp_reg[15][19] ) );
  FLIP_FLOP_D \scp_reg_reg[15][18]  ( .D(n749), .CK(clock), .Q(
        \scp_reg[15][18] ) );
  FLIP_FLOP_D \scp_reg_reg[15][17]  ( .D(n748), .CK(clock), .Q(
        \scp_reg[15][17] ) );
  FLIP_FLOP_D \scp_reg_reg[15][16]  ( .D(n747), .CK(clock), .Q(
        \scp_reg[15][16] ) );
  FLIP_FLOP_D \scp_reg_reg[15][15]  ( .D(n746), .CK(clock), .Q(
        \scp_reg[15][15] ) );
  FLIP_FLOP_D \scp_reg_reg[15][14]  ( .D(n745), .CK(clock), .Q(
        \scp_reg[15][14] ) );
  FLIP_FLOP_D \scp_reg_reg[15][13]  ( .D(n744), .CK(clock), .Q(
        \scp_reg[15][13] ) );
  FLIP_FLOP_D \scp_reg_reg[15][12]  ( .D(n743), .CK(clock), .Q(
        \scp_reg[15][12] ) );
  FLIP_FLOP_D \scp_reg_reg[15][11]  ( .D(n742), .CK(clock), .Q(
        \scp_reg[15][11] ) );
  FLIP_FLOP_D \scp_reg_reg[15][10]  ( .D(n741), .CK(clock), .Q(
        \scp_reg[15][10] ) );
  FLIP_FLOP_D \scp_reg_reg[15][9]  ( .D(n740), .CK(clock), .Q(\scp_reg[15][9] ) );
  FLIP_FLOP_D \scp_reg_reg[15][8]  ( .D(n739), .CK(clock), .Q(\scp_reg[15][8] ) );
  FLIP_FLOP_D \scp_reg_reg[15][7]  ( .D(n738), .CK(clock), .Q(\scp_reg[15][7] ) );
  FLIP_FLOP_D \scp_reg_reg[15][6]  ( .D(n737), .CK(clock), .Q(\scp_reg[15][6] ) );
  FLIP_FLOP_D \scp_reg_reg[15][5]  ( .D(n736), .CK(clock), .Q(\scp_reg[15][5] ) );
  FLIP_FLOP_D \scp_reg_reg[15][4]  ( .D(n735), .CK(clock), .Q(\scp_reg[15][4] ) );
  FLIP_FLOP_D \scp_reg_reg[15][3]  ( .D(n734), .CK(clock), .Q(\scp_reg[15][3] ) );
  FLIP_FLOP_D \scp_reg_reg[15][2]  ( .D(n733), .CK(clock), .Q(\scp_reg[15][2] ) );
  FLIP_FLOP_D \scp_reg_reg[15][1]  ( .D(n732), .CK(clock), .Q(\scp_reg[15][1] ) );
  FLIP_FLOP_D \scp_reg_reg[15][0]  ( .D(n731), .CK(clock), .Q(\scp_reg[15][0] ) );
  INV_GATE U3 ( .I1(n7), .O(n1) );
  INV_GATE U4 ( .I1(write_data[0]), .O(n2) );
  INV_GATE U5 ( .I1(write_data[2]), .O(n3) );
  INV_GATE U6 ( .I1(reset), .O(n4) );
  NAND_GATE U7 ( .I1(n5), .I2(n6), .O(vecteur_it[9]) );
  NAND_GATE U8 ( .I1(\scp_reg[14][9] ), .I2(n7), .O(n6) );
  NAND_GATE U9 ( .I1(\scp_reg[15][9] ), .I2(n1), .O(n5) );
  NAND_GATE U10 ( .I1(n8), .I2(n9), .O(vecteur_it[8]) );
  NAND_GATE U11 ( .I1(\scp_reg[14][8] ), .I2(n7), .O(n9) );
  NAND_GATE U12 ( .I1(\scp_reg[15][8] ), .I2(n1), .O(n8) );
  NAND_GATE U13 ( .I1(n10), .I2(n11), .O(vecteur_it[7]) );
  NAND_GATE U14 ( .I1(\scp_reg[14][7] ), .I2(n7), .O(n11) );
  NAND_GATE U15 ( .I1(\scp_reg[15][7] ), .I2(n1), .O(n10) );
  NAND_GATE U16 ( .I1(n12), .I2(n13), .O(vecteur_it[6]) );
  NAND_GATE U17 ( .I1(\scp_reg[14][6] ), .I2(n7), .O(n13) );
  NAND_GATE U18 ( .I1(\scp_reg[15][6] ), .I2(n1), .O(n12) );
  NAND_GATE U19 ( .I1(n14), .I2(n15), .O(vecteur_it[5]) );
  NAND_GATE U20 ( .I1(\scp_reg[14][5] ), .I2(n7), .O(n15) );
  NAND_GATE U21 ( .I1(\scp_reg[15][5] ), .I2(n1), .O(n14) );
  NAND_GATE U22 ( .I1(n16), .I2(n17), .O(vecteur_it[4]) );
  NAND_GATE U23 ( .I1(\scp_reg[14][4] ), .I2(n7), .O(n17) );
  NAND_GATE U24 ( .I1(\scp_reg[15][4] ), .I2(n1), .O(n16) );
  NAND_GATE U25 ( .I1(n18), .I2(n19), .O(vecteur_it[3]) );
  NAND_GATE U26 ( .I1(\scp_reg[14][3] ), .I2(n7), .O(n19) );
  NAND_GATE U27 ( .I1(\scp_reg[15][3] ), .I2(n1), .O(n18) );
  NAND_GATE U28 ( .I1(n20), .I2(n21), .O(vecteur_it[31]) );
  NAND_GATE U29 ( .I1(\scp_reg[14][31] ), .I2(n7), .O(n21) );
  NAND_GATE U30 ( .I1(\scp_reg[15][31] ), .I2(n1), .O(n20) );
  NAND_GATE U31 ( .I1(n22), .I2(n23), .O(vecteur_it[30]) );
  NAND_GATE U32 ( .I1(\scp_reg[14][30] ), .I2(n7), .O(n23) );
  NAND_GATE U33 ( .I1(\scp_reg[15][30] ), .I2(n1), .O(n22) );
  NAND_GATE U34 ( .I1(n24), .I2(n25), .O(vecteur_it[2]) );
  NAND_GATE U35 ( .I1(\scp_reg[14][2] ), .I2(n7), .O(n25) );
  NAND_GATE U36 ( .I1(\scp_reg[15][2] ), .I2(n1), .O(n24) );
  NAND_GATE U37 ( .I1(n26), .I2(n27), .O(vecteur_it[29]) );
  NAND_GATE U38 ( .I1(\scp_reg[14][29] ), .I2(n7), .O(n27) );
  NAND_GATE U39 ( .I1(\scp_reg[15][29] ), .I2(n1), .O(n26) );
  NAND_GATE U40 ( .I1(n28), .I2(n29), .O(vecteur_it[28]) );
  NAND_GATE U41 ( .I1(\scp_reg[14][28] ), .I2(n7), .O(n29) );
  NAND_GATE U42 ( .I1(\scp_reg[15][28] ), .I2(n1), .O(n28) );
  NAND_GATE U43 ( .I1(n30), .I2(n31), .O(vecteur_it[27]) );
  NAND_GATE U44 ( .I1(\scp_reg[14][27] ), .I2(n7), .O(n31) );
  NAND_GATE U45 ( .I1(\scp_reg[15][27] ), .I2(n1), .O(n30) );
  NAND_GATE U46 ( .I1(n32), .I2(n33), .O(vecteur_it[26]) );
  NAND_GATE U47 ( .I1(\scp_reg[14][26] ), .I2(n7), .O(n33) );
  NAND_GATE U48 ( .I1(\scp_reg[15][26] ), .I2(n1), .O(n32) );
  NAND_GATE U49 ( .I1(n34), .I2(n35), .O(vecteur_it[25]) );
  NAND_GATE U50 ( .I1(\scp_reg[14][25] ), .I2(n7), .O(n35) );
  NAND_GATE U51 ( .I1(\scp_reg[15][25] ), .I2(n1), .O(n34) );
  NAND_GATE U52 ( .I1(n36), .I2(n37), .O(vecteur_it[24]) );
  NAND_GATE U53 ( .I1(\scp_reg[14][24] ), .I2(n7), .O(n37) );
  NAND_GATE U54 ( .I1(\scp_reg[15][24] ), .I2(n1), .O(n36) );
  NAND_GATE U55 ( .I1(n38), .I2(n39), .O(vecteur_it[23]) );
  NAND_GATE U56 ( .I1(\scp_reg[14][23] ), .I2(n7), .O(n39) );
  NAND_GATE U57 ( .I1(\scp_reg[15][23] ), .I2(n1), .O(n38) );
  NAND_GATE U58 ( .I1(n40), .I2(n41), .O(vecteur_it[22]) );
  NAND_GATE U59 ( .I1(\scp_reg[14][22] ), .I2(n7), .O(n41) );
  NAND_GATE U60 ( .I1(\scp_reg[15][22] ), .I2(n1), .O(n40) );
  NAND_GATE U61 ( .I1(n42), .I2(n43), .O(vecteur_it[21]) );
  NAND_GATE U62 ( .I1(\scp_reg[14][21] ), .I2(n7), .O(n43) );
  NAND_GATE U63 ( .I1(\scp_reg[15][21] ), .I2(n1), .O(n42) );
  NAND_GATE U64 ( .I1(n44), .I2(n45), .O(vecteur_it[20]) );
  NAND_GATE U65 ( .I1(\scp_reg[14][20] ), .I2(n7), .O(n45) );
  NAND_GATE U66 ( .I1(\scp_reg[15][20] ), .I2(n1), .O(n44) );
  NAND_GATE U67 ( .I1(n46), .I2(n47), .O(vecteur_it[1]) );
  NAND_GATE U68 ( .I1(\scp_reg[14][1] ), .I2(n7), .O(n47) );
  NAND_GATE U69 ( .I1(\scp_reg[15][1] ), .I2(n1), .O(n46) );
  NAND_GATE U70 ( .I1(n48), .I2(n49), .O(vecteur_it[19]) );
  NAND_GATE U71 ( .I1(\scp_reg[14][19] ), .I2(n7), .O(n49) );
  NAND_GATE U72 ( .I1(\scp_reg[15][19] ), .I2(n1), .O(n48) );
  NAND_GATE U73 ( .I1(n50), .I2(n51), .O(vecteur_it[18]) );
  NAND_GATE U74 ( .I1(\scp_reg[14][18] ), .I2(n7), .O(n51) );
  NAND_GATE U75 ( .I1(\scp_reg[15][18] ), .I2(n1), .O(n50) );
  NAND_GATE U76 ( .I1(n52), .I2(n53), .O(vecteur_it[17]) );
  NAND_GATE U77 ( .I1(\scp_reg[14][17] ), .I2(n7), .O(n53) );
  NAND_GATE U78 ( .I1(\scp_reg[15][17] ), .I2(n1), .O(n52) );
  NAND_GATE U79 ( .I1(n54), .I2(n55), .O(vecteur_it[16]) );
  NAND_GATE U80 ( .I1(\scp_reg[14][16] ), .I2(n7), .O(n55) );
  NAND_GATE U81 ( .I1(\scp_reg[15][16] ), .I2(n1), .O(n54) );
  NAND_GATE U82 ( .I1(n56), .I2(n57), .O(vecteur_it[15]) );
  NAND_GATE U83 ( .I1(\scp_reg[14][15] ), .I2(n7), .O(n57) );
  NAND_GATE U84 ( .I1(\scp_reg[15][15] ), .I2(n1), .O(n56) );
  NAND_GATE U85 ( .I1(n58), .I2(n59), .O(vecteur_it[14]) );
  NAND_GATE U86 ( .I1(\scp_reg[14][14] ), .I2(n7), .O(n59) );
  NAND_GATE U87 ( .I1(\scp_reg[15][14] ), .I2(n1), .O(n58) );
  NAND_GATE U88 ( .I1(n60), .I2(n61), .O(vecteur_it[13]) );
  NAND_GATE U89 ( .I1(\scp_reg[14][13] ), .I2(n7), .O(n61) );
  NAND_GATE U90 ( .I1(\scp_reg[15][13] ), .I2(n1), .O(n60) );
  NAND_GATE U91 ( .I1(n62), .I2(n63), .O(vecteur_it[12]) );
  NAND_GATE U92 ( .I1(\scp_reg[14][12] ), .I2(n7), .O(n63) );
  NAND_GATE U93 ( .I1(\scp_reg[15][12] ), .I2(n1), .O(n62) );
  NAND_GATE U94 ( .I1(n64), .I2(n65), .O(vecteur_it[11]) );
  NAND_GATE U95 ( .I1(\scp_reg[14][11] ), .I2(n7), .O(n65) );
  NAND_GATE U96 ( .I1(\scp_reg[15][11] ), .I2(n1), .O(n64) );
  NAND_GATE U97 ( .I1(n66), .I2(n67), .O(vecteur_it[10]) );
  NAND_GATE U98 ( .I1(\scp_reg[14][10] ), .I2(n7), .O(n67) );
  NAND_GATE U99 ( .I1(\scp_reg[15][10] ), .I2(n1), .O(n66) );
  NAND_GATE U100 ( .I1(n68), .I2(n69), .O(vecteur_it[0]) );
  NAND_GATE U101 ( .I1(\scp_reg[14][0] ), .I2(n7), .O(n69) );
  NAND_GATE U102 ( .I1(\scp_reg[15][0] ), .I2(n1), .O(n68) );
  NAND4_GATE U103 ( .I1(n70), .I2(n71), .I3(n72), .I4(n73), .O(read_data2[9])
         );
  NAND_GATE U104 ( .I1(n74), .I2(\scp_reg[15][9] ), .O(n73) );
  NAND_GATE U105 ( .I1(n75), .I2(\scp_reg[14][9] ), .O(n72) );
  NAND_GATE U106 ( .I1(\scp_reg[13][9] ), .I2(n76), .O(n71) );
  NAND_GATE U107 ( .I1(\scp_reg[12][9] ), .I2(n77), .O(n70) );
  NAND4_GATE U108 ( .I1(n78), .I2(n79), .I3(n80), .I4(n81), .O(read_data2[8])
         );
  NAND_GATE U109 ( .I1(n74), .I2(\scp_reg[15][8] ), .O(n81) );
  NAND_GATE U110 ( .I1(n75), .I2(\scp_reg[14][8] ), .O(n80) );
  NAND_GATE U111 ( .I1(\scp_reg[13][8] ), .I2(n76), .O(n79) );
  NAND_GATE U112 ( .I1(\scp_reg[12][8] ), .I2(n77), .O(n78) );
  NAND4_GATE U113 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .O(read_data2[7])
         );
  NAND_GATE U114 ( .I1(n74), .I2(\scp_reg[15][7] ), .O(n85) );
  NAND_GATE U115 ( .I1(n75), .I2(\scp_reg[14][7] ), .O(n84) );
  NAND_GATE U116 ( .I1(\scp_reg[13][7] ), .I2(n76), .O(n83) );
  NAND_GATE U117 ( .I1(\scp_reg[12][7] ), .I2(n77), .O(n82) );
  NAND4_GATE U118 ( .I1(n86), .I2(n87), .I3(n88), .I4(n89), .O(read_data2[6])
         );
  NAND_GATE U119 ( .I1(n74), .I2(\scp_reg[15][6] ), .O(n89) );
  NAND_GATE U120 ( .I1(n75), .I2(\scp_reg[14][6] ), .O(n88) );
  NAND_GATE U121 ( .I1(\scp_reg[13][6] ), .I2(n76), .O(n87) );
  NAND_GATE U122 ( .I1(\scp_reg[12][6] ), .I2(n77), .O(n86) );
  NAND4_GATE U123 ( .I1(n90), .I2(n91), .I3(n92), .I4(n93), .O(read_data2[5])
         );
  NAND_GATE U124 ( .I1(n74), .I2(\scp_reg[15][5] ), .O(n93) );
  NAND_GATE U125 ( .I1(n75), .I2(\scp_reg[14][5] ), .O(n92) );
  NAND_GATE U126 ( .I1(\scp_reg[13][5] ), .I2(n76), .O(n91) );
  NAND_GATE U127 ( .I1(\scp_reg[12][5] ), .I2(n77), .O(n90) );
  NAND4_GATE U128 ( .I1(n94), .I2(n95), .I3(n96), .I4(n97), .O(read_data2[4])
         );
  NAND_GATE U129 ( .I1(n74), .I2(\scp_reg[15][4] ), .O(n97) );
  NAND_GATE U130 ( .I1(n75), .I2(\scp_reg[14][4] ), .O(n96) );
  NAND_GATE U131 ( .I1(\scp_reg[13][4] ), .I2(n76), .O(n95) );
  NAND_GATE U132 ( .I1(\scp_reg[12][4] ), .I2(n77), .O(n94) );
  NAND4_GATE U133 ( .I1(n98), .I2(n99), .I3(n100), .I4(n101), .O(read_data2[3]) );
  NAND_GATE U134 ( .I1(n74), .I2(\scp_reg[15][3] ), .O(n101) );
  NAND_GATE U135 ( .I1(n75), .I2(\scp_reg[14][3] ), .O(n100) );
  NAND_GATE U136 ( .I1(\scp_reg[13][3] ), .I2(n76), .O(n99) );
  NAND_GATE U137 ( .I1(\scp_reg[12][3] ), .I2(n77), .O(n98) );
  NAND4_GATE U138 ( .I1(n102), .I2(n103), .I3(n104), .I4(n105), .O(
        read_data2[31]) );
  NAND_GATE U139 ( .I1(n74), .I2(\scp_reg[15][31] ), .O(n105) );
  NAND_GATE U140 ( .I1(n75), .I2(\scp_reg[14][31] ), .O(n104) );
  NAND_GATE U141 ( .I1(\scp_reg[13][31] ), .I2(n76), .O(n103) );
  NAND_GATE U142 ( .I1(\scp_reg[12][31] ), .I2(n77), .O(n102) );
  NAND4_GATE U143 ( .I1(n106), .I2(n107), .I3(n108), .I4(n109), .O(
        read_data2[30]) );
  NAND_GATE U144 ( .I1(n74), .I2(\scp_reg[15][30] ), .O(n109) );
  NAND_GATE U145 ( .I1(n75), .I2(\scp_reg[14][30] ), .O(n108) );
  NAND_GATE U146 ( .I1(\scp_reg[13][30] ), .I2(n76), .O(n107) );
  NAND_GATE U147 ( .I1(\scp_reg[12][30] ), .I2(n77), .O(n106) );
  NAND4_GATE U148 ( .I1(n110), .I2(n111), .I3(n112), .I4(n113), .O(
        read_data2[2]) );
  NAND_GATE U149 ( .I1(n74), .I2(\scp_reg[15][2] ), .O(n113) );
  NAND_GATE U150 ( .I1(n75), .I2(\scp_reg[14][2] ), .O(n112) );
  NAND_GATE U151 ( .I1(\scp_reg[13][2] ), .I2(n76), .O(n111) );
  NAND_GATE U152 ( .I1(\scp_reg[12][2] ), .I2(n77), .O(n110) );
  NAND4_GATE U153 ( .I1(n114), .I2(n115), .I3(n116), .I4(n117), .O(
        read_data2[29]) );
  NAND_GATE U154 ( .I1(n74), .I2(\scp_reg[15][29] ), .O(n117) );
  NAND_GATE U155 ( .I1(n75), .I2(\scp_reg[14][29] ), .O(n116) );
  NAND_GATE U156 ( .I1(\scp_reg[13][29] ), .I2(n76), .O(n115) );
  NAND_GATE U157 ( .I1(\scp_reg[12][29] ), .I2(n77), .O(n114) );
  NAND4_GATE U158 ( .I1(n118), .I2(n119), .I3(n120), .I4(n121), .O(
        read_data2[28]) );
  NAND_GATE U159 ( .I1(n74), .I2(\scp_reg[15][28] ), .O(n121) );
  NAND_GATE U160 ( .I1(n75), .I2(\scp_reg[14][28] ), .O(n120) );
  NAND_GATE U161 ( .I1(\scp_reg[13][28] ), .I2(n76), .O(n119) );
  NAND_GATE U162 ( .I1(\scp_reg[12][28] ), .I2(n77), .O(n118) );
  NAND4_GATE U163 ( .I1(n122), .I2(n123), .I3(n124), .I4(n125), .O(
        read_data2[27]) );
  NAND_GATE U164 ( .I1(n74), .I2(\scp_reg[15][27] ), .O(n125) );
  NAND_GATE U165 ( .I1(n75), .I2(\scp_reg[14][27] ), .O(n124) );
  NAND_GATE U166 ( .I1(\scp_reg[13][27] ), .I2(n76), .O(n123) );
  NAND_GATE U167 ( .I1(\scp_reg[12][27] ), .I2(n77), .O(n122) );
  NAND4_GATE U168 ( .I1(n126), .I2(n127), .I3(n128), .I4(n129), .O(
        read_data2[26]) );
  NAND_GATE U169 ( .I1(n74), .I2(\scp_reg[15][26] ), .O(n129) );
  NAND_GATE U170 ( .I1(n75), .I2(\scp_reg[14][26] ), .O(n128) );
  NAND_GATE U171 ( .I1(\scp_reg[13][26] ), .I2(n76), .O(n127) );
  NAND_GATE U172 ( .I1(\scp_reg[12][26] ), .I2(n77), .O(n126) );
  NAND4_GATE U173 ( .I1(n130), .I2(n131), .I3(n132), .I4(n133), .O(
        read_data2[25]) );
  NAND_GATE U174 ( .I1(n74), .I2(\scp_reg[15][25] ), .O(n133) );
  NAND_GATE U175 ( .I1(n75), .I2(\scp_reg[14][25] ), .O(n132) );
  NAND_GATE U176 ( .I1(\scp_reg[13][25] ), .I2(n76), .O(n131) );
  NAND_GATE U177 ( .I1(\scp_reg[12][25] ), .I2(n77), .O(n130) );
  NAND4_GATE U178 ( .I1(n134), .I2(n135), .I3(n136), .I4(n137), .O(
        read_data2[24]) );
  NAND_GATE U179 ( .I1(n74), .I2(\scp_reg[15][24] ), .O(n137) );
  NAND_GATE U180 ( .I1(n75), .I2(\scp_reg[14][24] ), .O(n136) );
  NAND_GATE U181 ( .I1(\scp_reg[13][24] ), .I2(n76), .O(n135) );
  NAND_GATE U182 ( .I1(\scp_reg[12][24] ), .I2(n77), .O(n134) );
  NAND4_GATE U183 ( .I1(n138), .I2(n139), .I3(n140), .I4(n141), .O(
        read_data2[23]) );
  NAND_GATE U184 ( .I1(n74), .I2(\scp_reg[15][23] ), .O(n141) );
  NAND_GATE U185 ( .I1(n75), .I2(\scp_reg[14][23] ), .O(n140) );
  NAND_GATE U186 ( .I1(\scp_reg[13][23] ), .I2(n76), .O(n139) );
  NAND_GATE U187 ( .I1(\scp_reg[12][23] ), .I2(n77), .O(n138) );
  NAND4_GATE U188 ( .I1(n142), .I2(n143), .I3(n144), .I4(n145), .O(
        read_data2[22]) );
  NAND_GATE U189 ( .I1(n74), .I2(\scp_reg[15][22] ), .O(n145) );
  NAND_GATE U190 ( .I1(n75), .I2(\scp_reg[14][22] ), .O(n144) );
  NAND_GATE U191 ( .I1(\scp_reg[13][22] ), .I2(n76), .O(n143) );
  NAND_GATE U192 ( .I1(\scp_reg[12][22] ), .I2(n77), .O(n142) );
  NAND4_GATE U193 ( .I1(n146), .I2(n147), .I3(n148), .I4(n149), .O(
        read_data2[21]) );
  NAND_GATE U194 ( .I1(n74), .I2(\scp_reg[15][21] ), .O(n149) );
  NAND_GATE U195 ( .I1(n75), .I2(\scp_reg[14][21] ), .O(n148) );
  NAND_GATE U196 ( .I1(\scp_reg[13][21] ), .I2(n76), .O(n147) );
  NAND_GATE U197 ( .I1(\scp_reg[12][21] ), .I2(n77), .O(n146) );
  NAND4_GATE U198 ( .I1(n150), .I2(n151), .I3(n152), .I4(n153), .O(
        read_data2[20]) );
  NAND_GATE U199 ( .I1(n74), .I2(\scp_reg[15][20] ), .O(n153) );
  NAND_GATE U200 ( .I1(n75), .I2(\scp_reg[14][20] ), .O(n152) );
  NAND_GATE U201 ( .I1(\scp_reg[13][20] ), .I2(n76), .O(n151) );
  NAND_GATE U202 ( .I1(\scp_reg[12][20] ), .I2(n77), .O(n150) );
  NAND4_GATE U203 ( .I1(n154), .I2(n155), .I3(n156), .I4(n157), .O(
        read_data2[1]) );
  NAND_GATE U204 ( .I1(n74), .I2(\scp_reg[15][1] ), .O(n157) );
  NAND_GATE U205 ( .I1(n75), .I2(\scp_reg[14][1] ), .O(n156) );
  NAND_GATE U206 ( .I1(\scp_reg[13][1] ), .I2(n76), .O(n155) );
  NAND_GATE U207 ( .I1(\scp_reg[12][1] ), .I2(n77), .O(n154) );
  NAND4_GATE U208 ( .I1(n158), .I2(n159), .I3(n160), .I4(n161), .O(
        read_data2[19]) );
  NAND_GATE U209 ( .I1(n74), .I2(\scp_reg[15][19] ), .O(n161) );
  NAND_GATE U210 ( .I1(n75), .I2(\scp_reg[14][19] ), .O(n160) );
  NAND_GATE U211 ( .I1(\scp_reg[13][19] ), .I2(n76), .O(n159) );
  NAND_GATE U212 ( .I1(\scp_reg[12][19] ), .I2(n77), .O(n158) );
  NAND4_GATE U213 ( .I1(n162), .I2(n163), .I3(n164), .I4(n165), .O(
        read_data2[18]) );
  NAND_GATE U214 ( .I1(n74), .I2(\scp_reg[15][18] ), .O(n165) );
  NAND_GATE U215 ( .I1(n75), .I2(\scp_reg[14][18] ), .O(n164) );
  NAND_GATE U216 ( .I1(\scp_reg[13][18] ), .I2(n76), .O(n163) );
  NAND_GATE U217 ( .I1(\scp_reg[12][18] ), .I2(n77), .O(n162) );
  NAND4_GATE U218 ( .I1(n166), .I2(n167), .I3(n168), .I4(n169), .O(
        read_data2[17]) );
  NAND_GATE U219 ( .I1(n74), .I2(\scp_reg[15][17] ), .O(n169) );
  NAND_GATE U220 ( .I1(n75), .I2(\scp_reg[14][17] ), .O(n168) );
  NAND_GATE U221 ( .I1(\scp_reg[13][17] ), .I2(n76), .O(n167) );
  NAND_GATE U222 ( .I1(\scp_reg[12][17] ), .I2(n77), .O(n166) );
  NAND4_GATE U223 ( .I1(n170), .I2(n171), .I3(n172), .I4(n173), .O(
        read_data2[16]) );
  NAND_GATE U224 ( .I1(n74), .I2(\scp_reg[15][16] ), .O(n173) );
  NAND_GATE U225 ( .I1(n75), .I2(\scp_reg[14][16] ), .O(n172) );
  NAND_GATE U226 ( .I1(\scp_reg[13][16] ), .I2(n76), .O(n171) );
  NAND_GATE U227 ( .I1(\scp_reg[12][16] ), .I2(n77), .O(n170) );
  NAND4_GATE U228 ( .I1(n174), .I2(n175), .I3(n176), .I4(n177), .O(
        read_data2[15]) );
  NAND_GATE U229 ( .I1(n74), .I2(\scp_reg[15][15] ), .O(n177) );
  NAND_GATE U230 ( .I1(n75), .I2(\scp_reg[14][15] ), .O(n176) );
  NAND_GATE U231 ( .I1(\scp_reg[13][15] ), .I2(n76), .O(n175) );
  NAND_GATE U232 ( .I1(\scp_reg[12][15] ), .I2(n77), .O(n174) );
  NAND4_GATE U233 ( .I1(n178), .I2(n179), .I3(n180), .I4(n181), .O(
        read_data2[14]) );
  NAND_GATE U234 ( .I1(n74), .I2(\scp_reg[15][14] ), .O(n181) );
  NAND_GATE U235 ( .I1(n75), .I2(\scp_reg[14][14] ), .O(n180) );
  NAND_GATE U236 ( .I1(\scp_reg[13][14] ), .I2(n76), .O(n179) );
  NAND_GATE U237 ( .I1(\scp_reg[12][14] ), .I2(n77), .O(n178) );
  NAND4_GATE U238 ( .I1(n182), .I2(n183), .I3(n184), .I4(n185), .O(
        read_data2[13]) );
  NAND_GATE U239 ( .I1(n74), .I2(\scp_reg[15][13] ), .O(n185) );
  NAND_GATE U240 ( .I1(n75), .I2(\scp_reg[14][13] ), .O(n184) );
  NAND_GATE U241 ( .I1(\scp_reg[13][13] ), .I2(n76), .O(n183) );
  NAND_GATE U242 ( .I1(\scp_reg[12][13] ), .I2(n77), .O(n182) );
  NAND4_GATE U243 ( .I1(n186), .I2(n187), .I3(n188), .I4(n189), .O(
        read_data2[12]) );
  NAND_GATE U244 ( .I1(n74), .I2(\scp_reg[15][12] ), .O(n189) );
  NAND_GATE U245 ( .I1(n75), .I2(\scp_reg[14][12] ), .O(n188) );
  NAND_GATE U246 ( .I1(\scp_reg[13][12] ), .I2(n76), .O(n187) );
  NAND_GATE U247 ( .I1(\scp_reg[12][12] ), .I2(n77), .O(n186) );
  NAND4_GATE U248 ( .I1(n190), .I2(n191), .I3(n192), .I4(n193), .O(
        read_data2[11]) );
  NAND_GATE U249 ( .I1(n74), .I2(\scp_reg[15][11] ), .O(n193) );
  NAND_GATE U250 ( .I1(n75), .I2(\scp_reg[14][11] ), .O(n192) );
  NAND_GATE U251 ( .I1(\scp_reg[13][11] ), .I2(n76), .O(n191) );
  NAND_GATE U252 ( .I1(\scp_reg[12][11] ), .I2(n77), .O(n190) );
  NAND4_GATE U253 ( .I1(n194), .I2(n195), .I3(n196), .I4(n197), .O(
        read_data2[10]) );
  NAND_GATE U254 ( .I1(n74), .I2(\scp_reg[15][10] ), .O(n197) );
  NAND_GATE U255 ( .I1(n75), .I2(\scp_reg[14][10] ), .O(n196) );
  NAND_GATE U256 ( .I1(\scp_reg[13][10] ), .I2(n76), .O(n195) );
  NAND_GATE U257 ( .I1(\scp_reg[12][10] ), .I2(n77), .O(n194) );
  NAND4_GATE U258 ( .I1(n198), .I2(n199), .I3(n200), .I4(n201), .O(
        read_data2[0]) );
  NAND_GATE U259 ( .I1(n74), .I2(\scp_reg[15][0] ), .O(n201) );
  AND3_GATE U260 ( .I1(read_adr2[0]), .I2(n202), .I3(read_adr2[1]), .O(n74) );
  NAND_GATE U261 ( .I1(n75), .I2(\scp_reg[14][0] ), .O(n200) );
  AND3_GATE U262 ( .I1(n202), .I2(n203), .I3(read_adr2[1]), .O(n75) );
  NAND_GATE U263 ( .I1(\scp_reg[13][0] ), .I2(n76), .O(n199) );
  AND3_GATE U264 ( .I1(n202), .I2(n204), .I3(read_adr2[0]), .O(n76) );
  NAND_GATE U265 ( .I1(n77), .I2(\scp_reg[12][0] ), .O(n198) );
  AND3_GATE U266 ( .I1(n203), .I2(n204), .I3(n202), .O(n77) );
  AND3_GATE U267 ( .I1(read_adr2[2]), .I2(n205), .I3(read_adr2[3]), .O(n202)
         );
  INV_GATE U268 ( .I1(N72), .O(n205) );
  INV_GATE U269 ( .I1(read_adr2[1]), .O(n204) );
  INV_GATE U270 ( .I1(read_adr2[0]), .O(n203) );
  NAND4_GATE U271 ( .I1(n206), .I2(n207), .I3(n208), .I4(n209), .O(
        read_data1[9]) );
  NAND_GATE U272 ( .I1(n210), .I2(\scp_reg[15][9] ), .O(n209) );
  NAND_GATE U273 ( .I1(n211), .I2(\scp_reg[14][9] ), .O(n208) );
  NAND_GATE U274 ( .I1(n212), .I2(\scp_reg[13][9] ), .O(n207) );
  NAND_GATE U275 ( .I1(n213), .I2(\scp_reg[12][9] ), .O(n206) );
  NAND4_GATE U276 ( .I1(n214), .I2(n215), .I3(n216), .I4(n217), .O(
        read_data1[8]) );
  NAND_GATE U277 ( .I1(n210), .I2(\scp_reg[15][8] ), .O(n217) );
  NAND_GATE U278 ( .I1(n211), .I2(\scp_reg[14][8] ), .O(n216) );
  NAND_GATE U279 ( .I1(n212), .I2(\scp_reg[13][8] ), .O(n215) );
  NAND_GATE U280 ( .I1(n213), .I2(\scp_reg[12][8] ), .O(n214) );
  NAND4_GATE U281 ( .I1(n218), .I2(n219), .I3(n220), .I4(n221), .O(
        read_data1[7]) );
  NAND_GATE U282 ( .I1(n210), .I2(\scp_reg[15][7] ), .O(n221) );
  NAND_GATE U283 ( .I1(n211), .I2(\scp_reg[14][7] ), .O(n220) );
  NAND_GATE U284 ( .I1(n212), .I2(\scp_reg[13][7] ), .O(n219) );
  NAND_GATE U285 ( .I1(n213), .I2(\scp_reg[12][7] ), .O(n218) );
  NAND4_GATE U286 ( .I1(n222), .I2(n223), .I3(n224), .I4(n225), .O(
        read_data1[6]) );
  NAND_GATE U287 ( .I1(n210), .I2(\scp_reg[15][6] ), .O(n225) );
  NAND_GATE U288 ( .I1(n211), .I2(\scp_reg[14][6] ), .O(n224) );
  NAND_GATE U289 ( .I1(n212), .I2(\scp_reg[13][6] ), .O(n223) );
  NAND_GATE U290 ( .I1(n213), .I2(\scp_reg[12][6] ), .O(n222) );
  NAND4_GATE U291 ( .I1(n226), .I2(n227), .I3(n228), .I4(n229), .O(
        read_data1[5]) );
  NAND_GATE U292 ( .I1(n210), .I2(\scp_reg[15][5] ), .O(n229) );
  NAND_GATE U293 ( .I1(n211), .I2(\scp_reg[14][5] ), .O(n228) );
  NAND_GATE U294 ( .I1(n212), .I2(\scp_reg[13][5] ), .O(n227) );
  NAND_GATE U295 ( .I1(n213), .I2(\scp_reg[12][5] ), .O(n226) );
  NAND4_GATE U296 ( .I1(n230), .I2(n231), .I3(n232), .I4(n233), .O(
        read_data1[4]) );
  NAND_GATE U297 ( .I1(n210), .I2(\scp_reg[15][4] ), .O(n233) );
  NAND_GATE U298 ( .I1(n211), .I2(\scp_reg[14][4] ), .O(n232) );
  NAND_GATE U299 ( .I1(n212), .I2(\scp_reg[13][4] ), .O(n231) );
  NAND_GATE U300 ( .I1(n213), .I2(\scp_reg[12][4] ), .O(n230) );
  NAND4_GATE U301 ( .I1(n234), .I2(n235), .I3(n236), .I4(n237), .O(
        read_data1[3]) );
  NAND_GATE U302 ( .I1(n210), .I2(\scp_reg[15][3] ), .O(n237) );
  NAND_GATE U303 ( .I1(n211), .I2(\scp_reg[14][3] ), .O(n236) );
  NAND_GATE U304 ( .I1(n212), .I2(\scp_reg[13][3] ), .O(n235) );
  NAND_GATE U305 ( .I1(n213), .I2(\scp_reg[12][3] ), .O(n234) );
  NAND4_GATE U306 ( .I1(n238), .I2(n239), .I3(n240), .I4(n241), .O(
        read_data1[31]) );
  NAND_GATE U307 ( .I1(n210), .I2(\scp_reg[15][31] ), .O(n241) );
  NAND_GATE U308 ( .I1(n211), .I2(\scp_reg[14][31] ), .O(n240) );
  NAND_GATE U309 ( .I1(n212), .I2(\scp_reg[13][31] ), .O(n239) );
  NAND_GATE U310 ( .I1(n213), .I2(\scp_reg[12][31] ), .O(n238) );
  NAND4_GATE U311 ( .I1(n242), .I2(n243), .I3(n244), .I4(n245), .O(
        read_data1[30]) );
  NAND_GATE U312 ( .I1(n210), .I2(\scp_reg[15][30] ), .O(n245) );
  NAND_GATE U313 ( .I1(n211), .I2(\scp_reg[14][30] ), .O(n244) );
  NAND_GATE U314 ( .I1(n212), .I2(\scp_reg[13][30] ), .O(n243) );
  NAND_GATE U315 ( .I1(n213), .I2(\scp_reg[12][30] ), .O(n242) );
  NAND4_GATE U316 ( .I1(n246), .I2(n247), .I3(n248), .I4(n249), .O(
        read_data1[2]) );
  NAND_GATE U317 ( .I1(n210), .I2(\scp_reg[15][2] ), .O(n249) );
  NAND_GATE U318 ( .I1(n211), .I2(\scp_reg[14][2] ), .O(n248) );
  NAND_GATE U319 ( .I1(n212), .I2(\scp_reg[13][2] ), .O(n247) );
  NAND_GATE U320 ( .I1(n213), .I2(\scp_reg[12][2] ), .O(n246) );
  NAND4_GATE U321 ( .I1(n250), .I2(n251), .I3(n252), .I4(n253), .O(
        read_data1[29]) );
  NAND_GATE U322 ( .I1(n210), .I2(\scp_reg[15][29] ), .O(n253) );
  NAND_GATE U323 ( .I1(n211), .I2(\scp_reg[14][29] ), .O(n252) );
  NAND_GATE U324 ( .I1(n212), .I2(\scp_reg[13][29] ), .O(n251) );
  NAND_GATE U325 ( .I1(n213), .I2(\scp_reg[12][29] ), .O(n250) );
  NAND4_GATE U326 ( .I1(n254), .I2(n255), .I3(n256), .I4(n257), .O(
        read_data1[28]) );
  NAND_GATE U327 ( .I1(n210), .I2(\scp_reg[15][28] ), .O(n257) );
  NAND_GATE U328 ( .I1(n211), .I2(\scp_reg[14][28] ), .O(n256) );
  NAND_GATE U329 ( .I1(n212), .I2(\scp_reg[13][28] ), .O(n255) );
  NAND_GATE U330 ( .I1(n213), .I2(\scp_reg[12][28] ), .O(n254) );
  NAND4_GATE U331 ( .I1(n258), .I2(n259), .I3(n260), .I4(n261), .O(
        read_data1[27]) );
  NAND_GATE U332 ( .I1(n210), .I2(\scp_reg[15][27] ), .O(n261) );
  NAND_GATE U333 ( .I1(n211), .I2(\scp_reg[14][27] ), .O(n260) );
  NAND_GATE U334 ( .I1(n212), .I2(\scp_reg[13][27] ), .O(n259) );
  NAND_GATE U335 ( .I1(n213), .I2(\scp_reg[12][27] ), .O(n258) );
  NAND4_GATE U336 ( .I1(n262), .I2(n263), .I3(n264), .I4(n265), .O(
        read_data1[26]) );
  NAND_GATE U337 ( .I1(n210), .I2(\scp_reg[15][26] ), .O(n265) );
  NAND_GATE U338 ( .I1(n211), .I2(\scp_reg[14][26] ), .O(n264) );
  NAND_GATE U339 ( .I1(n212), .I2(\scp_reg[13][26] ), .O(n263) );
  NAND_GATE U340 ( .I1(n213), .I2(\scp_reg[12][26] ), .O(n262) );
  NAND4_GATE U341 ( .I1(n266), .I2(n267), .I3(n268), .I4(n269), .O(
        read_data1[25]) );
  NAND_GATE U342 ( .I1(n210), .I2(\scp_reg[15][25] ), .O(n269) );
  NAND_GATE U343 ( .I1(n211), .I2(\scp_reg[14][25] ), .O(n268) );
  NAND_GATE U344 ( .I1(n212), .I2(\scp_reg[13][25] ), .O(n267) );
  NAND_GATE U345 ( .I1(n213), .I2(\scp_reg[12][25] ), .O(n266) );
  NAND4_GATE U346 ( .I1(n270), .I2(n271), .I3(n272), .I4(n273), .O(
        read_data1[24]) );
  NAND_GATE U347 ( .I1(n210), .I2(\scp_reg[15][24] ), .O(n273) );
  NAND_GATE U348 ( .I1(n211), .I2(\scp_reg[14][24] ), .O(n272) );
  NAND_GATE U349 ( .I1(n212), .I2(\scp_reg[13][24] ), .O(n271) );
  NAND_GATE U350 ( .I1(n213), .I2(\scp_reg[12][24] ), .O(n270) );
  NAND4_GATE U351 ( .I1(n274), .I2(n275), .I3(n276), .I4(n277), .O(
        read_data1[23]) );
  NAND_GATE U352 ( .I1(n210), .I2(\scp_reg[15][23] ), .O(n277) );
  NAND_GATE U353 ( .I1(n211), .I2(\scp_reg[14][23] ), .O(n276) );
  NAND_GATE U354 ( .I1(n212), .I2(\scp_reg[13][23] ), .O(n275) );
  NAND_GATE U355 ( .I1(n213), .I2(\scp_reg[12][23] ), .O(n274) );
  NAND4_GATE U356 ( .I1(n278), .I2(n279), .I3(n280), .I4(n281), .O(
        read_data1[22]) );
  NAND_GATE U357 ( .I1(n210), .I2(\scp_reg[15][22] ), .O(n281) );
  NAND_GATE U358 ( .I1(n211), .I2(\scp_reg[14][22] ), .O(n280) );
  NAND_GATE U359 ( .I1(n212), .I2(\scp_reg[13][22] ), .O(n279) );
  NAND_GATE U360 ( .I1(n213), .I2(\scp_reg[12][22] ), .O(n278) );
  NAND4_GATE U361 ( .I1(n282), .I2(n283), .I3(n284), .I4(n285), .O(
        read_data1[21]) );
  NAND_GATE U362 ( .I1(n210), .I2(\scp_reg[15][21] ), .O(n285) );
  NAND_GATE U363 ( .I1(n211), .I2(\scp_reg[14][21] ), .O(n284) );
  NAND_GATE U364 ( .I1(n212), .I2(\scp_reg[13][21] ), .O(n283) );
  NAND_GATE U365 ( .I1(n213), .I2(\scp_reg[12][21] ), .O(n282) );
  NAND4_GATE U366 ( .I1(n286), .I2(n287), .I3(n288), .I4(n289), .O(
        read_data1[20]) );
  NAND_GATE U367 ( .I1(n210), .I2(\scp_reg[15][20] ), .O(n289) );
  NAND_GATE U368 ( .I1(n211), .I2(\scp_reg[14][20] ), .O(n288) );
  NAND_GATE U369 ( .I1(n212), .I2(\scp_reg[13][20] ), .O(n287) );
  NAND_GATE U370 ( .I1(n213), .I2(\scp_reg[12][20] ), .O(n286) );
  NAND4_GATE U371 ( .I1(n290), .I2(n291), .I3(n292), .I4(n293), .O(
        read_data1[1]) );
  NAND_GATE U372 ( .I1(n210), .I2(\scp_reg[15][1] ), .O(n293) );
  NAND_GATE U373 ( .I1(n211), .I2(\scp_reg[14][1] ), .O(n292) );
  NAND_GATE U374 ( .I1(n212), .I2(\scp_reg[13][1] ), .O(n291) );
  NAND_GATE U375 ( .I1(n213), .I2(\scp_reg[12][1] ), .O(n290) );
  NAND4_GATE U376 ( .I1(n294), .I2(n295), .I3(n296), .I4(n297), .O(
        read_data1[19]) );
  NAND_GATE U377 ( .I1(n210), .I2(\scp_reg[15][19] ), .O(n297) );
  NAND_GATE U378 ( .I1(n211), .I2(\scp_reg[14][19] ), .O(n296) );
  NAND_GATE U379 ( .I1(n212), .I2(\scp_reg[13][19] ), .O(n295) );
  NAND_GATE U380 ( .I1(n213), .I2(\scp_reg[12][19] ), .O(n294) );
  NAND4_GATE U381 ( .I1(n298), .I2(n299), .I3(n300), .I4(n301), .O(
        read_data1[18]) );
  NAND_GATE U382 ( .I1(n210), .I2(\scp_reg[15][18] ), .O(n301) );
  NAND_GATE U383 ( .I1(n211), .I2(\scp_reg[14][18] ), .O(n300) );
  NAND_GATE U384 ( .I1(n212), .I2(\scp_reg[13][18] ), .O(n299) );
  NAND_GATE U385 ( .I1(n213), .I2(\scp_reg[12][18] ), .O(n298) );
  NAND4_GATE U386 ( .I1(n302), .I2(n303), .I3(n304), .I4(n305), .O(
        read_data1[17]) );
  NAND_GATE U387 ( .I1(n210), .I2(\scp_reg[15][17] ), .O(n305) );
  NAND_GATE U388 ( .I1(n211), .I2(\scp_reg[14][17] ), .O(n304) );
  NAND_GATE U389 ( .I1(n212), .I2(\scp_reg[13][17] ), .O(n303) );
  NAND_GATE U390 ( .I1(n213), .I2(\scp_reg[12][17] ), .O(n302) );
  NAND4_GATE U391 ( .I1(n306), .I2(n307), .I3(n308), .I4(n309), .O(
        read_data1[16]) );
  NAND_GATE U392 ( .I1(n210), .I2(\scp_reg[15][16] ), .O(n309) );
  NAND_GATE U393 ( .I1(n211), .I2(\scp_reg[14][16] ), .O(n308) );
  NAND_GATE U394 ( .I1(n212), .I2(\scp_reg[13][16] ), .O(n307) );
  NAND_GATE U395 ( .I1(n213), .I2(\scp_reg[12][16] ), .O(n306) );
  NAND4_GATE U396 ( .I1(n310), .I2(n311), .I3(n312), .I4(n313), .O(
        read_data1[15]) );
  NAND_GATE U397 ( .I1(n210), .I2(\scp_reg[15][15] ), .O(n313) );
  NAND_GATE U398 ( .I1(n211), .I2(\scp_reg[14][15] ), .O(n312) );
  NAND_GATE U399 ( .I1(n212), .I2(\scp_reg[13][15] ), .O(n311) );
  NAND_GATE U400 ( .I1(n213), .I2(\scp_reg[12][15] ), .O(n310) );
  NAND4_GATE U401 ( .I1(n314), .I2(n315), .I3(n316), .I4(n317), .O(
        read_data1[14]) );
  NAND_GATE U402 ( .I1(n210), .I2(\scp_reg[15][14] ), .O(n317) );
  NAND_GATE U403 ( .I1(n211), .I2(\scp_reg[14][14] ), .O(n316) );
  NAND_GATE U404 ( .I1(n212), .I2(\scp_reg[13][14] ), .O(n315) );
  NAND_GATE U405 ( .I1(n213), .I2(\scp_reg[12][14] ), .O(n314) );
  NAND4_GATE U406 ( .I1(n318), .I2(n319), .I3(n320), .I4(n321), .O(
        read_data1[13]) );
  NAND_GATE U407 ( .I1(n210), .I2(\scp_reg[15][13] ), .O(n321) );
  NAND_GATE U408 ( .I1(n211), .I2(\scp_reg[14][13] ), .O(n320) );
  NAND_GATE U409 ( .I1(n212), .I2(\scp_reg[13][13] ), .O(n319) );
  NAND_GATE U410 ( .I1(n213), .I2(\scp_reg[12][13] ), .O(n318) );
  NAND4_GATE U411 ( .I1(n322), .I2(n323), .I3(n324), .I4(n325), .O(
        read_data1[12]) );
  NAND_GATE U412 ( .I1(n210), .I2(\scp_reg[15][12] ), .O(n325) );
  NAND_GATE U413 ( .I1(n211), .I2(\scp_reg[14][12] ), .O(n324) );
  NAND_GATE U414 ( .I1(n212), .I2(\scp_reg[13][12] ), .O(n323) );
  NAND_GATE U415 ( .I1(n213), .I2(\scp_reg[12][12] ), .O(n322) );
  NAND4_GATE U416 ( .I1(n326), .I2(n327), .I3(n328), .I4(n329), .O(
        read_data1[11]) );
  NAND_GATE U417 ( .I1(n210), .I2(\scp_reg[15][11] ), .O(n329) );
  NAND_GATE U418 ( .I1(n211), .I2(\scp_reg[14][11] ), .O(n328) );
  NAND_GATE U419 ( .I1(n212), .I2(\scp_reg[13][11] ), .O(n327) );
  NAND_GATE U420 ( .I1(n213), .I2(\scp_reg[12][11] ), .O(n326) );
  NAND4_GATE U421 ( .I1(n330), .I2(n331), .I3(n332), .I4(n333), .O(
        read_data1[10]) );
  NAND_GATE U422 ( .I1(n210), .I2(\scp_reg[15][10] ), .O(n333) );
  NAND_GATE U423 ( .I1(n211), .I2(\scp_reg[14][10] ), .O(n332) );
  NAND_GATE U424 ( .I1(n212), .I2(\scp_reg[13][10] ), .O(n331) );
  NAND_GATE U425 ( .I1(n213), .I2(\scp_reg[12][10] ), .O(n330) );
  NAND4_GATE U426 ( .I1(n334), .I2(n335), .I3(n336), .I4(n337), .O(
        read_data1[0]) );
  NAND_GATE U427 ( .I1(n210), .I2(\scp_reg[15][0] ), .O(n337) );
  AND3_GATE U428 ( .I1(read_adr1[0]), .I2(n338), .I3(read_adr1[1]), .O(n210)
         );
  NAND_GATE U429 ( .I1(n211), .I2(\scp_reg[14][0] ), .O(n336) );
  AND3_GATE U430 ( .I1(n338), .I2(n339), .I3(read_adr1[1]), .O(n211) );
  NAND_GATE U431 ( .I1(n212), .I2(\scp_reg[13][0] ), .O(n335) );
  AND3_GATE U432 ( .I1(n338), .I2(n340), .I3(read_adr1[0]), .O(n212) );
  NAND_GATE U433 ( .I1(n213), .I2(\scp_reg[12][0] ), .O(n334) );
  AND3_GATE U434 ( .I1(n339), .I2(n340), .I3(n338), .O(n213) );
  AND3_GATE U435 ( .I1(read_adr1[2]), .I2(n341), .I3(read_adr1[3]), .O(n338)
         );
  INV_GATE U436 ( .I1(N30), .O(n341) );
  INV_GATE U437 ( .I1(read_adr1[1]), .O(n340) );
  INV_GATE U438 ( .I1(read_adr1[0]), .O(n339) );
  NAND3_GATE U439 ( .I1(n342), .I2(n343), .I3(n344), .O(\pre_reg[14][9] ) );
  NAND_GATE U440 ( .I1(n345), .I2(\scp_reg[14][9] ), .O(n344) );
  NAND_GATE U441 ( .I1(MEM_adr[9]), .I2(n346), .O(n343) );
  NAND_GATE U442 ( .I1(write_data[9]), .I2(n347), .O(n342) );
  NAND3_GATE U443 ( .I1(n348), .I2(n349), .I3(n350), .O(\pre_reg[14][8] ) );
  NAND_GATE U444 ( .I1(n345), .I2(\scp_reg[14][8] ), .O(n350) );
  NAND_GATE U445 ( .I1(MEM_adr[8]), .I2(n346), .O(n349) );
  NAND_GATE U446 ( .I1(write_data[8]), .I2(n347), .O(n348) );
  NAND3_GATE U447 ( .I1(n351), .I2(n352), .I3(n353), .O(\pre_reg[14][7] ) );
  NAND_GATE U448 ( .I1(n345), .I2(\scp_reg[14][7] ), .O(n353) );
  NAND_GATE U449 ( .I1(MEM_adr[7]), .I2(n346), .O(n352) );
  NAND_GATE U450 ( .I1(write_data[7]), .I2(n347), .O(n351) );
  NAND3_GATE U451 ( .I1(n354), .I2(n355), .I3(n356), .O(\pre_reg[14][6] ) );
  NAND_GATE U452 ( .I1(n345), .I2(\scp_reg[14][6] ), .O(n356) );
  NAND_GATE U453 ( .I1(MEM_adr[6]), .I2(n346), .O(n355) );
  NAND_GATE U454 ( .I1(write_data[6]), .I2(n347), .O(n354) );
  NAND3_GATE U455 ( .I1(n357), .I2(n358), .I3(n359), .O(\pre_reg[14][5] ) );
  NAND_GATE U456 ( .I1(n345), .I2(\scp_reg[14][5] ), .O(n359) );
  NAND_GATE U457 ( .I1(MEM_adr[5]), .I2(n346), .O(n358) );
  NAND_GATE U458 ( .I1(write_data[5]), .I2(n347), .O(n357) );
  NAND3_GATE U459 ( .I1(n360), .I2(n361), .I3(n362), .O(\pre_reg[14][4] ) );
  NAND_GATE U460 ( .I1(n345), .I2(\scp_reg[14][4] ), .O(n362) );
  NAND_GATE U461 ( .I1(MEM_adr[4]), .I2(n346), .O(n361) );
  NAND_GATE U462 ( .I1(write_data[4]), .I2(n347), .O(n360) );
  NAND3_GATE U463 ( .I1(n363), .I2(n364), .I3(n365), .O(\pre_reg[14][3] ) );
  NAND_GATE U464 ( .I1(n345), .I2(\scp_reg[14][3] ), .O(n365) );
  NAND_GATE U465 ( .I1(MEM_adr[3]), .I2(n346), .O(n364) );
  NAND_GATE U466 ( .I1(write_data[3]), .I2(n347), .O(n363) );
  NAND3_GATE U467 ( .I1(n366), .I2(n367), .I3(n368), .O(\pre_reg[14][31] ) );
  NAND_GATE U468 ( .I1(n345), .I2(\scp_reg[14][31] ), .O(n368) );
  NAND_GATE U469 ( .I1(MEM_adr[31]), .I2(n346), .O(n367) );
  NAND_GATE U470 ( .I1(write_data[31]), .I2(n347), .O(n366) );
  NAND3_GATE U471 ( .I1(n369), .I2(n370), .I3(n371), .O(\pre_reg[14][30] ) );
  NAND_GATE U472 ( .I1(n345), .I2(\scp_reg[14][30] ), .O(n371) );
  NAND_GATE U473 ( .I1(MEM_adr[30]), .I2(n346), .O(n370) );
  NAND_GATE U474 ( .I1(write_data[30]), .I2(n347), .O(n369) );
  NAND3_GATE U475 ( .I1(n372), .I2(n373), .I3(n374), .O(\pre_reg[14][2] ) );
  NAND_GATE U476 ( .I1(n345), .I2(\scp_reg[14][2] ), .O(n374) );
  NAND_GATE U477 ( .I1(MEM_adr[2]), .I2(n346), .O(n373) );
  NAND_GATE U478 ( .I1(n347), .I2(write_data[2]), .O(n372) );
  NAND3_GATE U479 ( .I1(n375), .I2(n376), .I3(n377), .O(\pre_reg[14][29] ) );
  NAND_GATE U480 ( .I1(n345), .I2(\scp_reg[14][29] ), .O(n377) );
  NAND_GATE U481 ( .I1(MEM_adr[29]), .I2(n346), .O(n376) );
  NAND_GATE U482 ( .I1(write_data[29]), .I2(n347), .O(n375) );
  NAND3_GATE U483 ( .I1(n378), .I2(n379), .I3(n380), .O(\pre_reg[14][28] ) );
  NAND_GATE U484 ( .I1(n345), .I2(\scp_reg[14][28] ), .O(n380) );
  NAND_GATE U485 ( .I1(MEM_adr[28]), .I2(n346), .O(n379) );
  NAND_GATE U486 ( .I1(write_data[28]), .I2(n347), .O(n378) );
  NAND3_GATE U487 ( .I1(n381), .I2(n382), .I3(n383), .O(\pre_reg[14][27] ) );
  NAND_GATE U488 ( .I1(n345), .I2(\scp_reg[14][27] ), .O(n383) );
  NAND_GATE U489 ( .I1(MEM_adr[27]), .I2(n346), .O(n382) );
  NAND_GATE U490 ( .I1(write_data[27]), .I2(n347), .O(n381) );
  NAND3_GATE U491 ( .I1(n384), .I2(n385), .I3(n386), .O(\pre_reg[14][26] ) );
  NAND_GATE U492 ( .I1(n345), .I2(\scp_reg[14][26] ), .O(n386) );
  NAND_GATE U493 ( .I1(MEM_adr[26]), .I2(n346), .O(n385) );
  NAND_GATE U494 ( .I1(write_data[26]), .I2(n347), .O(n384) );
  NAND3_GATE U495 ( .I1(n387), .I2(n388), .I3(n389), .O(\pre_reg[14][25] ) );
  NAND_GATE U496 ( .I1(n345), .I2(\scp_reg[14][25] ), .O(n389) );
  NAND_GATE U497 ( .I1(MEM_adr[25]), .I2(n346), .O(n388) );
  NAND_GATE U498 ( .I1(write_data[25]), .I2(n347), .O(n387) );
  NAND3_GATE U499 ( .I1(n390), .I2(n391), .I3(n392), .O(\pre_reg[14][24] ) );
  NAND_GATE U500 ( .I1(n345), .I2(\scp_reg[14][24] ), .O(n392) );
  NAND_GATE U501 ( .I1(MEM_adr[24]), .I2(n346), .O(n391) );
  NAND_GATE U502 ( .I1(write_data[24]), .I2(n347), .O(n390) );
  NAND3_GATE U503 ( .I1(n393), .I2(n394), .I3(n395), .O(\pre_reg[14][23] ) );
  NAND_GATE U504 ( .I1(n345), .I2(\scp_reg[14][23] ), .O(n395) );
  NAND_GATE U505 ( .I1(MEM_adr[23]), .I2(n346), .O(n394) );
  NAND_GATE U506 ( .I1(write_data[23]), .I2(n347), .O(n393) );
  NAND3_GATE U507 ( .I1(n396), .I2(n397), .I3(n398), .O(\pre_reg[14][22] ) );
  NAND_GATE U508 ( .I1(n345), .I2(\scp_reg[14][22] ), .O(n398) );
  NAND_GATE U509 ( .I1(MEM_adr[22]), .I2(n346), .O(n397) );
  NAND_GATE U510 ( .I1(write_data[22]), .I2(n347), .O(n396) );
  NAND3_GATE U511 ( .I1(n399), .I2(n400), .I3(n401), .O(\pre_reg[14][21] ) );
  NAND_GATE U512 ( .I1(n345), .I2(\scp_reg[14][21] ), .O(n401) );
  NAND_GATE U513 ( .I1(MEM_adr[21]), .I2(n346), .O(n400) );
  NAND_GATE U514 ( .I1(write_data[21]), .I2(n347), .O(n399) );
  NAND3_GATE U515 ( .I1(n402), .I2(n403), .I3(n404), .O(\pre_reg[14][20] ) );
  NAND_GATE U516 ( .I1(n345), .I2(\scp_reg[14][20] ), .O(n404) );
  NAND_GATE U517 ( .I1(MEM_adr[20]), .I2(n346), .O(n403) );
  NAND_GATE U518 ( .I1(write_data[20]), .I2(n347), .O(n402) );
  NAND3_GATE U519 ( .I1(n405), .I2(n406), .I3(n407), .O(\pre_reg[14][1] ) );
  NAND_GATE U520 ( .I1(n345), .I2(\scp_reg[14][1] ), .O(n407) );
  NAND_GATE U521 ( .I1(MEM_adr[1]), .I2(n346), .O(n406) );
  NAND_GATE U522 ( .I1(write_data[1]), .I2(n347), .O(n405) );
  NAND3_GATE U523 ( .I1(n408), .I2(n409), .I3(n410), .O(\pre_reg[14][19] ) );
  NAND_GATE U524 ( .I1(n345), .I2(\scp_reg[14][19] ), .O(n410) );
  NAND_GATE U525 ( .I1(MEM_adr[19]), .I2(n346), .O(n409) );
  NAND_GATE U526 ( .I1(write_data[19]), .I2(n347), .O(n408) );
  NAND3_GATE U527 ( .I1(n411), .I2(n412), .I3(n413), .O(\pre_reg[14][18] ) );
  NAND_GATE U528 ( .I1(n345), .I2(\scp_reg[14][18] ), .O(n413) );
  NAND_GATE U529 ( .I1(MEM_adr[18]), .I2(n346), .O(n412) );
  NAND_GATE U530 ( .I1(write_data[18]), .I2(n347), .O(n411) );
  NAND3_GATE U531 ( .I1(n414), .I2(n415), .I3(n416), .O(\pre_reg[14][17] ) );
  NAND_GATE U532 ( .I1(n345), .I2(\scp_reg[14][17] ), .O(n416) );
  NAND_GATE U533 ( .I1(MEM_adr[17]), .I2(n346), .O(n415) );
  NAND_GATE U534 ( .I1(write_data[17]), .I2(n347), .O(n414) );
  NAND3_GATE U535 ( .I1(n417), .I2(n418), .I3(n419), .O(\pre_reg[14][16] ) );
  NAND_GATE U536 ( .I1(n345), .I2(\scp_reg[14][16] ), .O(n419) );
  NAND_GATE U537 ( .I1(MEM_adr[16]), .I2(n346), .O(n418) );
  NAND_GATE U538 ( .I1(write_data[16]), .I2(n347), .O(n417) );
  NAND3_GATE U539 ( .I1(n420), .I2(n421), .I3(n422), .O(\pre_reg[14][15] ) );
  NAND_GATE U540 ( .I1(n345), .I2(\scp_reg[14][15] ), .O(n422) );
  NAND_GATE U541 ( .I1(MEM_adr[15]), .I2(n346), .O(n421) );
  NAND_GATE U542 ( .I1(write_data[15]), .I2(n347), .O(n420) );
  NAND3_GATE U543 ( .I1(n423), .I2(n424), .I3(n425), .O(\pre_reg[14][14] ) );
  NAND_GATE U544 ( .I1(n345), .I2(\scp_reg[14][14] ), .O(n425) );
  NAND_GATE U545 ( .I1(MEM_adr[14]), .I2(n346), .O(n424) );
  NAND_GATE U546 ( .I1(write_data[14]), .I2(n347), .O(n423) );
  NAND3_GATE U547 ( .I1(n426), .I2(n427), .I3(n428), .O(\pre_reg[14][13] ) );
  NAND_GATE U548 ( .I1(n345), .I2(\scp_reg[14][13] ), .O(n428) );
  NAND_GATE U549 ( .I1(MEM_adr[13]), .I2(n346), .O(n427) );
  NAND_GATE U550 ( .I1(write_data[13]), .I2(n347), .O(n426) );
  NAND3_GATE U551 ( .I1(n429), .I2(n430), .I3(n431), .O(\pre_reg[14][12] ) );
  NAND_GATE U552 ( .I1(n345), .I2(\scp_reg[14][12] ), .O(n431) );
  NAND_GATE U553 ( .I1(MEM_adr[12]), .I2(n346), .O(n430) );
  NAND_GATE U554 ( .I1(write_data[12]), .I2(n347), .O(n429) );
  NAND3_GATE U555 ( .I1(n432), .I2(n433), .I3(n434), .O(\pre_reg[14][11] ) );
  NAND_GATE U556 ( .I1(n345), .I2(\scp_reg[14][11] ), .O(n434) );
  NAND_GATE U557 ( .I1(MEM_adr[11]), .I2(n346), .O(n433) );
  NAND_GATE U558 ( .I1(write_data[11]), .I2(n347), .O(n432) );
  NAND3_GATE U559 ( .I1(n435), .I2(n436), .I3(n437), .O(\pre_reg[14][10] ) );
  NAND_GATE U560 ( .I1(n345), .I2(\scp_reg[14][10] ), .O(n437) );
  NAND_GATE U561 ( .I1(MEM_adr[10]), .I2(n346), .O(n436) );
  NAND_GATE U562 ( .I1(write_data[10]), .I2(n347), .O(n435) );
  NAND3_GATE U563 ( .I1(n438), .I2(n439), .I3(n440), .O(\pre_reg[14][0] ) );
  NAND_GATE U564 ( .I1(n345), .I2(\scp_reg[14][0] ), .O(n440) );
  AND_GATE U565 ( .I1(n441), .I2(n442), .O(n345) );
  NAND_GATE U566 ( .I1(n443), .I2(n444), .O(n442) );
  NAND_GATE U567 ( .I1(MEM_adr[0]), .I2(n346), .O(n439) );
  AND_GATE U568 ( .I1(interrupt), .I2(n4), .O(n346) );
  NAND_GATE U569 ( .I1(write_data[0]), .I2(n347), .O(n438) );
  AND3_GATE U570 ( .I1(n443), .I2(n444), .I3(n441), .O(n347) );
  NAND3_GATE U571 ( .I1(n445), .I2(n446), .I3(n447), .O(\pre_reg[13][9] ) );
  NAND_GATE U572 ( .I1(MEM_exc_cause[9]), .I2(n4), .O(n447) );
  NAND_GATE U573 ( .I1(n448), .I2(write_data[9]), .O(n446) );
  NAND_GATE U574 ( .I1(n449), .I2(\scp_reg[13][9] ), .O(n445) );
  NAND3_GATE U575 ( .I1(n450), .I2(n451), .I3(n452), .O(\pre_reg[13][8] ) );
  NAND_GATE U576 ( .I1(MEM_exc_cause[8]), .I2(n4), .O(n452) );
  NAND_GATE U577 ( .I1(n448), .I2(write_data[8]), .O(n451) );
  NAND_GATE U578 ( .I1(n449), .I2(\scp_reg[13][8] ), .O(n450) );
  NAND3_GATE U579 ( .I1(n453), .I2(n454), .I3(n455), .O(\pre_reg[13][7] ) );
  NAND_GATE U580 ( .I1(MEM_exc_cause[7]), .I2(n4), .O(n455) );
  NAND_GATE U581 ( .I1(n448), .I2(write_data[7]), .O(n454) );
  NAND_GATE U582 ( .I1(n449), .I2(\scp_reg[13][7] ), .O(n453) );
  NAND3_GATE U583 ( .I1(n456), .I2(n457), .I3(n458), .O(\pre_reg[13][6] ) );
  NAND_GATE U584 ( .I1(MEM_exc_cause[6]), .I2(n4), .O(n458) );
  NAND_GATE U585 ( .I1(n448), .I2(write_data[6]), .O(n457) );
  NAND_GATE U586 ( .I1(n449), .I2(\scp_reg[13][6] ), .O(n456) );
  NAND3_GATE U587 ( .I1(n459), .I2(n460), .I3(n461), .O(\pre_reg[13][5] ) );
  NAND_GATE U588 ( .I1(MEM_exc_cause[5]), .I2(n4), .O(n461) );
  NAND_GATE U589 ( .I1(n448), .I2(write_data[5]), .O(n460) );
  NAND_GATE U590 ( .I1(n449), .I2(\scp_reg[13][5] ), .O(n459) );
  NAND3_GATE U591 ( .I1(n462), .I2(n463), .I3(n464), .O(\pre_reg[13][4] ) );
  NAND_GATE U592 ( .I1(MEM_exc_cause[4]), .I2(n4), .O(n464) );
  NAND_GATE U593 ( .I1(n448), .I2(write_data[4]), .O(n463) );
  NAND_GATE U594 ( .I1(n449), .I2(\scp_reg[13][4] ), .O(n462) );
  NAND3_GATE U595 ( .I1(n465), .I2(n466), .I3(n467), .O(\pre_reg[13][3] ) );
  NAND_GATE U596 ( .I1(MEM_exc_cause[3]), .I2(n4), .O(n467) );
  NAND_GATE U597 ( .I1(n448), .I2(write_data[3]), .O(n466) );
  NAND_GATE U598 ( .I1(n449), .I2(\scp_reg[13][3] ), .O(n465) );
  NAND3_GATE U599 ( .I1(n468), .I2(n469), .I3(n470), .O(\pre_reg[13][31] ) );
  NAND_GATE U600 ( .I1(MEM_exc_cause[31]), .I2(n4), .O(n470) );
  NAND_GATE U601 ( .I1(n448), .I2(write_data[31]), .O(n469) );
  NAND_GATE U602 ( .I1(n449), .I2(\scp_reg[13][31] ), .O(n468) );
  NAND3_GATE U603 ( .I1(n471), .I2(n472), .I3(n473), .O(\pre_reg[13][30] ) );
  NAND_GATE U604 ( .I1(MEM_exc_cause[30]), .I2(n4), .O(n473) );
  NAND_GATE U605 ( .I1(n448), .I2(write_data[30]), .O(n472) );
  NAND_GATE U606 ( .I1(n449), .I2(\scp_reg[13][30] ), .O(n471) );
  NAND3_GATE U607 ( .I1(n474), .I2(n475), .I3(n476), .O(\pre_reg[13][2] ) );
  NAND_GATE U608 ( .I1(MEM_exc_cause[2]), .I2(n4), .O(n476) );
  NAND_GATE U609 ( .I1(n448), .I2(write_data[2]), .O(n475) );
  NAND_GATE U610 ( .I1(n449), .I2(\scp_reg[13][2] ), .O(n474) );
  NAND3_GATE U611 ( .I1(n477), .I2(n478), .I3(n479), .O(\pre_reg[13][29] ) );
  NAND_GATE U612 ( .I1(MEM_exc_cause[29]), .I2(n4), .O(n479) );
  NAND_GATE U613 ( .I1(n448), .I2(write_data[29]), .O(n478) );
  NAND_GATE U614 ( .I1(n449), .I2(\scp_reg[13][29] ), .O(n477) );
  NAND3_GATE U615 ( .I1(n480), .I2(n481), .I3(n482), .O(\pre_reg[13][28] ) );
  NAND_GATE U616 ( .I1(MEM_exc_cause[28]), .I2(n4), .O(n482) );
  NAND_GATE U617 ( .I1(n448), .I2(write_data[28]), .O(n481) );
  NAND_GATE U618 ( .I1(n449), .I2(\scp_reg[13][28] ), .O(n480) );
  NAND3_GATE U619 ( .I1(n483), .I2(n484), .I3(n485), .O(\pre_reg[13][27] ) );
  NAND_GATE U620 ( .I1(MEM_exc_cause[27]), .I2(n4), .O(n485) );
  NAND_GATE U621 ( .I1(n448), .I2(write_data[27]), .O(n484) );
  NAND_GATE U622 ( .I1(n449), .I2(\scp_reg[13][27] ), .O(n483) );
  NAND3_GATE U623 ( .I1(n486), .I2(n487), .I3(n488), .O(\pre_reg[13][26] ) );
  NAND_GATE U624 ( .I1(MEM_exc_cause[26]), .I2(n4), .O(n488) );
  NAND_GATE U625 ( .I1(n448), .I2(write_data[26]), .O(n487) );
  NAND_GATE U626 ( .I1(n449), .I2(\scp_reg[13][26] ), .O(n486) );
  NAND3_GATE U627 ( .I1(n489), .I2(n490), .I3(n491), .O(\pre_reg[13][25] ) );
  NAND_GATE U628 ( .I1(MEM_exc_cause[25]), .I2(n4), .O(n491) );
  NAND_GATE U629 ( .I1(n448), .I2(write_data[25]), .O(n490) );
  NAND_GATE U630 ( .I1(n449), .I2(\scp_reg[13][25] ), .O(n489) );
  NAND3_GATE U631 ( .I1(n492), .I2(n493), .I3(n494), .O(\pre_reg[13][24] ) );
  NAND_GATE U632 ( .I1(MEM_exc_cause[24]), .I2(n4), .O(n494) );
  NAND_GATE U633 ( .I1(n448), .I2(write_data[24]), .O(n493) );
  NAND_GATE U634 ( .I1(n449), .I2(\scp_reg[13][24] ), .O(n492) );
  NAND3_GATE U635 ( .I1(n495), .I2(n496), .I3(n497), .O(\pre_reg[13][23] ) );
  NAND_GATE U636 ( .I1(MEM_exc_cause[23]), .I2(n4), .O(n497) );
  NAND_GATE U637 ( .I1(n448), .I2(write_data[23]), .O(n496) );
  NAND_GATE U638 ( .I1(n449), .I2(\scp_reg[13][23] ), .O(n495) );
  NAND3_GATE U639 ( .I1(n498), .I2(n499), .I3(n500), .O(\pre_reg[13][22] ) );
  NAND_GATE U640 ( .I1(MEM_exc_cause[22]), .I2(n4), .O(n500) );
  NAND_GATE U641 ( .I1(n448), .I2(write_data[22]), .O(n499) );
  NAND_GATE U642 ( .I1(n449), .I2(\scp_reg[13][22] ), .O(n498) );
  NAND3_GATE U643 ( .I1(n501), .I2(n502), .I3(n503), .O(\pre_reg[13][21] ) );
  NAND_GATE U644 ( .I1(MEM_exc_cause[21]), .I2(n4), .O(n503) );
  NAND_GATE U645 ( .I1(n448), .I2(write_data[21]), .O(n502) );
  NAND_GATE U646 ( .I1(n449), .I2(\scp_reg[13][21] ), .O(n501) );
  NAND3_GATE U647 ( .I1(n504), .I2(n505), .I3(n506), .O(\pre_reg[13][20] ) );
  NAND_GATE U648 ( .I1(MEM_exc_cause[20]), .I2(n4), .O(n506) );
  NAND_GATE U649 ( .I1(n448), .I2(write_data[20]), .O(n505) );
  NAND_GATE U650 ( .I1(n449), .I2(\scp_reg[13][20] ), .O(n504) );
  NAND3_GATE U651 ( .I1(n507), .I2(n508), .I3(n509), .O(\pre_reg[13][1] ) );
  NAND_GATE U652 ( .I1(MEM_exc_cause[1]), .I2(n4), .O(n509) );
  NAND_GATE U653 ( .I1(n448), .I2(write_data[1]), .O(n508) );
  NAND_GATE U654 ( .I1(n449), .I2(\scp_reg[13][1] ), .O(n507) );
  NAND3_GATE U655 ( .I1(n510), .I2(n511), .I3(n512), .O(\pre_reg[13][19] ) );
  NAND_GATE U656 ( .I1(MEM_exc_cause[19]), .I2(n4), .O(n512) );
  NAND_GATE U657 ( .I1(n448), .I2(write_data[19]), .O(n511) );
  NAND_GATE U658 ( .I1(n449), .I2(\scp_reg[13][19] ), .O(n510) );
  NAND3_GATE U659 ( .I1(n513), .I2(n514), .I3(n515), .O(\pre_reg[13][18] ) );
  NAND_GATE U660 ( .I1(MEM_exc_cause[18]), .I2(n4), .O(n515) );
  NAND_GATE U661 ( .I1(n448), .I2(write_data[18]), .O(n514) );
  NAND_GATE U662 ( .I1(n449), .I2(\scp_reg[13][18] ), .O(n513) );
  NAND3_GATE U663 ( .I1(n516), .I2(n517), .I3(n518), .O(\pre_reg[13][17] ) );
  NAND_GATE U664 ( .I1(MEM_exc_cause[17]), .I2(n4), .O(n518) );
  NAND_GATE U665 ( .I1(n448), .I2(write_data[17]), .O(n517) );
  NAND_GATE U666 ( .I1(n449), .I2(\scp_reg[13][17] ), .O(n516) );
  NAND3_GATE U667 ( .I1(n519), .I2(n520), .I3(n521), .O(\pre_reg[13][16] ) );
  NAND_GATE U668 ( .I1(MEM_exc_cause[16]), .I2(n4), .O(n521) );
  NAND_GATE U669 ( .I1(n448), .I2(write_data[16]), .O(n520) );
  NAND_GATE U670 ( .I1(n449), .I2(\scp_reg[13][16] ), .O(n519) );
  NAND3_GATE U671 ( .I1(n522), .I2(n523), .I3(n524), .O(\pre_reg[13][15] ) );
  NAND_GATE U672 ( .I1(MEM_exc_cause[15]), .I2(n4), .O(n524) );
  NAND_GATE U673 ( .I1(n448), .I2(write_data[15]), .O(n523) );
  NAND_GATE U674 ( .I1(n449), .I2(\scp_reg[13][15] ), .O(n522) );
  NAND3_GATE U675 ( .I1(n525), .I2(n526), .I3(n527), .O(\pre_reg[13][14] ) );
  NAND_GATE U676 ( .I1(MEM_exc_cause[14]), .I2(n4), .O(n527) );
  NAND_GATE U677 ( .I1(n448), .I2(write_data[14]), .O(n526) );
  NAND_GATE U678 ( .I1(n449), .I2(\scp_reg[13][14] ), .O(n525) );
  NAND3_GATE U679 ( .I1(n528), .I2(n529), .I3(n530), .O(\pre_reg[13][13] ) );
  NAND_GATE U680 ( .I1(MEM_exc_cause[13]), .I2(n4), .O(n530) );
  NAND_GATE U681 ( .I1(n448), .I2(write_data[13]), .O(n529) );
  NAND_GATE U682 ( .I1(n449), .I2(\scp_reg[13][13] ), .O(n528) );
  NAND3_GATE U683 ( .I1(n531), .I2(n532), .I3(n533), .O(\pre_reg[13][12] ) );
  NAND_GATE U684 ( .I1(MEM_exc_cause[12]), .I2(n4), .O(n533) );
  NAND_GATE U685 ( .I1(n448), .I2(write_data[12]), .O(n532) );
  NAND_GATE U686 ( .I1(n449), .I2(\scp_reg[13][12] ), .O(n531) );
  NAND3_GATE U687 ( .I1(n534), .I2(n535), .I3(n536), .O(\pre_reg[13][11] ) );
  NAND_GATE U688 ( .I1(MEM_exc_cause[11]), .I2(n4), .O(n536) );
  NAND_GATE U689 ( .I1(n448), .I2(write_data[11]), .O(n535) );
  NAND_GATE U690 ( .I1(n449), .I2(\scp_reg[13][11] ), .O(n534) );
  NAND3_GATE U691 ( .I1(n537), .I2(n538), .I3(n539), .O(\pre_reg[13][10] ) );
  NAND_GATE U692 ( .I1(MEM_exc_cause[10]), .I2(n4), .O(n539) );
  NAND_GATE U693 ( .I1(n448), .I2(write_data[10]), .O(n538) );
  NOR_GATE U694 ( .I1(n540), .I2(n541), .O(n448) );
  INV_GATE U695 ( .I1(n441), .O(n541) );
  NAND_GATE U696 ( .I1(n449), .I2(\scp_reg[13][10] ), .O(n537) );
  AND_GATE U697 ( .I1(n441), .I2(n540), .O(n449) );
  AND_GATE U698 ( .I1(n542), .I2(n4), .O(\pre_reg[13][0] ) );
  OR_GATE U699 ( .I1(MEM_exc_cause[0]), .I2(n543), .O(n542) );
  AND_GATE U700 ( .I1(n544), .I2(n545), .O(n543) );
  NAND3_GATE U701 ( .I1(n546), .I2(n547), .I3(n548), .O(n545) );
  OR_GATE U702 ( .I1(n540), .I2(n2), .O(n547) );
  NAND_GATE U703 ( .I1(\scp_reg[13][0] ), .I2(n540), .O(n546) );
  NAND3_GATE U704 ( .I1(n549), .I2(n550), .I3(write_adr[0]), .O(n540) );
  AND_GATE U705 ( .I1(n441), .I2(n551), .O(\pre_reg[12][0] ) );
  NAND3_GATE U706 ( .I1(n552), .I2(n553), .I3(n554), .O(n551) );
  NAND_GATE U707 ( .I1(save_msk), .I2(n7), .O(n554) );
  NOR4_GATE U708 ( .I1(n3), .I2(n555), .I3(write_data[0]), .I4(write_data[1]), 
        .O(n7) );
  OR_GATE U709 ( .I1(n555), .I2(n556), .O(n553) );
  AND_GATE U710 ( .I1(n557), .I2(n558), .O(n556) );
  NAND3_GATE U711 ( .I1(n2), .I2(n3), .I3(write_data[1]), .O(n558) );
  NAND_GATE U712 ( .I1(\scp_reg[12][0] ), .I2(n559), .O(n557) );
  OR_GATE U713 ( .I1(n560), .I2(write_data[1]), .O(n559) );
  AND_GATE U714 ( .I1(n561), .I2(n562), .O(n560) );
  OR_GATE U715 ( .I1(n3), .I2(write_data[0]), .O(n562) );
  OR_GATE U716 ( .I1(n2), .I2(write_data[2]), .O(n561) );
  NAND_GATE U717 ( .I1(n563), .I2(n555), .O(n552) );
  NAND4_GATE U718 ( .I1(n564), .I2(n565), .I3(n566), .I4(n567), .O(n555) );
  NOR5_GATE U719 ( .I1(write_data[30]), .I2(write_data[31]), .I3(write_data[3]), .I4(write_data[4]), .I5(n568), .O(n567) );
  OR5_GATE U720 ( .I1(write_data[6]), .I2(write_data[5]), .I3(write_data[7]), 
        .I4(write_data[9]), .I5(write_data[8]), .O(n568) );
  NOR5_GATE U721 ( .I1(write_data[21]), .I2(write_data[22]), .I3(
        write_data[23]), .I4(write_data[24]), .I5(n569), .O(n566) );
  OR5_GATE U722 ( .I1(write_data[26]), .I2(write_data[25]), .I3(write_data[27]), .I4(write_data[29]), .I5(write_data[28]), .O(n569) );
  NOR5_GATE U723 ( .I1(write_data[12]), .I2(write_data[13]), .I3(
        write_data[14]), .I4(write_data[15]), .I5(n570), .O(n565) );
  OR5_GATE U724 ( .I1(write_data[17]), .I2(write_data[16]), .I3(write_data[18]), .I4(write_data[20]), .I5(write_data[19]), .O(n570) );
  AND5_GATE U725 ( .I1(write_SCP), .I2(n444), .I3(n550), .I4(n571), .I5(n572), 
        .O(n564) );
  NOR4_GATE U726 ( .I1(write_data[11]), .I2(write_data[10]), .I3(write_adr[4]), 
        .I4(write_adr[3]), .O(n572) );
  INV_GATE U727 ( .I1(write_adr[2]), .O(n571) );
  NAND_GATE U728 ( .I1(n573), .I2(n574), .O(n563) );
  OR_GATE U729 ( .I1(n575), .I2(n2), .O(n574) );
  NAND_GATE U730 ( .I1(\scp_reg[12][0] ), .I2(n575), .O(n573) );
  AND_GATE U731 ( .I1(n576), .I2(n4), .O(n441) );
  NAND_GATE U732 ( .I1(n577), .I2(n578), .O(n794) );
  NAND_GATE U733 ( .I1(save_msk), .I2(n576), .O(n578) );
  NAND_GATE U734 ( .I1(\scp_reg[12][0] ), .I2(interrupt), .O(n577) );
  NAND_GATE U735 ( .I1(n579), .I2(n580), .O(n793) );
  NAND_GATE U736 ( .I1(n581), .I2(write_data[1]), .O(n580) );
  NAND_GATE U737 ( .I1(n582), .I2(\scp_reg[12][1] ), .O(n579) );
  NAND_GATE U738 ( .I1(n583), .I2(n584), .O(n792) );
  NAND_GATE U739 ( .I1(n581), .I2(write_data[2]), .O(n584) );
  NAND_GATE U740 ( .I1(n582), .I2(\scp_reg[12][2] ), .O(n583) );
  NAND_GATE U741 ( .I1(n585), .I2(n586), .O(n791) );
  NAND_GATE U742 ( .I1(n581), .I2(write_data[3]), .O(n586) );
  NAND_GATE U743 ( .I1(n582), .I2(\scp_reg[12][3] ), .O(n585) );
  NAND_GATE U744 ( .I1(n587), .I2(n588), .O(n790) );
  NAND_GATE U745 ( .I1(n581), .I2(write_data[4]), .O(n588) );
  NAND_GATE U746 ( .I1(n582), .I2(\scp_reg[12][4] ), .O(n587) );
  NAND_GATE U747 ( .I1(n589), .I2(n590), .O(n789) );
  NAND_GATE U748 ( .I1(n581), .I2(write_data[5]), .O(n590) );
  NAND_GATE U749 ( .I1(n582), .I2(\scp_reg[12][5] ), .O(n589) );
  NAND_GATE U750 ( .I1(n591), .I2(n592), .O(n788) );
  NAND_GATE U751 ( .I1(n581), .I2(write_data[6]), .O(n592) );
  NAND_GATE U752 ( .I1(n582), .I2(\scp_reg[12][6] ), .O(n591) );
  NAND_GATE U753 ( .I1(n593), .I2(n594), .O(n787) );
  NAND_GATE U754 ( .I1(n581), .I2(write_data[7]), .O(n594) );
  NAND_GATE U755 ( .I1(n582), .I2(\scp_reg[12][7] ), .O(n593) );
  NAND_GATE U756 ( .I1(n595), .I2(n596), .O(n786) );
  NAND_GATE U757 ( .I1(n581), .I2(write_data[8]), .O(n596) );
  NAND_GATE U758 ( .I1(n582), .I2(\scp_reg[12][8] ), .O(n595) );
  NAND_GATE U759 ( .I1(n597), .I2(n598), .O(n785) );
  NAND_GATE U760 ( .I1(n581), .I2(write_data[9]), .O(n598) );
  NAND_GATE U761 ( .I1(n582), .I2(\scp_reg[12][9] ), .O(n597) );
  NAND_GATE U762 ( .I1(n599), .I2(n600), .O(n784) );
  NAND_GATE U763 ( .I1(n581), .I2(write_data[10]), .O(n600) );
  NAND_GATE U764 ( .I1(n582), .I2(\scp_reg[12][10] ), .O(n599) );
  NAND_GATE U765 ( .I1(n601), .I2(n602), .O(n783) );
  NAND_GATE U766 ( .I1(n581), .I2(write_data[11]), .O(n602) );
  NAND_GATE U767 ( .I1(n582), .I2(\scp_reg[12][11] ), .O(n601) );
  NAND_GATE U768 ( .I1(n603), .I2(n604), .O(n782) );
  NAND_GATE U769 ( .I1(n581), .I2(write_data[12]), .O(n604) );
  NAND_GATE U770 ( .I1(n582), .I2(\scp_reg[12][12] ), .O(n603) );
  NAND_GATE U771 ( .I1(n605), .I2(n606), .O(n781) );
  NAND_GATE U772 ( .I1(n581), .I2(write_data[13]), .O(n606) );
  NAND_GATE U773 ( .I1(n582), .I2(\scp_reg[12][13] ), .O(n605) );
  NAND_GATE U774 ( .I1(n607), .I2(n608), .O(n780) );
  NAND_GATE U775 ( .I1(n581), .I2(write_data[14]), .O(n608) );
  NAND_GATE U776 ( .I1(n582), .I2(\scp_reg[12][14] ), .O(n607) );
  NAND_GATE U777 ( .I1(n609), .I2(n610), .O(n779) );
  NAND_GATE U778 ( .I1(n581), .I2(write_data[15]), .O(n610) );
  NAND_GATE U779 ( .I1(n582), .I2(\scp_reg[12][15] ), .O(n609) );
  NAND_GATE U780 ( .I1(n611), .I2(n612), .O(n778) );
  NAND_GATE U781 ( .I1(n581), .I2(write_data[16]), .O(n612) );
  NAND_GATE U782 ( .I1(n582), .I2(\scp_reg[12][16] ), .O(n611) );
  NAND_GATE U783 ( .I1(n613), .I2(n614), .O(n777) );
  NAND_GATE U784 ( .I1(n581), .I2(write_data[17]), .O(n614) );
  NAND_GATE U785 ( .I1(n582), .I2(\scp_reg[12][17] ), .O(n613) );
  NAND_GATE U786 ( .I1(n615), .I2(n616), .O(n776) );
  NAND_GATE U787 ( .I1(n581), .I2(write_data[18]), .O(n616) );
  NAND_GATE U788 ( .I1(n582), .I2(\scp_reg[12][18] ), .O(n615) );
  NAND_GATE U789 ( .I1(n617), .I2(n618), .O(n775) );
  NAND_GATE U790 ( .I1(n581), .I2(write_data[19]), .O(n618) );
  NAND_GATE U791 ( .I1(n582), .I2(\scp_reg[12][19] ), .O(n617) );
  NAND_GATE U792 ( .I1(n619), .I2(n620), .O(n774) );
  NAND_GATE U793 ( .I1(n581), .I2(write_data[20]), .O(n620) );
  NAND_GATE U794 ( .I1(n582), .I2(\scp_reg[12][20] ), .O(n619) );
  NAND_GATE U795 ( .I1(n621), .I2(n622), .O(n773) );
  NAND_GATE U796 ( .I1(n581), .I2(write_data[21]), .O(n622) );
  NAND_GATE U797 ( .I1(n582), .I2(\scp_reg[12][21] ), .O(n621) );
  NAND_GATE U798 ( .I1(n623), .I2(n624), .O(n772) );
  NAND_GATE U799 ( .I1(n581), .I2(write_data[22]), .O(n624) );
  NAND_GATE U800 ( .I1(n582), .I2(\scp_reg[12][22] ), .O(n623) );
  NAND_GATE U801 ( .I1(n625), .I2(n626), .O(n771) );
  NAND_GATE U802 ( .I1(n581), .I2(write_data[23]), .O(n626) );
  NAND_GATE U803 ( .I1(n582), .I2(\scp_reg[12][23] ), .O(n625) );
  NAND_GATE U804 ( .I1(n627), .I2(n628), .O(n770) );
  NAND_GATE U805 ( .I1(n581), .I2(write_data[24]), .O(n628) );
  NAND_GATE U806 ( .I1(n582), .I2(\scp_reg[12][24] ), .O(n627) );
  NAND_GATE U807 ( .I1(n629), .I2(n630), .O(n769) );
  NAND_GATE U808 ( .I1(n581), .I2(write_data[25]), .O(n630) );
  NAND_GATE U809 ( .I1(n582), .I2(\scp_reg[12][25] ), .O(n629) );
  NAND_GATE U810 ( .I1(n631), .I2(n632), .O(n768) );
  NAND_GATE U811 ( .I1(n581), .I2(write_data[26]), .O(n632) );
  NAND_GATE U812 ( .I1(n582), .I2(\scp_reg[12][26] ), .O(n631) );
  NAND_GATE U813 ( .I1(n633), .I2(n634), .O(n767) );
  NAND_GATE U814 ( .I1(n581), .I2(write_data[27]), .O(n634) );
  NAND_GATE U815 ( .I1(n582), .I2(\scp_reg[12][27] ), .O(n633) );
  NAND_GATE U816 ( .I1(n635), .I2(n636), .O(n766) );
  NAND_GATE U817 ( .I1(n581), .I2(write_data[28]), .O(n636) );
  NAND_GATE U818 ( .I1(n582), .I2(\scp_reg[12][28] ), .O(n635) );
  NAND_GATE U819 ( .I1(n637), .I2(n638), .O(n765) );
  NAND_GATE U820 ( .I1(n581), .I2(write_data[29]), .O(n638) );
  NAND_GATE U821 ( .I1(n582), .I2(\scp_reg[12][29] ), .O(n637) );
  NAND_GATE U822 ( .I1(n639), .I2(n640), .O(n764) );
  NAND_GATE U823 ( .I1(n581), .I2(write_data[30]), .O(n640) );
  NAND_GATE U824 ( .I1(n582), .I2(\scp_reg[12][30] ), .O(n639) );
  NAND_GATE U825 ( .I1(n641), .I2(n642), .O(n763) );
  NAND_GATE U826 ( .I1(n581), .I2(write_data[31]), .O(n642) );
  AND_GATE U827 ( .I1(n643), .I2(n4), .O(n581) );
  NAND_GATE U828 ( .I1(n582), .I2(\scp_reg[12][31] ), .O(n641) );
  AND_GATE U829 ( .I1(n575), .I2(n4), .O(n582) );
  INV_GATE U830 ( .I1(n643), .O(n575) );
  AND3_GATE U831 ( .I1(n444), .I2(n550), .I3(n549), .O(n643) );
  INV_GATE U832 ( .I1(write_adr[1]), .O(n550) );
  INV_GATE U833 ( .I1(write_adr[0]), .O(n444) );
  NAND_GATE U834 ( .I1(n644), .I2(n645), .O(n762) );
  NAND_GATE U835 ( .I1(n646), .I2(write_data[31]), .O(n645) );
  NAND_GATE U836 ( .I1(n647), .I2(\scp_reg[15][31] ), .O(n644) );
  NAND_GATE U837 ( .I1(n648), .I2(n649), .O(n761) );
  NAND_GATE U838 ( .I1(n646), .I2(write_data[30]), .O(n649) );
  NAND_GATE U839 ( .I1(n647), .I2(\scp_reg[15][30] ), .O(n648) );
  NAND_GATE U840 ( .I1(n650), .I2(n651), .O(n760) );
  NAND_GATE U841 ( .I1(n646), .I2(write_data[29]), .O(n651) );
  NAND_GATE U842 ( .I1(n647), .I2(\scp_reg[15][29] ), .O(n650) );
  NAND_GATE U843 ( .I1(n652), .I2(n653), .O(n759) );
  NAND_GATE U844 ( .I1(n646), .I2(write_data[28]), .O(n653) );
  NAND_GATE U845 ( .I1(n647), .I2(\scp_reg[15][28] ), .O(n652) );
  NAND_GATE U846 ( .I1(n654), .I2(n655), .O(n758) );
  NAND_GATE U847 ( .I1(n646), .I2(write_data[27]), .O(n655) );
  NAND_GATE U848 ( .I1(n647), .I2(\scp_reg[15][27] ), .O(n654) );
  NAND_GATE U849 ( .I1(n656), .I2(n657), .O(n757) );
  NAND_GATE U850 ( .I1(n646), .I2(write_data[26]), .O(n657) );
  NAND_GATE U851 ( .I1(n647), .I2(\scp_reg[15][26] ), .O(n656) );
  NAND_GATE U852 ( .I1(n658), .I2(n659), .O(n756) );
  NAND_GATE U853 ( .I1(n646), .I2(write_data[25]), .O(n659) );
  NAND_GATE U854 ( .I1(n647), .I2(\scp_reg[15][25] ), .O(n658) );
  NAND_GATE U855 ( .I1(n660), .I2(n661), .O(n755) );
  NAND_GATE U856 ( .I1(n646), .I2(write_data[24]), .O(n661) );
  NAND_GATE U857 ( .I1(n647), .I2(\scp_reg[15][24] ), .O(n660) );
  NAND_GATE U858 ( .I1(n662), .I2(n663), .O(n754) );
  NAND_GATE U859 ( .I1(n646), .I2(write_data[23]), .O(n663) );
  NAND_GATE U860 ( .I1(n647), .I2(\scp_reg[15][23] ), .O(n662) );
  NAND_GATE U861 ( .I1(n664), .I2(n665), .O(n753) );
  NAND_GATE U862 ( .I1(n646), .I2(write_data[22]), .O(n665) );
  NAND_GATE U863 ( .I1(n647), .I2(\scp_reg[15][22] ), .O(n664) );
  NAND_GATE U864 ( .I1(n666), .I2(n667), .O(n752) );
  NAND_GATE U865 ( .I1(n646), .I2(write_data[21]), .O(n667) );
  NAND_GATE U866 ( .I1(n647), .I2(\scp_reg[15][21] ), .O(n666) );
  NAND_GATE U867 ( .I1(n668), .I2(n669), .O(n751) );
  NAND_GATE U868 ( .I1(n646), .I2(write_data[20]), .O(n669) );
  NAND_GATE U869 ( .I1(n647), .I2(\scp_reg[15][20] ), .O(n668) );
  NAND_GATE U870 ( .I1(n670), .I2(n671), .O(n750) );
  NAND_GATE U871 ( .I1(n646), .I2(write_data[19]), .O(n671) );
  NAND_GATE U872 ( .I1(n647), .I2(\scp_reg[15][19] ), .O(n670) );
  NAND_GATE U873 ( .I1(n672), .I2(n673), .O(n749) );
  NAND_GATE U874 ( .I1(n646), .I2(write_data[18]), .O(n673) );
  NAND_GATE U875 ( .I1(n647), .I2(\scp_reg[15][18] ), .O(n672) );
  NAND_GATE U876 ( .I1(n674), .I2(n675), .O(n748) );
  NAND_GATE U877 ( .I1(n646), .I2(write_data[17]), .O(n675) );
  NAND_GATE U878 ( .I1(n647), .I2(\scp_reg[15][17] ), .O(n674) );
  NAND_GATE U879 ( .I1(n676), .I2(n677), .O(n747) );
  NAND_GATE U880 ( .I1(n646), .I2(write_data[16]), .O(n677) );
  NAND_GATE U881 ( .I1(n647), .I2(\scp_reg[15][16] ), .O(n676) );
  NAND_GATE U882 ( .I1(n678), .I2(n679), .O(n746) );
  NAND_GATE U883 ( .I1(n646), .I2(write_data[15]), .O(n679) );
  NAND_GATE U884 ( .I1(n647), .I2(\scp_reg[15][15] ), .O(n678) );
  NAND_GATE U885 ( .I1(n680), .I2(n681), .O(n745) );
  NAND_GATE U886 ( .I1(n646), .I2(write_data[14]), .O(n681) );
  NAND_GATE U887 ( .I1(n647), .I2(\scp_reg[15][14] ), .O(n680) );
  NAND_GATE U888 ( .I1(n682), .I2(n683), .O(n744) );
  NAND_GATE U889 ( .I1(n646), .I2(write_data[13]), .O(n683) );
  NAND_GATE U890 ( .I1(n647), .I2(\scp_reg[15][13] ), .O(n682) );
  NAND_GATE U891 ( .I1(n684), .I2(n685), .O(n743) );
  NAND_GATE U892 ( .I1(n646), .I2(write_data[12]), .O(n685) );
  NAND_GATE U893 ( .I1(n647), .I2(\scp_reg[15][12] ), .O(n684) );
  NAND_GATE U894 ( .I1(n686), .I2(n687), .O(n742) );
  NAND_GATE U895 ( .I1(n646), .I2(write_data[11]), .O(n687) );
  NAND_GATE U896 ( .I1(n647), .I2(\scp_reg[15][11] ), .O(n686) );
  NAND_GATE U897 ( .I1(n688), .I2(n689), .O(n741) );
  NAND_GATE U898 ( .I1(n646), .I2(write_data[10]), .O(n689) );
  NAND_GATE U899 ( .I1(n647), .I2(\scp_reg[15][10] ), .O(n688) );
  NAND_GATE U900 ( .I1(n690), .I2(n691), .O(n740) );
  NAND_GATE U901 ( .I1(n646), .I2(write_data[9]), .O(n691) );
  NAND_GATE U902 ( .I1(n647), .I2(\scp_reg[15][9] ), .O(n690) );
  NAND_GATE U903 ( .I1(n692), .I2(n693), .O(n739) );
  NAND_GATE U904 ( .I1(n646), .I2(write_data[8]), .O(n693) );
  NAND_GATE U905 ( .I1(n647), .I2(\scp_reg[15][8] ), .O(n692) );
  NAND_GATE U906 ( .I1(n694), .I2(n695), .O(n738) );
  NAND_GATE U907 ( .I1(n646), .I2(write_data[7]), .O(n695) );
  NAND_GATE U908 ( .I1(n647), .I2(\scp_reg[15][7] ), .O(n694) );
  NAND_GATE U909 ( .I1(n696), .I2(n697), .O(n737) );
  NAND_GATE U910 ( .I1(n646), .I2(write_data[6]), .O(n697) );
  NAND_GATE U911 ( .I1(n647), .I2(\scp_reg[15][6] ), .O(n696) );
  NAND_GATE U912 ( .I1(n698), .I2(n699), .O(n736) );
  NAND_GATE U913 ( .I1(n646), .I2(write_data[5]), .O(n699) );
  NAND_GATE U914 ( .I1(n647), .I2(\scp_reg[15][5] ), .O(n698) );
  NAND_GATE U915 ( .I1(n700), .I2(n701), .O(n735) );
  NAND_GATE U916 ( .I1(n646), .I2(write_data[4]), .O(n701) );
  NAND_GATE U917 ( .I1(n647), .I2(\scp_reg[15][4] ), .O(n700) );
  NAND_GATE U918 ( .I1(n702), .I2(n703), .O(n734) );
  NAND_GATE U919 ( .I1(n646), .I2(write_data[3]), .O(n703) );
  NAND_GATE U920 ( .I1(n647), .I2(\scp_reg[15][3] ), .O(n702) );
  NAND_GATE U921 ( .I1(n704), .I2(n705), .O(n733) );
  NAND_GATE U922 ( .I1(n646), .I2(write_data[2]), .O(n705) );
  NAND_GATE U923 ( .I1(n647), .I2(\scp_reg[15][2] ), .O(n704) );
  NAND_GATE U924 ( .I1(n706), .I2(n707), .O(n732) );
  NAND_GATE U925 ( .I1(n646), .I2(write_data[1]), .O(n707) );
  NAND_GATE U926 ( .I1(n647), .I2(\scp_reg[15][1] ), .O(n706) );
  NAND_GATE U927 ( .I1(n708), .I2(n709), .O(n731) );
  NAND_GATE U928 ( .I1(n646), .I2(write_data[0]), .O(n709) );
  AND3_GATE U929 ( .I1(n443), .I2(n4), .I3(write_adr[0]), .O(n646) );
  NAND_GATE U930 ( .I1(n647), .I2(\scp_reg[15][0] ), .O(n708) );
  AND_GATE U931 ( .I1(n710), .I2(n4), .O(n647) );
  NAND_GATE U932 ( .I1(write_adr[0]), .I2(n443), .O(n710) );
  AND_GATE U933 ( .I1(write_adr[1]), .I2(n549), .O(n443) );
  AND4_GATE U934 ( .I1(write_adr[3]), .I2(write_adr[2]), .I3(write_SCP), .I4(
        n711), .O(n549) );
  INV_GATE U935 ( .I1(write_adr[4]), .O(n711) );
  INV_GATE U936 ( .I1(n576), .O(interrupt) );
  AND_GATE U937 ( .I1(n544), .I2(n548), .O(n576) );
  NAND3_GATE U938 ( .I1(MEM_it_ok), .I2(\scp_reg[12][0] ), .I3(it_mat), .O(
        n548) );
  AND4_GATE U939 ( .I1(n712), .I2(n713), .I3(n714), .I4(n715), .O(n544) );
  NOR5_GATE U940 ( .I1(MEM_exc_cause[31]), .I2(MEM_exc_cause[3]), .I3(
        MEM_exc_cause[4]), .I4(MEM_exc_cause[5]), .I5(n716), .O(n715) );
  OR4_GATE U941 ( .I1(MEM_exc_cause[9]), .I2(MEM_exc_cause[8]), .I3(
        MEM_exc_cause[7]), .I4(MEM_exc_cause[6]), .O(n716) );
  NOR5_GATE U942 ( .I1(MEM_exc_cause[24]), .I2(MEM_exc_cause[25]), .I3(
        MEM_exc_cause[26]), .I4(MEM_exc_cause[27]), .I5(n717), .O(n714) );
  OR4_GATE U943 ( .I1(MEM_exc_cause[30]), .I2(MEM_exc_cause[2]), .I3(
        MEM_exc_cause[29]), .I4(MEM_exc_cause[28]), .O(n717) );
  NOR5_GATE U944 ( .I1(MEM_exc_cause[17]), .I2(MEM_exc_cause[18]), .I3(
        MEM_exc_cause[19]), .I4(MEM_exc_cause[1]), .I5(n718), .O(n713) );
  OR4_GATE U945 ( .I1(MEM_exc_cause[23]), .I2(MEM_exc_cause[22]), .I3(
        MEM_exc_cause[21]), .I4(MEM_exc_cause[20]), .O(n718) );
  NOR5_GATE U946 ( .I1(MEM_exc_cause[0]), .I2(MEM_exc_cause[10]), .I3(
        MEM_exc_cause[11]), .I4(MEM_exc_cause[12]), .I5(n719), .O(n712) );
  OR4_GATE U947 ( .I1(MEM_exc_cause[16]), .I2(MEM_exc_cause[15]), .I3(
        MEM_exc_cause[14]), .I4(MEM_exc_cause[13]), .O(n719) );
endmodule


module banc ( clock, reset, reg_src1, reg_src2, reg_dest, donnee, cmd_ecr, 
        data_src1, data_src2 );
  input [4:0] reg_src1;
  input [4:0] reg_src2;
  input [4:0] reg_dest;
  input [31:0] donnee;
  output [31:0] data_src1;
  output [31:0] data_src2;
  input clock, reset, cmd_ecr;
  wire   \registres[1][31] , \registres[1][30] , \registres[1][29] ,
         \registres[1][28] , \registres[1][27] , \registres[1][26] ,
         \registres[1][25] , \registres[1][24] , \registres[1][23] ,
         \registres[1][22] , \registres[1][21] , \registres[1][20] ,
         \registres[1][19] , \registres[1][18] , \registres[1][17] ,
         \registres[1][16] , \registres[1][15] , \registres[1][14] ,
         \registres[1][13] , \registres[1][12] , \registres[1][11] ,
         \registres[1][10] , \registres[1][9] , \registres[1][8] ,
         \registres[1][7] , \registres[1][6] , \registres[1][5] ,
         \registres[1][4] , \registres[1][3] , \registres[1][2] ,
         \registres[1][1] , \registres[1][0] , \registres[2][31] ,
         \registres[2][30] , \registres[2][29] , \registres[2][28] ,
         \registres[2][27] , \registres[2][26] , \registres[2][25] ,
         \registres[2][24] , \registres[2][23] , \registres[2][22] ,
         \registres[2][21] , \registres[2][20] , \registres[2][19] ,
         \registres[2][18] , \registres[2][17] , \registres[2][16] ,
         \registres[2][15] , \registres[2][14] , \registres[2][13] ,
         \registres[2][12] , \registres[2][11] , \registres[2][10] ,
         \registres[2][9] , \registres[2][8] , \registres[2][7] ,
         \registres[2][6] , \registres[2][5] , \registres[2][4] ,
         \registres[2][3] , \registres[2][2] , \registres[2][1] ,
         \registres[2][0] , \registres[3][31] , \registres[3][30] ,
         \registres[3][29] , \registres[3][28] , \registres[3][27] ,
         \registres[3][26] , \registres[3][25] , \registres[3][24] ,
         \registres[3][23] , \registres[3][22] , \registres[3][21] ,
         \registres[3][20] , \registres[3][19] , \registres[3][18] ,
         \registres[3][17] , \registres[3][16] , \registres[3][15] ,
         \registres[3][14] , \registres[3][13] , \registres[3][12] ,
         \registres[3][11] , \registres[3][10] , \registres[3][9] ,
         \registres[3][8] , \registres[3][7] , \registres[3][6] ,
         \registres[3][5] , \registres[3][4] , \registres[3][3] ,
         \registres[3][2] , \registres[3][1] , \registres[3][0] ,
         \registres[4][31] , \registres[4][30] , \registres[4][29] ,
         \registres[4][28] , \registres[4][27] , \registres[4][26] ,
         \registres[4][25] , \registres[4][24] , \registres[4][23] ,
         \registres[4][22] , \registres[4][21] , \registres[4][20] ,
         \registres[4][19] , \registres[4][18] , \registres[4][17] ,
         \registres[4][16] , \registres[4][15] , \registres[4][14] ,
         \registres[4][13] , \registres[4][12] , \registres[4][11] ,
         \registres[4][10] , \registres[4][9] , \registres[4][8] ,
         \registres[4][7] , \registres[4][6] , \registres[4][5] ,
         \registres[4][4] , \registres[4][3] , \registres[4][2] ,
         \registres[4][1] , \registres[4][0] , \registres[5][31] ,
         \registres[5][30] , \registres[5][29] , \registres[5][28] ,
         \registres[5][27] , \registres[5][26] , \registres[5][25] ,
         \registres[5][24] , \registres[5][23] , \registres[5][22] ,
         \registres[5][21] , \registres[5][20] , \registres[5][19] ,
         \registres[5][18] , \registres[5][17] , \registres[5][16] ,
         \registres[5][15] , \registres[5][14] , \registres[5][13] ,
         \registres[5][12] , \registres[5][11] , \registres[5][10] ,
         \registres[5][9] , \registres[5][8] , \registres[5][7] ,
         \registres[5][6] , \registres[5][5] , \registres[5][4] ,
         \registres[5][3] , \registres[5][2] , \registres[5][1] ,
         \registres[5][0] , \registres[6][31] , \registres[6][30] ,
         \registres[6][29] , \registres[6][28] , \registres[6][27] ,
         \registres[6][26] , \registres[6][25] , \registres[6][24] ,
         \registres[6][23] , \registres[6][22] , \registres[6][21] ,
         \registres[6][20] , \registres[6][19] , \registres[6][18] ,
         \registres[6][17] , \registres[6][16] , \registres[6][15] ,
         \registres[6][14] , \registres[6][13] , \registres[6][12] ,
         \registres[6][11] , \registres[6][10] , \registres[6][9] ,
         \registres[6][8] , \registres[6][7] , \registres[6][6] ,
         \registres[6][5] , \registres[6][4] , \registres[6][3] ,
         \registres[6][2] , \registres[6][1] , \registres[6][0] ,
         \registres[7][31] , \registres[7][30] , \registres[7][29] ,
         \registres[7][28] , \registres[7][27] , \registres[7][26] ,
         \registres[7][25] , \registres[7][24] , \registres[7][23] ,
         \registres[7][22] , \registres[7][21] , \registres[7][20] ,
         \registres[7][19] , \registres[7][18] , \registres[7][17] ,
         \registres[7][16] , \registres[7][15] , \registres[7][14] ,
         \registres[7][13] , \registres[7][12] , \registres[7][11] ,
         \registres[7][10] , \registres[7][9] , \registres[7][8] ,
         \registres[7][7] , \registres[7][6] , \registres[7][5] ,
         \registres[7][4] , \registres[7][3] , \registres[7][2] ,
         \registres[7][1] , \registres[7][0] , \registres[8][31] ,
         \registres[8][30] , \registres[8][29] , \registres[8][28] ,
         \registres[8][27] , \registres[8][26] , \registres[8][25] ,
         \registres[8][24] , \registres[8][23] , \registres[8][22] ,
         \registres[8][21] , \registres[8][20] , \registres[8][19] ,
         \registres[8][18] , \registres[8][17] , \registres[8][16] ,
         \registres[8][15] , \registres[8][14] , \registres[8][13] ,
         \registres[8][12] , \registres[8][11] , \registres[8][10] ,
         \registres[8][9] , \registres[8][8] , \registres[8][7] ,
         \registres[8][6] , \registres[8][5] , \registres[8][4] ,
         \registres[8][3] , \registres[8][2] , \registres[8][1] ,
         \registres[8][0] , \registres[9][31] , \registres[9][30] ,
         \registres[9][29] , \registres[9][28] , \registres[9][27] ,
         \registres[9][26] , \registres[9][25] , \registres[9][24] ,
         \registres[9][23] , \registres[9][22] , \registres[9][21] ,
         \registres[9][20] , \registres[9][19] , \registres[9][18] ,
         \registres[9][17] , \registres[9][16] , \registres[9][15] ,
         \registres[9][14] , \registres[9][13] , \registres[9][12] ,
         \registres[9][11] , \registres[9][10] , \registres[9][9] ,
         \registres[9][8] , \registres[9][7] , \registres[9][6] ,
         \registres[9][5] , \registres[9][4] , \registres[9][3] ,
         \registres[9][2] , \registres[9][1] , \registres[9][0] ,
         \registres[10][31] , \registres[10][30] , \registres[10][29] ,
         \registres[10][28] , \registres[10][27] , \registres[10][26] ,
         \registres[10][25] , \registres[10][24] , \registres[10][23] ,
         \registres[10][22] , \registres[10][21] , \registres[10][20] ,
         \registres[10][19] , \registres[10][18] , \registres[10][17] ,
         \registres[10][16] , \registres[10][15] , \registres[10][14] ,
         \registres[10][13] , \registres[10][12] , \registres[10][11] ,
         \registres[10][10] , \registres[10][9] , \registres[10][8] ,
         \registres[10][7] , \registres[10][6] , \registres[10][5] ,
         \registres[10][4] , \registres[10][3] , \registres[10][2] ,
         \registres[10][1] , \registres[10][0] , \registres[11][31] ,
         \registres[11][30] , \registres[11][29] , \registres[11][28] ,
         \registres[11][27] , \registres[11][26] , \registres[11][25] ,
         \registres[11][24] , \registres[11][23] , \registres[11][22] ,
         \registres[11][21] , \registres[11][20] , \registres[11][19] ,
         \registres[11][18] , \registres[11][17] , \registres[11][16] ,
         \registres[11][15] , \registres[11][14] , \registres[11][13] ,
         \registres[11][12] , \registres[11][11] , \registres[11][10] ,
         \registres[11][9] , \registres[11][8] , \registres[11][7] ,
         \registres[11][6] , \registres[11][5] , \registres[11][4] ,
         \registres[11][3] , \registres[11][2] , \registres[11][1] ,
         \registres[11][0] , \registres[12][31] , \registres[12][30] ,
         \registres[12][29] , \registres[12][28] , \registres[12][27] ,
         \registres[12][26] , \registres[12][25] , \registres[12][24] ,
         \registres[12][23] , \registres[12][22] , \registres[12][21] ,
         \registres[12][20] , \registres[12][19] , \registres[12][18] ,
         \registres[12][17] , \registres[12][16] , \registres[12][15] ,
         \registres[12][14] , \registres[12][13] , \registres[12][12] ,
         \registres[12][11] , \registres[12][10] , \registres[12][9] ,
         \registres[12][8] , \registres[12][7] , \registres[12][6] ,
         \registres[12][5] , \registres[12][4] , \registres[12][3] ,
         \registres[12][2] , \registres[12][1] , \registres[12][0] ,
         \registres[13][31] , \registres[13][30] , \registres[13][29] ,
         \registres[13][28] , \registres[13][27] , \registres[13][26] ,
         \registres[13][25] , \registres[13][24] , \registres[13][23] ,
         \registres[13][22] , \registres[13][21] , \registres[13][20] ,
         \registres[13][19] , \registres[13][18] , \registres[13][17] ,
         \registres[13][16] , \registres[13][15] , \registres[13][14] ,
         \registres[13][13] , \registres[13][12] , \registres[13][11] ,
         \registres[13][10] , \registres[13][9] , \registres[13][8] ,
         \registres[13][7] , \registres[13][6] , \registres[13][5] ,
         \registres[13][4] , \registres[13][3] , \registres[13][2] ,
         \registres[13][1] , \registres[13][0] , \registres[14][31] ,
         \registres[14][30] , \registres[14][29] , \registres[14][28] ,
         \registres[14][27] , \registres[14][26] , \registres[14][25] ,
         \registres[14][24] , \registres[14][23] , \registres[14][22] ,
         \registres[14][21] , \registres[14][20] , \registres[14][19] ,
         \registres[14][18] , \registres[14][17] , \registres[14][16] ,
         \registres[14][15] , \registres[14][14] , \registres[14][13] ,
         \registres[14][12] , \registres[14][11] , \registres[14][10] ,
         \registres[14][9] , \registres[14][8] , \registres[14][7] ,
         \registres[14][6] , \registres[14][5] , \registres[14][4] ,
         \registres[14][3] , \registres[14][2] , \registres[14][1] ,
         \registres[14][0] , \registres[15][31] , \registres[15][30] ,
         \registres[15][29] , \registres[15][28] , \registres[15][27] ,
         \registres[15][26] , \registres[15][25] , \registres[15][24] ,
         \registres[15][23] , \registres[15][22] , \registres[15][21] ,
         \registres[15][20] , \registres[15][19] , \registres[15][18] ,
         \registres[15][17] , \registres[15][16] , \registres[15][15] ,
         \registres[15][14] , \registres[15][13] , \registres[15][12] ,
         \registres[15][11] , \registres[15][10] , \registres[15][9] ,
         \registres[15][8] , \registres[15][7] , \registres[15][6] ,
         \registres[15][5] , \registres[15][4] , \registres[15][3] ,
         \registres[15][2] , \registres[15][1] , \registres[15][0] ,
         \registres[16][31] , \registres[16][30] , \registres[16][29] ,
         \registres[16][28] , \registres[16][27] , \registres[16][26] ,
         \registres[16][25] , \registres[16][24] , \registres[16][23] ,
         \registres[16][22] , \registres[16][21] , \registres[16][20] ,
         \registres[16][19] , \registres[16][18] , \registres[16][17] ,
         \registres[16][16] , \registres[16][15] , \registres[16][14] ,
         \registres[16][13] , \registres[16][12] , \registres[16][11] ,
         \registres[16][10] , \registres[16][9] , \registres[16][8] ,
         \registres[16][7] , \registres[16][6] , \registres[16][5] ,
         \registres[16][4] , \registres[16][3] , \registres[16][2] ,
         \registres[16][1] , \registres[16][0] , \registres[17][31] ,
         \registres[17][30] , \registres[17][29] , \registres[17][28] ,
         \registres[17][27] , \registres[17][26] , \registres[17][25] ,
         \registres[17][24] , \registres[17][23] , \registres[17][22] ,
         \registres[17][21] , \registres[17][20] , \registres[17][19] ,
         \registres[17][18] , \registres[17][17] , \registres[17][16] ,
         \registres[17][15] , \registres[17][14] , \registres[17][13] ,
         \registres[17][12] , \registres[17][11] , \registres[17][10] ,
         \registres[17][9] , \registres[17][8] , \registres[17][7] ,
         \registres[17][6] , \registres[17][5] , \registres[17][4] ,
         \registres[17][3] , \registres[17][2] , \registres[17][1] ,
         \registres[17][0] , \registres[18][31] , \registres[18][30] ,
         \registres[18][29] , \registres[18][28] , \registres[18][27] ,
         \registres[18][26] , \registres[18][25] , \registres[18][24] ,
         \registres[18][23] , \registres[18][22] , \registres[18][21] ,
         \registres[18][20] , \registres[18][19] , \registres[18][18] ,
         \registres[18][17] , \registres[18][16] , \registres[18][15] ,
         \registres[18][14] , \registres[18][13] , \registres[18][12] ,
         \registres[18][11] , \registres[18][10] , \registres[18][9] ,
         \registres[18][8] , \registres[18][7] , \registres[18][6] ,
         \registres[18][5] , \registres[18][4] , \registres[18][3] ,
         \registres[18][2] , \registres[18][1] , \registres[18][0] ,
         \registres[19][31] , \registres[19][30] , \registres[19][29] ,
         \registres[19][28] , \registres[19][27] , \registres[19][26] ,
         \registres[19][25] , \registres[19][24] , \registres[19][23] ,
         \registres[19][22] , \registres[19][21] , \registres[19][20] ,
         \registres[19][19] , \registres[19][18] , \registres[19][17] ,
         \registres[19][16] , \registres[19][15] , \registres[19][14] ,
         \registres[19][13] , \registres[19][12] , \registres[19][11] ,
         \registres[19][10] , \registres[19][9] , \registres[19][8] ,
         \registres[19][7] , \registres[19][6] , \registres[19][5] ,
         \registres[19][4] , \registres[19][3] , \registres[19][2] ,
         \registres[19][1] , \registres[19][0] , \registres[20][31] ,
         \registres[20][30] , \registres[20][29] , \registres[20][28] ,
         \registres[20][27] , \registres[20][26] , \registres[20][25] ,
         \registres[20][24] , \registres[20][23] , \registres[20][22] ,
         \registres[20][21] , \registres[20][20] , \registres[20][19] ,
         \registres[20][18] , \registres[20][17] , \registres[20][16] ,
         \registres[20][15] , \registres[20][14] , \registres[20][13] ,
         \registres[20][12] , \registres[20][11] , \registres[20][10] ,
         \registres[20][9] , \registres[20][8] , \registres[20][7] ,
         \registres[20][6] , \registres[20][5] , \registres[20][4] ,
         \registres[20][3] , \registres[20][2] , \registres[20][1] ,
         \registres[20][0] , \registres[21][31] , \registres[21][30] ,
         \registres[21][29] , \registres[21][28] , \registres[21][27] ,
         \registres[21][26] , \registres[21][25] , \registres[21][24] ,
         \registres[21][23] , \registres[21][22] , \registres[21][21] ,
         \registres[21][20] , \registres[21][19] , \registres[21][18] ,
         \registres[21][17] , \registres[21][16] , \registres[21][15] ,
         \registres[21][14] , \registres[21][13] , \registres[21][12] ,
         \registres[21][11] , \registres[21][10] , \registres[21][9] ,
         \registres[21][8] , \registres[21][7] , \registres[21][6] ,
         \registres[21][5] , \registres[21][4] , \registres[21][3] ,
         \registres[21][2] , \registres[21][1] , \registres[21][0] ,
         \registres[22][31] , \registres[22][30] , \registres[22][29] ,
         \registres[22][28] , \registres[22][27] , \registres[22][26] ,
         \registres[22][25] , \registres[22][24] , \registres[22][23] ,
         \registres[22][22] , \registres[22][21] , \registres[22][20] ,
         \registres[22][19] , \registres[22][18] , \registres[22][17] ,
         \registres[22][16] , \registres[22][15] , \registres[22][14] ,
         \registres[22][13] , \registres[22][12] , \registres[22][11] ,
         \registres[22][10] , \registres[22][9] , \registres[22][8] ,
         \registres[22][7] , \registres[22][6] , \registres[22][5] ,
         \registres[22][4] , \registres[22][3] , \registres[22][2] ,
         \registres[22][1] , \registres[22][0] , \registres[23][31] ,
         \registres[23][30] , \registres[23][29] , \registres[23][28] ,
         \registres[23][27] , \registres[23][26] , \registres[23][25] ,
         \registres[23][24] , \registres[23][23] , \registres[23][22] ,
         \registres[23][21] , \registres[23][20] , \registres[23][19] ,
         \registres[23][18] , \registres[23][17] , \registres[23][16] ,
         \registres[23][15] , \registres[23][14] , \registres[23][13] ,
         \registres[23][12] , \registres[23][11] , \registres[23][10] ,
         \registres[23][9] , \registres[23][8] , \registres[23][7] ,
         \registres[23][6] , \registres[23][5] , \registres[23][4] ,
         \registres[23][3] , \registres[23][2] , \registres[23][1] ,
         \registres[23][0] , \registres[24][31] , \registres[24][30] ,
         \registres[24][29] , \registres[24][28] , \registres[24][27] ,
         \registres[24][26] , \registres[24][25] , \registres[24][24] ,
         \registres[24][23] , \registres[24][22] , \registres[24][21] ,
         \registres[24][20] , \registres[24][19] , \registres[24][18] ,
         \registres[24][17] , \registres[24][16] , \registres[24][15] ,
         \registres[24][14] , \registres[24][13] , \registres[24][12] ,
         \registres[24][11] , \registres[24][10] , \registres[24][9] ,
         \registres[24][8] , \registres[24][7] , \registres[24][6] ,
         \registres[24][5] , \registres[24][4] , \registres[24][3] ,
         \registres[24][2] , \registres[24][1] , \registres[24][0] ,
         \registres[25][31] , \registres[25][30] , \registres[25][29] ,
         \registres[25][28] , \registres[25][27] , \registres[25][26] ,
         \registres[25][25] , \registres[25][24] , \registres[25][23] ,
         \registres[25][22] , \registres[25][21] , \registres[25][20] ,
         \registres[25][19] , \registres[25][18] , \registres[25][17] ,
         \registres[25][16] , \registres[25][15] , \registres[25][14] ,
         \registres[25][13] , \registres[25][12] , \registres[25][11] ,
         \registres[25][10] , \registres[25][9] , \registres[25][8] ,
         \registres[25][7] , \registres[25][6] , \registres[25][5] ,
         \registres[25][4] , \registres[25][3] , \registres[25][2] ,
         \registres[25][1] , \registres[25][0] , \registres[26][31] ,
         \registres[26][30] , \registres[26][29] , \registres[26][28] ,
         \registres[26][27] , \registres[26][26] , \registres[26][25] ,
         \registres[26][24] , \registres[26][23] , \registres[26][22] ,
         \registres[26][21] , \registres[26][20] , \registres[26][19] ,
         \registres[26][18] , \registres[26][17] , \registres[26][16] ,
         \registres[26][15] , \registres[26][14] , \registres[26][13] ,
         \registres[26][12] , \registres[26][11] , \registres[26][10] ,
         \registres[26][9] , \registres[26][8] , \registres[26][7] ,
         \registres[26][6] , \registres[26][5] , \registres[26][4] ,
         \registres[26][3] , \registres[26][2] , \registres[26][1] ,
         \registres[26][0] , \registres[27][31] , \registres[27][30] ,
         \registres[27][29] , \registres[27][28] , \registres[27][27] ,
         \registres[27][26] , \registres[27][25] , \registres[27][24] ,
         \registres[27][23] , \registres[27][22] , \registres[27][21] ,
         \registres[27][20] , \registres[27][19] , \registres[27][18] ,
         \registres[27][17] , \registres[27][16] , \registres[27][15] ,
         \registres[27][14] , \registres[27][13] , \registres[27][12] ,
         \registres[27][11] , \registres[27][10] , \registres[27][9] ,
         \registres[27][8] , \registres[27][7] , \registres[27][6] ,
         \registres[27][5] , \registres[27][4] , \registres[27][3] ,
         \registres[27][2] , \registres[27][1] , \registres[27][0] ,
         \registres[28][31] , \registres[28][30] , \registres[28][29] ,
         \registres[28][28] , \registres[28][27] , \registres[28][26] ,
         \registres[28][25] , \registres[28][24] , \registres[28][23] ,
         \registres[28][22] , \registres[28][21] , \registres[28][20] ,
         \registres[28][19] , \registres[28][18] , \registres[28][17] ,
         \registres[28][16] , \registres[28][15] , \registres[28][14] ,
         \registres[28][13] , \registres[28][12] , \registres[28][11] ,
         \registres[28][10] , \registres[28][9] , \registres[28][8] ,
         \registres[28][7] , \registres[28][6] , \registres[28][5] ,
         \registres[28][4] , \registres[28][3] , \registres[28][2] ,
         \registres[28][1] , \registres[28][0] , \registres[29][31] ,
         \registres[29][30] , \registres[29][29] , \registres[29][28] ,
         \registres[29][27] , \registres[29][26] , \registres[29][25] ,
         \registres[29][24] , \registres[29][23] , \registres[29][22] ,
         \registres[29][21] , \registres[29][20] , \registres[29][19] ,
         \registres[29][18] , \registres[29][17] , \registres[29][16] ,
         \registres[29][15] , \registres[29][14] , \registres[29][13] ,
         \registres[29][12] , \registres[29][11] , \registres[29][10] ,
         \registres[29][9] , \registres[29][8] , \registres[29][7] ,
         \registres[29][6] , \registres[29][5] , \registres[29][4] ,
         \registres[29][3] , \registres[29][2] , \registres[29][1] ,
         \registres[29][0] , \registres[30][31] , \registres[30][30] ,
         \registres[30][29] , \registres[30][28] , \registres[30][27] ,
         \registres[30][26] , \registres[30][25] , \registres[30][24] ,
         \registres[30][23] , \registres[30][22] , \registres[30][21] ,
         \registres[30][20] , \registres[30][19] , \registres[30][18] ,
         \registres[30][17] , \registres[30][16] , \registres[30][15] ,
         \registres[30][14] , \registres[30][13] , \registres[30][12] ,
         \registres[30][11] , \registres[30][10] , \registres[30][9] ,
         \registres[30][8] , \registres[30][7] , \registres[30][6] ,
         \registres[30][5] , \registres[30][4] , \registres[30][3] ,
         \registres[30][2] , \registres[30][1] , \registres[30][0] ,
         \registres[31][31] , \registres[31][30] , \registres[31][29] ,
         \registres[31][28] , \registres[31][27] , \registres[31][26] ,
         \registres[31][25] , \registres[31][24] , \registres[31][23] ,
         \registres[31][22] , \registres[31][21] , \registres[31][20] ,
         \registres[31][19] , \registres[31][18] , \registres[31][17] ,
         \registres[31][16] , \registres[31][15] , \registres[31][14] ,
         \registres[31][13] , \registres[31][12] , \registres[31][11] ,
         \registres[31][10] , \registres[31][9] , \registres[31][8] ,
         \registres[31][7] , \registres[31][6] , \registres[31][5] ,
         \registres[31][4] , \registres[31][3] , \registres[31][2] ,
         \registres[31][1] , \registres[31][0] , n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14;

  FLIP_FLOP_D \registres_reg[1][31]  ( .D(n5750), .CK(clock), .Q(
        \registres[1][31] ) );
  FLIP_FLOP_D \registres_reg[1][30]  ( .D(n5749), .CK(clock), .Q(
        \registres[1][30] ) );
  FLIP_FLOP_D \registres_reg[1][29]  ( .D(n5748), .CK(clock), .Q(
        \registres[1][29] ) );
  FLIP_FLOP_D \registres_reg[1][28]  ( .D(n5747), .CK(clock), .Q(
        \registres[1][28] ) );
  FLIP_FLOP_D \registres_reg[1][27]  ( .D(n5746), .CK(clock), .Q(
        \registres[1][27] ) );
  FLIP_FLOP_D \registres_reg[1][26]  ( .D(n5745), .CK(clock), .Q(
        \registres[1][26] ) );
  FLIP_FLOP_D \registres_reg[1][25]  ( .D(n5744), .CK(clock), .Q(
        \registres[1][25] ) );
  FLIP_FLOP_D \registres_reg[1][24]  ( .D(n5743), .CK(clock), .Q(
        \registres[1][24] ) );
  FLIP_FLOP_D \registres_reg[1][23]  ( .D(n5742), .CK(clock), .Q(
        \registres[1][23] ) );
  FLIP_FLOP_D \registres_reg[1][22]  ( .D(n5741), .CK(clock), .Q(
        \registres[1][22] ) );
  FLIP_FLOP_D \registres_reg[1][21]  ( .D(n5740), .CK(clock), .Q(
        \registres[1][21] ) );
  FLIP_FLOP_D \registres_reg[1][20]  ( .D(n5739), .CK(clock), .Q(
        \registres[1][20] ) );
  FLIP_FLOP_D \registres_reg[1][19]  ( .D(n5738), .CK(clock), .Q(
        \registres[1][19] ) );
  FLIP_FLOP_D \registres_reg[1][18]  ( .D(n5737), .CK(clock), .Q(
        \registres[1][18] ) );
  FLIP_FLOP_D \registres_reg[1][17]  ( .D(n5736), .CK(clock), .Q(
        \registres[1][17] ) );
  FLIP_FLOP_D \registres_reg[1][16]  ( .D(n5735), .CK(clock), .Q(
        \registres[1][16] ) );
  FLIP_FLOP_D \registres_reg[1][15]  ( .D(n5734), .CK(clock), .Q(
        \registres[1][15] ) );
  FLIP_FLOP_D \registres_reg[1][14]  ( .D(n5733), .CK(clock), .Q(
        \registres[1][14] ) );
  FLIP_FLOP_D \registres_reg[1][13]  ( .D(n5732), .CK(clock), .Q(
        \registres[1][13] ) );
  FLIP_FLOP_D \registres_reg[1][12]  ( .D(n5731), .CK(clock), .Q(
        \registres[1][12] ) );
  FLIP_FLOP_D \registres_reg[1][11]  ( .D(n5730), .CK(clock), .Q(
        \registres[1][11] ) );
  FLIP_FLOP_D \registres_reg[1][10]  ( .D(n5729), .CK(clock), .Q(
        \registres[1][10] ) );
  FLIP_FLOP_D \registres_reg[1][9]  ( .D(n5728), .CK(clock), .Q(
        \registres[1][9] ) );
  FLIP_FLOP_D \registres_reg[1][8]  ( .D(n5727), .CK(clock), .Q(
        \registres[1][8] ) );
  FLIP_FLOP_D \registres_reg[1][7]  ( .D(n5726), .CK(clock), .Q(
        \registres[1][7] ) );
  FLIP_FLOP_D \registres_reg[1][6]  ( .D(n5725), .CK(clock), .Q(
        \registres[1][6] ) );
  FLIP_FLOP_D \registres_reg[1][5]  ( .D(n5724), .CK(clock), .Q(
        \registres[1][5] ) );
  FLIP_FLOP_D \registres_reg[1][4]  ( .D(n5723), .CK(clock), .Q(
        \registres[1][4] ) );
  FLIP_FLOP_D \registres_reg[1][3]  ( .D(n5722), .CK(clock), .Q(
        \registres[1][3] ) );
  FLIP_FLOP_D \registres_reg[1][2]  ( .D(n5721), .CK(clock), .Q(
        \registres[1][2] ) );
  FLIP_FLOP_D \registres_reg[1][1]  ( .D(n5720), .CK(clock), .Q(
        \registres[1][1] ) );
  FLIP_FLOP_D \registres_reg[1][0]  ( .D(n5719), .CK(clock), .Q(
        \registres[1][0] ) );
  FLIP_FLOP_D \registres_reg[2][31]  ( .D(n5718), .CK(clock), .Q(
        \registres[2][31] ) );
  FLIP_FLOP_D \registres_reg[2][30]  ( .D(n5717), .CK(clock), .Q(
        \registres[2][30] ) );
  FLIP_FLOP_D \registres_reg[2][29]  ( .D(n5716), .CK(clock), .Q(
        \registres[2][29] ) );
  FLIP_FLOP_D \registres_reg[2][28]  ( .D(n5715), .CK(clock), .Q(
        \registres[2][28] ) );
  FLIP_FLOP_D \registres_reg[2][27]  ( .D(n5714), .CK(clock), .Q(
        \registres[2][27] ) );
  FLIP_FLOP_D \registres_reg[2][26]  ( .D(n5713), .CK(clock), .Q(
        \registres[2][26] ) );
  FLIP_FLOP_D \registres_reg[2][25]  ( .D(n5712), .CK(clock), .Q(
        \registres[2][25] ) );
  FLIP_FLOP_D \registres_reg[2][24]  ( .D(n5711), .CK(clock), .Q(
        \registres[2][24] ) );
  FLIP_FLOP_D \registres_reg[2][23]  ( .D(n5710), .CK(clock), .Q(
        \registres[2][23] ) );
  FLIP_FLOP_D \registres_reg[2][22]  ( .D(n5709), .CK(clock), .Q(
        \registres[2][22] ) );
  FLIP_FLOP_D \registres_reg[2][21]  ( .D(n5708), .CK(clock), .Q(
        \registres[2][21] ) );
  FLIP_FLOP_D \registres_reg[2][20]  ( .D(n5707), .CK(clock), .Q(
        \registres[2][20] ) );
  FLIP_FLOP_D \registres_reg[2][19]  ( .D(n5706), .CK(clock), .Q(
        \registres[2][19] ) );
  FLIP_FLOP_D \registres_reg[2][18]  ( .D(n5705), .CK(clock), .Q(
        \registres[2][18] ) );
  FLIP_FLOP_D \registres_reg[2][17]  ( .D(n5704), .CK(clock), .Q(
        \registres[2][17] ) );
  FLIP_FLOP_D \registres_reg[2][16]  ( .D(n5703), .CK(clock), .Q(
        \registres[2][16] ) );
  FLIP_FLOP_D \registres_reg[2][15]  ( .D(n5702), .CK(clock), .Q(
        \registres[2][15] ) );
  FLIP_FLOP_D \registres_reg[2][14]  ( .D(n5701), .CK(clock), .Q(
        \registres[2][14] ) );
  FLIP_FLOP_D \registres_reg[2][13]  ( .D(n5700), .CK(clock), .Q(
        \registres[2][13] ) );
  FLIP_FLOP_D \registres_reg[2][12]  ( .D(n5699), .CK(clock), .Q(
        \registres[2][12] ) );
  FLIP_FLOP_D \registres_reg[2][11]  ( .D(n5698), .CK(clock), .Q(
        \registres[2][11] ) );
  FLIP_FLOP_D \registres_reg[2][10]  ( .D(n5697), .CK(clock), .Q(
        \registres[2][10] ) );
  FLIP_FLOP_D \registres_reg[2][9]  ( .D(n5696), .CK(clock), .Q(
        \registres[2][9] ) );
  FLIP_FLOP_D \registres_reg[2][8]  ( .D(n5695), .CK(clock), .Q(
        \registres[2][8] ) );
  FLIP_FLOP_D \registres_reg[2][7]  ( .D(n5694), .CK(clock), .Q(
        \registres[2][7] ) );
  FLIP_FLOP_D \registres_reg[2][6]  ( .D(n5693), .CK(clock), .Q(
        \registres[2][6] ) );
  FLIP_FLOP_D \registres_reg[2][5]  ( .D(n5692), .CK(clock), .Q(
        \registres[2][5] ) );
  FLIP_FLOP_D \registres_reg[2][4]  ( .D(n5691), .CK(clock), .Q(
        \registres[2][4] ) );
  FLIP_FLOP_D \registres_reg[2][3]  ( .D(n5690), .CK(clock), .Q(
        \registres[2][3] ) );
  FLIP_FLOP_D \registres_reg[2][2]  ( .D(n5689), .CK(clock), .Q(
        \registres[2][2] ) );
  FLIP_FLOP_D \registres_reg[2][1]  ( .D(n5688), .CK(clock), .Q(
        \registres[2][1] ) );
  FLIP_FLOP_D \registres_reg[2][0]  ( .D(n5687), .CK(clock), .Q(
        \registres[2][0] ) );
  FLIP_FLOP_D \registres_reg[3][31]  ( .D(n5686), .CK(clock), .Q(
        \registres[3][31] ) );
  FLIP_FLOP_D \registres_reg[3][30]  ( .D(n5685), .CK(clock), .Q(
        \registres[3][30] ) );
  FLIP_FLOP_D \registres_reg[3][29]  ( .D(n5684), .CK(clock), .Q(
        \registres[3][29] ) );
  FLIP_FLOP_D \registres_reg[3][28]  ( .D(n5683), .CK(clock), .Q(
        \registres[3][28] ) );
  FLIP_FLOP_D \registres_reg[3][27]  ( .D(n5682), .CK(clock), .Q(
        \registres[3][27] ) );
  FLIP_FLOP_D \registres_reg[3][26]  ( .D(n5681), .CK(clock), .Q(
        \registres[3][26] ) );
  FLIP_FLOP_D \registres_reg[3][25]  ( .D(n5680), .CK(clock), .Q(
        \registres[3][25] ) );
  FLIP_FLOP_D \registres_reg[3][24]  ( .D(n5679), .CK(clock), .Q(
        \registres[3][24] ) );
  FLIP_FLOP_D \registres_reg[3][23]  ( .D(n5678), .CK(clock), .Q(
        \registres[3][23] ) );
  FLIP_FLOP_D \registres_reg[3][22]  ( .D(n5677), .CK(clock), .Q(
        \registres[3][22] ) );
  FLIP_FLOP_D \registres_reg[3][21]  ( .D(n5676), .CK(clock), .Q(
        \registres[3][21] ) );
  FLIP_FLOP_D \registres_reg[3][20]  ( .D(n5675), .CK(clock), .Q(
        \registres[3][20] ) );
  FLIP_FLOP_D \registres_reg[3][19]  ( .D(n5674), .CK(clock), .Q(
        \registres[3][19] ) );
  FLIP_FLOP_D \registres_reg[3][18]  ( .D(n5673), .CK(clock), .Q(
        \registres[3][18] ) );
  FLIP_FLOP_D \registres_reg[3][17]  ( .D(n5672), .CK(clock), .Q(
        \registres[3][17] ) );
  FLIP_FLOP_D \registres_reg[3][16]  ( .D(n5671), .CK(clock), .Q(
        \registres[3][16] ) );
  FLIP_FLOP_D \registres_reg[3][15]  ( .D(n5670), .CK(clock), .Q(
        \registres[3][15] ) );
  FLIP_FLOP_D \registres_reg[3][14]  ( .D(n5669), .CK(clock), .Q(
        \registres[3][14] ) );
  FLIP_FLOP_D \registres_reg[3][13]  ( .D(n5668), .CK(clock), .Q(
        \registres[3][13] ) );
  FLIP_FLOP_D \registres_reg[3][12]  ( .D(n5667), .CK(clock), .Q(
        \registres[3][12] ) );
  FLIP_FLOP_D \registres_reg[3][11]  ( .D(n5666), .CK(clock), .Q(
        \registres[3][11] ) );
  FLIP_FLOP_D \registres_reg[3][10]  ( .D(n5665), .CK(clock), .Q(
        \registres[3][10] ) );
  FLIP_FLOP_D \registres_reg[3][9]  ( .D(n5664), .CK(clock), .Q(
        \registres[3][9] ) );
  FLIP_FLOP_D \registres_reg[3][8]  ( .D(n5663), .CK(clock), .Q(
        \registres[3][8] ) );
  FLIP_FLOP_D \registres_reg[3][7]  ( .D(n5662), .CK(clock), .Q(
        \registres[3][7] ) );
  FLIP_FLOP_D \registres_reg[3][6]  ( .D(n5661), .CK(clock), .Q(
        \registres[3][6] ) );
  FLIP_FLOP_D \registres_reg[3][5]  ( .D(n5660), .CK(clock), .Q(
        \registres[3][5] ) );
  FLIP_FLOP_D \registres_reg[3][4]  ( .D(n5659), .CK(clock), .Q(
        \registres[3][4] ) );
  FLIP_FLOP_D \registres_reg[3][3]  ( .D(n5658), .CK(clock), .Q(
        \registres[3][3] ) );
  FLIP_FLOP_D \registres_reg[3][2]  ( .D(n5657), .CK(clock), .Q(
        \registres[3][2] ) );
  FLIP_FLOP_D \registres_reg[3][1]  ( .D(n5656), .CK(clock), .Q(
        \registres[3][1] ) );
  FLIP_FLOP_D \registres_reg[3][0]  ( .D(n5655), .CK(clock), .Q(
        \registres[3][0] ) );
  FLIP_FLOP_D \registres_reg[4][31]  ( .D(n5654), .CK(clock), .Q(
        \registres[4][31] ) );
  FLIP_FLOP_D \registres_reg[4][30]  ( .D(n5653), .CK(clock), .Q(
        \registres[4][30] ) );
  FLIP_FLOP_D \registres_reg[4][29]  ( .D(n5652), .CK(clock), .Q(
        \registres[4][29] ) );
  FLIP_FLOP_D \registres_reg[4][28]  ( .D(n5651), .CK(clock), .Q(
        \registres[4][28] ) );
  FLIP_FLOP_D \registres_reg[4][27]  ( .D(n5650), .CK(clock), .Q(
        \registres[4][27] ) );
  FLIP_FLOP_D \registres_reg[4][26]  ( .D(n5649), .CK(clock), .Q(
        \registres[4][26] ) );
  FLIP_FLOP_D \registres_reg[4][25]  ( .D(n5648), .CK(clock), .Q(
        \registres[4][25] ) );
  FLIP_FLOP_D \registres_reg[4][24]  ( .D(n5647), .CK(clock), .Q(
        \registres[4][24] ) );
  FLIP_FLOP_D \registres_reg[4][23]  ( .D(n5646), .CK(clock), .Q(
        \registres[4][23] ) );
  FLIP_FLOP_D \registres_reg[4][22]  ( .D(n5645), .CK(clock), .Q(
        \registres[4][22] ) );
  FLIP_FLOP_D \registres_reg[4][21]  ( .D(n5644), .CK(clock), .Q(
        \registres[4][21] ) );
  FLIP_FLOP_D \registres_reg[4][20]  ( .D(n5643), .CK(clock), .Q(
        \registres[4][20] ) );
  FLIP_FLOP_D \registres_reg[4][19]  ( .D(n5642), .CK(clock), .Q(
        \registres[4][19] ) );
  FLIP_FLOP_D \registres_reg[4][18]  ( .D(n5641), .CK(clock), .Q(
        \registres[4][18] ) );
  FLIP_FLOP_D \registres_reg[4][17]  ( .D(n5640), .CK(clock), .Q(
        \registres[4][17] ) );
  FLIP_FLOP_D \registres_reg[4][16]  ( .D(n5639), .CK(clock), .Q(
        \registres[4][16] ) );
  FLIP_FLOP_D \registres_reg[4][15]  ( .D(n5638), .CK(clock), .Q(
        \registres[4][15] ) );
  FLIP_FLOP_D \registres_reg[4][14]  ( .D(n5637), .CK(clock), .Q(
        \registres[4][14] ) );
  FLIP_FLOP_D \registres_reg[4][13]  ( .D(n5636), .CK(clock), .Q(
        \registres[4][13] ) );
  FLIP_FLOP_D \registres_reg[4][12]  ( .D(n5635), .CK(clock), .Q(
        \registres[4][12] ) );
  FLIP_FLOP_D \registres_reg[4][11]  ( .D(n5634), .CK(clock), .Q(
        \registres[4][11] ) );
  FLIP_FLOP_D \registres_reg[4][10]  ( .D(n5633), .CK(clock), .Q(
        \registres[4][10] ) );
  FLIP_FLOP_D \registres_reg[4][9]  ( .D(n5632), .CK(clock), .Q(
        \registres[4][9] ) );
  FLIP_FLOP_D \registres_reg[4][8]  ( .D(n5631), .CK(clock), .Q(
        \registres[4][8] ) );
  FLIP_FLOP_D \registres_reg[4][7]  ( .D(n5630), .CK(clock), .Q(
        \registres[4][7] ) );
  FLIP_FLOP_D \registres_reg[4][6]  ( .D(n5629), .CK(clock), .Q(
        \registres[4][6] ) );
  FLIP_FLOP_D \registres_reg[4][5]  ( .D(n5628), .CK(clock), .Q(
        \registres[4][5] ) );
  FLIP_FLOP_D \registres_reg[4][4]  ( .D(n5627), .CK(clock), .Q(
        \registres[4][4] ) );
  FLIP_FLOP_D \registres_reg[4][3]  ( .D(n5626), .CK(clock), .Q(
        \registres[4][3] ) );
  FLIP_FLOP_D \registres_reg[4][2]  ( .D(n5625), .CK(clock), .Q(
        \registres[4][2] ) );
  FLIP_FLOP_D \registres_reg[4][1]  ( .D(n5624), .CK(clock), .Q(
        \registres[4][1] ) );
  FLIP_FLOP_D \registres_reg[4][0]  ( .D(n5623), .CK(clock), .Q(
        \registres[4][0] ) );
  FLIP_FLOP_D \registres_reg[5][31]  ( .D(n5622), .CK(clock), .Q(
        \registres[5][31] ) );
  FLIP_FLOP_D \registres_reg[5][30]  ( .D(n5621), .CK(clock), .Q(
        \registres[5][30] ) );
  FLIP_FLOP_D \registres_reg[5][29]  ( .D(n5620), .CK(clock), .Q(
        \registres[5][29] ) );
  FLIP_FLOP_D \registres_reg[5][28]  ( .D(n5619), .CK(clock), .Q(
        \registres[5][28] ) );
  FLIP_FLOP_D \registres_reg[5][27]  ( .D(n5618), .CK(clock), .Q(
        \registres[5][27] ) );
  FLIP_FLOP_D \registres_reg[5][26]  ( .D(n5617), .CK(clock), .Q(
        \registres[5][26] ) );
  FLIP_FLOP_D \registres_reg[5][25]  ( .D(n5616), .CK(clock), .Q(
        \registres[5][25] ) );
  FLIP_FLOP_D \registres_reg[5][24]  ( .D(n5615), .CK(clock), .Q(
        \registres[5][24] ) );
  FLIP_FLOP_D \registres_reg[5][23]  ( .D(n5614), .CK(clock), .Q(
        \registres[5][23] ) );
  FLIP_FLOP_D \registres_reg[5][22]  ( .D(n5613), .CK(clock), .Q(
        \registres[5][22] ) );
  FLIP_FLOP_D \registres_reg[5][21]  ( .D(n5612), .CK(clock), .Q(
        \registres[5][21] ) );
  FLIP_FLOP_D \registres_reg[5][20]  ( .D(n5611), .CK(clock), .Q(
        \registres[5][20] ) );
  FLIP_FLOP_D \registres_reg[5][19]  ( .D(n5610), .CK(clock), .Q(
        \registres[5][19] ) );
  FLIP_FLOP_D \registres_reg[5][18]  ( .D(n5609), .CK(clock), .Q(
        \registres[5][18] ) );
  FLIP_FLOP_D \registres_reg[5][17]  ( .D(n5608), .CK(clock), .Q(
        \registres[5][17] ) );
  FLIP_FLOP_D \registres_reg[5][16]  ( .D(n5607), .CK(clock), .Q(
        \registres[5][16] ) );
  FLIP_FLOP_D \registres_reg[5][15]  ( .D(n5606), .CK(clock), .Q(
        \registres[5][15] ) );
  FLIP_FLOP_D \registres_reg[5][14]  ( .D(n5605), .CK(clock), .Q(
        \registres[5][14] ) );
  FLIP_FLOP_D \registres_reg[5][13]  ( .D(n5604), .CK(clock), .Q(
        \registres[5][13] ) );
  FLIP_FLOP_D \registres_reg[5][12]  ( .D(n5603), .CK(clock), .Q(
        \registres[5][12] ) );
  FLIP_FLOP_D \registres_reg[5][11]  ( .D(n5602), .CK(clock), .Q(
        \registres[5][11] ) );
  FLIP_FLOP_D \registres_reg[5][10]  ( .D(n5601), .CK(clock), .Q(
        \registres[5][10] ) );
  FLIP_FLOP_D \registres_reg[5][9]  ( .D(n5600), .CK(clock), .Q(
        \registres[5][9] ) );
  FLIP_FLOP_D \registres_reg[5][8]  ( .D(n5599), .CK(clock), .Q(
        \registres[5][8] ) );
  FLIP_FLOP_D \registres_reg[5][7]  ( .D(n5598), .CK(clock), .Q(
        \registres[5][7] ) );
  FLIP_FLOP_D \registres_reg[5][6]  ( .D(n5597), .CK(clock), .Q(
        \registres[5][6] ) );
  FLIP_FLOP_D \registres_reg[5][5]  ( .D(n5596), .CK(clock), .Q(
        \registres[5][5] ) );
  FLIP_FLOP_D \registres_reg[5][4]  ( .D(n5595), .CK(clock), .Q(
        \registres[5][4] ) );
  FLIP_FLOP_D \registres_reg[5][3]  ( .D(n5594), .CK(clock), .Q(
        \registres[5][3] ) );
  FLIP_FLOP_D \registres_reg[5][2]  ( .D(n5593), .CK(clock), .Q(
        \registres[5][2] ) );
  FLIP_FLOP_D \registres_reg[5][1]  ( .D(n5592), .CK(clock), .Q(
        \registres[5][1] ) );
  FLIP_FLOP_D \registres_reg[5][0]  ( .D(n5591), .CK(clock), .Q(
        \registres[5][0] ) );
  FLIP_FLOP_D \registres_reg[6][31]  ( .D(n5590), .CK(clock), .Q(
        \registres[6][31] ) );
  FLIP_FLOP_D \registres_reg[6][30]  ( .D(n5589), .CK(clock), .Q(
        \registres[6][30] ) );
  FLIP_FLOP_D \registres_reg[6][29]  ( .D(n5588), .CK(clock), .Q(
        \registres[6][29] ) );
  FLIP_FLOP_D \registres_reg[6][28]  ( .D(n5587), .CK(clock), .Q(
        \registres[6][28] ) );
  FLIP_FLOP_D \registres_reg[6][27]  ( .D(n5586), .CK(clock), .Q(
        \registres[6][27] ) );
  FLIP_FLOP_D \registres_reg[6][26]  ( .D(n5585), .CK(clock), .Q(
        \registres[6][26] ) );
  FLIP_FLOP_D \registres_reg[6][25]  ( .D(n5584), .CK(clock), .Q(
        \registres[6][25] ) );
  FLIP_FLOP_D \registres_reg[6][24]  ( .D(n5583), .CK(clock), .Q(
        \registres[6][24] ) );
  FLIP_FLOP_D \registres_reg[6][23]  ( .D(n5582), .CK(clock), .Q(
        \registres[6][23] ) );
  FLIP_FLOP_D \registres_reg[6][22]  ( .D(n5581), .CK(clock), .Q(
        \registres[6][22] ) );
  FLIP_FLOP_D \registres_reg[6][21]  ( .D(n5580), .CK(clock), .Q(
        \registres[6][21] ) );
  FLIP_FLOP_D \registres_reg[6][20]  ( .D(n5579), .CK(clock), .Q(
        \registres[6][20] ) );
  FLIP_FLOP_D \registres_reg[6][19]  ( .D(n5578), .CK(clock), .Q(
        \registres[6][19] ) );
  FLIP_FLOP_D \registres_reg[6][18]  ( .D(n5577), .CK(clock), .Q(
        \registres[6][18] ) );
  FLIP_FLOP_D \registres_reg[6][17]  ( .D(n5576), .CK(clock), .Q(
        \registres[6][17] ) );
  FLIP_FLOP_D \registres_reg[6][16]  ( .D(n5575), .CK(clock), .Q(
        \registres[6][16] ) );
  FLIP_FLOP_D \registres_reg[6][15]  ( .D(n5574), .CK(clock), .Q(
        \registres[6][15] ) );
  FLIP_FLOP_D \registres_reg[6][14]  ( .D(n5573), .CK(clock), .Q(
        \registres[6][14] ) );
  FLIP_FLOP_D \registres_reg[6][13]  ( .D(n5572), .CK(clock), .Q(
        \registres[6][13] ) );
  FLIP_FLOP_D \registres_reg[6][12]  ( .D(n5571), .CK(clock), .Q(
        \registres[6][12] ) );
  FLIP_FLOP_D \registres_reg[6][11]  ( .D(n5570), .CK(clock), .Q(
        \registres[6][11] ) );
  FLIP_FLOP_D \registres_reg[6][10]  ( .D(n5569), .CK(clock), .Q(
        \registres[6][10] ) );
  FLIP_FLOP_D \registres_reg[6][9]  ( .D(n5568), .CK(clock), .Q(
        \registres[6][9] ) );
  FLIP_FLOP_D \registres_reg[6][8]  ( .D(n5567), .CK(clock), .Q(
        \registres[6][8] ) );
  FLIP_FLOP_D \registres_reg[6][7]  ( .D(n5566), .CK(clock), .Q(
        \registres[6][7] ) );
  FLIP_FLOP_D \registres_reg[6][6]  ( .D(n5565), .CK(clock), .Q(
        \registres[6][6] ) );
  FLIP_FLOP_D \registres_reg[6][5]  ( .D(n5564), .CK(clock), .Q(
        \registres[6][5] ) );
  FLIP_FLOP_D \registres_reg[6][4]  ( .D(n5563), .CK(clock), .Q(
        \registres[6][4] ) );
  FLIP_FLOP_D \registres_reg[6][3]  ( .D(n5562), .CK(clock), .Q(
        \registres[6][3] ) );
  FLIP_FLOP_D \registres_reg[6][2]  ( .D(n5561), .CK(clock), .Q(
        \registres[6][2] ) );
  FLIP_FLOP_D \registres_reg[6][1]  ( .D(n5560), .CK(clock), .Q(
        \registres[6][1] ) );
  FLIP_FLOP_D \registres_reg[6][0]  ( .D(n5559), .CK(clock), .Q(
        \registres[6][0] ) );
  FLIP_FLOP_D \registres_reg[7][31]  ( .D(n5558), .CK(clock), .Q(
        \registres[7][31] ) );
  FLIP_FLOP_D \registres_reg[7][30]  ( .D(n5557), .CK(clock), .Q(
        \registres[7][30] ) );
  FLIP_FLOP_D \registres_reg[7][29]  ( .D(n5556), .CK(clock), .Q(
        \registres[7][29] ) );
  FLIP_FLOP_D \registres_reg[7][28]  ( .D(n5555), .CK(clock), .Q(
        \registres[7][28] ) );
  FLIP_FLOP_D \registres_reg[7][27]  ( .D(n5554), .CK(clock), .Q(
        \registres[7][27] ) );
  FLIP_FLOP_D \registres_reg[7][26]  ( .D(n5553), .CK(clock), .Q(
        \registres[7][26] ) );
  FLIP_FLOP_D \registres_reg[7][25]  ( .D(n5552), .CK(clock), .Q(
        \registres[7][25] ) );
  FLIP_FLOP_D \registres_reg[7][24]  ( .D(n5551), .CK(clock), .Q(
        \registres[7][24] ) );
  FLIP_FLOP_D \registres_reg[7][23]  ( .D(n5550), .CK(clock), .Q(
        \registres[7][23] ) );
  FLIP_FLOP_D \registres_reg[7][22]  ( .D(n5549), .CK(clock), .Q(
        \registres[7][22] ) );
  FLIP_FLOP_D \registres_reg[7][21]  ( .D(n5548), .CK(clock), .Q(
        \registres[7][21] ) );
  FLIP_FLOP_D \registres_reg[7][20]  ( .D(n5547), .CK(clock), .Q(
        \registres[7][20] ) );
  FLIP_FLOP_D \registres_reg[7][19]  ( .D(n5546), .CK(clock), .Q(
        \registres[7][19] ) );
  FLIP_FLOP_D \registres_reg[7][18]  ( .D(n5545), .CK(clock), .Q(
        \registres[7][18] ) );
  FLIP_FLOP_D \registres_reg[7][17]  ( .D(n5544), .CK(clock), .Q(
        \registres[7][17] ) );
  FLIP_FLOP_D \registres_reg[7][16]  ( .D(n5543), .CK(clock), .Q(
        \registres[7][16] ) );
  FLIP_FLOP_D \registres_reg[7][15]  ( .D(n5542), .CK(clock), .Q(
        \registres[7][15] ) );
  FLIP_FLOP_D \registres_reg[7][14]  ( .D(n5541), .CK(clock), .Q(
        \registres[7][14] ) );
  FLIP_FLOP_D \registres_reg[7][13]  ( .D(n5540), .CK(clock), .Q(
        \registres[7][13] ) );
  FLIP_FLOP_D \registres_reg[7][12]  ( .D(n5539), .CK(clock), .Q(
        \registres[7][12] ) );
  FLIP_FLOP_D \registres_reg[7][11]  ( .D(n5538), .CK(clock), .Q(
        \registres[7][11] ) );
  FLIP_FLOP_D \registres_reg[7][10]  ( .D(n5537), .CK(clock), .Q(
        \registres[7][10] ) );
  FLIP_FLOP_D \registres_reg[7][9]  ( .D(n5536), .CK(clock), .Q(
        \registres[7][9] ) );
  FLIP_FLOP_D \registres_reg[7][8]  ( .D(n5535), .CK(clock), .Q(
        \registres[7][8] ) );
  FLIP_FLOP_D \registres_reg[7][7]  ( .D(n5534), .CK(clock), .Q(
        \registres[7][7] ) );
  FLIP_FLOP_D \registres_reg[7][6]  ( .D(n5533), .CK(clock), .Q(
        \registres[7][6] ) );
  FLIP_FLOP_D \registres_reg[7][5]  ( .D(n5532), .CK(clock), .Q(
        \registres[7][5] ) );
  FLIP_FLOP_D \registres_reg[7][4]  ( .D(n5531), .CK(clock), .Q(
        \registres[7][4] ) );
  FLIP_FLOP_D \registres_reg[7][3]  ( .D(n5530), .CK(clock), .Q(
        \registres[7][3] ) );
  FLIP_FLOP_D \registres_reg[7][2]  ( .D(n5529), .CK(clock), .Q(
        \registres[7][2] ) );
  FLIP_FLOP_D \registres_reg[7][1]  ( .D(n5528), .CK(clock), .Q(
        \registres[7][1] ) );
  FLIP_FLOP_D \registres_reg[7][0]  ( .D(n5527), .CK(clock), .Q(
        \registres[7][0] ) );
  FLIP_FLOP_D \registres_reg[8][31]  ( .D(n5526), .CK(clock), .Q(
        \registres[8][31] ) );
  FLIP_FLOP_D \registres_reg[8][30]  ( .D(n5525), .CK(clock), .Q(
        \registres[8][30] ) );
  FLIP_FLOP_D \registres_reg[8][29]  ( .D(n5524), .CK(clock), .Q(
        \registres[8][29] ) );
  FLIP_FLOP_D \registres_reg[8][28]  ( .D(n5523), .CK(clock), .Q(
        \registres[8][28] ) );
  FLIP_FLOP_D \registres_reg[8][27]  ( .D(n5522), .CK(clock), .Q(
        \registres[8][27] ) );
  FLIP_FLOP_D \registres_reg[8][26]  ( .D(n5521), .CK(clock), .Q(
        \registres[8][26] ) );
  FLIP_FLOP_D \registres_reg[8][25]  ( .D(n5520), .CK(clock), .Q(
        \registres[8][25] ) );
  FLIP_FLOP_D \registres_reg[8][24]  ( .D(n5519), .CK(clock), .Q(
        \registres[8][24] ) );
  FLIP_FLOP_D \registres_reg[8][23]  ( .D(n5518), .CK(clock), .Q(
        \registres[8][23] ) );
  FLIP_FLOP_D \registres_reg[8][22]  ( .D(n5517), .CK(clock), .Q(
        \registres[8][22] ) );
  FLIP_FLOP_D \registres_reg[8][21]  ( .D(n5516), .CK(clock), .Q(
        \registres[8][21] ) );
  FLIP_FLOP_D \registres_reg[8][20]  ( .D(n5515), .CK(clock), .Q(
        \registres[8][20] ) );
  FLIP_FLOP_D \registres_reg[8][19]  ( .D(n5514), .CK(clock), .Q(
        \registres[8][19] ) );
  FLIP_FLOP_D \registres_reg[8][18]  ( .D(n5513), .CK(clock), .Q(
        \registres[8][18] ) );
  FLIP_FLOP_D \registres_reg[8][17]  ( .D(n5512), .CK(clock), .Q(
        \registres[8][17] ) );
  FLIP_FLOP_D \registres_reg[8][16]  ( .D(n5511), .CK(clock), .Q(
        \registres[8][16] ) );
  FLIP_FLOP_D \registres_reg[8][15]  ( .D(n5510), .CK(clock), .Q(
        \registres[8][15] ) );
  FLIP_FLOP_D \registres_reg[8][14]  ( .D(n5509), .CK(clock), .Q(
        \registres[8][14] ) );
  FLIP_FLOP_D \registres_reg[8][13]  ( .D(n5508), .CK(clock), .Q(
        \registres[8][13] ) );
  FLIP_FLOP_D \registres_reg[8][12]  ( .D(n5507), .CK(clock), .Q(
        \registres[8][12] ) );
  FLIP_FLOP_D \registres_reg[8][11]  ( .D(n5506), .CK(clock), .Q(
        \registres[8][11] ) );
  FLIP_FLOP_D \registres_reg[8][10]  ( .D(n5505), .CK(clock), .Q(
        \registres[8][10] ) );
  FLIP_FLOP_D \registres_reg[8][9]  ( .D(n5504), .CK(clock), .Q(
        \registres[8][9] ) );
  FLIP_FLOP_D \registres_reg[8][8]  ( .D(n5503), .CK(clock), .Q(
        \registres[8][8] ) );
  FLIP_FLOP_D \registres_reg[8][7]  ( .D(n5502), .CK(clock), .Q(
        \registres[8][7] ) );
  FLIP_FLOP_D \registres_reg[8][6]  ( .D(n5501), .CK(clock), .Q(
        \registres[8][6] ) );
  FLIP_FLOP_D \registres_reg[8][5]  ( .D(n5500), .CK(clock), .Q(
        \registres[8][5] ) );
  FLIP_FLOP_D \registres_reg[8][4]  ( .D(n5499), .CK(clock), .Q(
        \registres[8][4] ) );
  FLIP_FLOP_D \registres_reg[8][3]  ( .D(n5498), .CK(clock), .Q(
        \registres[8][3] ) );
  FLIP_FLOP_D \registres_reg[8][2]  ( .D(n5497), .CK(clock), .Q(
        \registres[8][2] ) );
  FLIP_FLOP_D \registres_reg[8][1]  ( .D(n5496), .CK(clock), .Q(
        \registres[8][1] ) );
  FLIP_FLOP_D \registres_reg[8][0]  ( .D(n5495), .CK(clock), .Q(
        \registres[8][0] ) );
  FLIP_FLOP_D \registres_reg[9][31]  ( .D(n5494), .CK(clock), .Q(
        \registres[9][31] ) );
  FLIP_FLOP_D \registres_reg[9][30]  ( .D(n5493), .CK(clock), .Q(
        \registres[9][30] ) );
  FLIP_FLOP_D \registres_reg[9][29]  ( .D(n5492), .CK(clock), .Q(
        \registres[9][29] ) );
  FLIP_FLOP_D \registres_reg[9][28]  ( .D(n5491), .CK(clock), .Q(
        \registres[9][28] ) );
  FLIP_FLOP_D \registres_reg[9][27]  ( .D(n5490), .CK(clock), .Q(
        \registres[9][27] ) );
  FLIP_FLOP_D \registres_reg[9][26]  ( .D(n5489), .CK(clock), .Q(
        \registres[9][26] ) );
  FLIP_FLOP_D \registres_reg[9][25]  ( .D(n5488), .CK(clock), .Q(
        \registres[9][25] ) );
  FLIP_FLOP_D \registres_reg[9][24]  ( .D(n5487), .CK(clock), .Q(
        \registres[9][24] ) );
  FLIP_FLOP_D \registres_reg[9][23]  ( .D(n5486), .CK(clock), .Q(
        \registres[9][23] ) );
  FLIP_FLOP_D \registres_reg[9][22]  ( .D(n5485), .CK(clock), .Q(
        \registres[9][22] ) );
  FLIP_FLOP_D \registres_reg[9][21]  ( .D(n5484), .CK(clock), .Q(
        \registres[9][21] ) );
  FLIP_FLOP_D \registres_reg[9][20]  ( .D(n5483), .CK(clock), .Q(
        \registres[9][20] ) );
  FLIP_FLOP_D \registres_reg[9][19]  ( .D(n5482), .CK(clock), .Q(
        \registres[9][19] ) );
  FLIP_FLOP_D \registres_reg[9][18]  ( .D(n5481), .CK(clock), .Q(
        \registres[9][18] ) );
  FLIP_FLOP_D \registres_reg[9][17]  ( .D(n5480), .CK(clock), .Q(
        \registres[9][17] ) );
  FLIP_FLOP_D \registres_reg[9][16]  ( .D(n5479), .CK(clock), .Q(
        \registres[9][16] ) );
  FLIP_FLOP_D \registres_reg[9][15]  ( .D(n5478), .CK(clock), .Q(
        \registres[9][15] ) );
  FLIP_FLOP_D \registres_reg[9][14]  ( .D(n5477), .CK(clock), .Q(
        \registres[9][14] ) );
  FLIP_FLOP_D \registres_reg[9][13]  ( .D(n5476), .CK(clock), .Q(
        \registres[9][13] ) );
  FLIP_FLOP_D \registres_reg[9][12]  ( .D(n5475), .CK(clock), .Q(
        \registres[9][12] ) );
  FLIP_FLOP_D \registres_reg[9][11]  ( .D(n5474), .CK(clock), .Q(
        \registres[9][11] ) );
  FLIP_FLOP_D \registres_reg[9][10]  ( .D(n5473), .CK(clock), .Q(
        \registres[9][10] ) );
  FLIP_FLOP_D \registres_reg[9][9]  ( .D(n5472), .CK(clock), .Q(
        \registres[9][9] ) );
  FLIP_FLOP_D \registres_reg[9][8]  ( .D(n5471), .CK(clock), .Q(
        \registres[9][8] ) );
  FLIP_FLOP_D \registres_reg[9][7]  ( .D(n5470), .CK(clock), .Q(
        \registres[9][7] ) );
  FLIP_FLOP_D \registres_reg[9][6]  ( .D(n5469), .CK(clock), .Q(
        \registres[9][6] ) );
  FLIP_FLOP_D \registres_reg[9][5]  ( .D(n5468), .CK(clock), .Q(
        \registres[9][5] ) );
  FLIP_FLOP_D \registres_reg[9][4]  ( .D(n5467), .CK(clock), .Q(
        \registres[9][4] ) );
  FLIP_FLOP_D \registres_reg[9][3]  ( .D(n5466), .CK(clock), .Q(
        \registres[9][3] ) );
  FLIP_FLOP_D \registres_reg[9][2]  ( .D(n5465), .CK(clock), .Q(
        \registres[9][2] ) );
  FLIP_FLOP_D \registres_reg[9][1]  ( .D(n5464), .CK(clock), .Q(
        \registres[9][1] ) );
  FLIP_FLOP_D \registres_reg[9][0]  ( .D(n5463), .CK(clock), .Q(
        \registres[9][0] ) );
  FLIP_FLOP_D \registres_reg[10][31]  ( .D(n5462), .CK(clock), .Q(
        \registres[10][31] ) );
  FLIP_FLOP_D \registres_reg[10][30]  ( .D(n5461), .CK(clock), .Q(
        \registres[10][30] ) );
  FLIP_FLOP_D \registres_reg[10][29]  ( .D(n5460), .CK(clock), .Q(
        \registres[10][29] ) );
  FLIP_FLOP_D \registres_reg[10][28]  ( .D(n5459), .CK(clock), .Q(
        \registres[10][28] ) );
  FLIP_FLOP_D \registres_reg[10][27]  ( .D(n5458), .CK(clock), .Q(
        \registres[10][27] ) );
  FLIP_FLOP_D \registres_reg[10][26]  ( .D(n5457), .CK(clock), .Q(
        \registres[10][26] ) );
  FLIP_FLOP_D \registres_reg[10][25]  ( .D(n5456), .CK(clock), .Q(
        \registres[10][25] ) );
  FLIP_FLOP_D \registres_reg[10][24]  ( .D(n5455), .CK(clock), .Q(
        \registres[10][24] ) );
  FLIP_FLOP_D \registres_reg[10][23]  ( .D(n5454), .CK(clock), .Q(
        \registres[10][23] ) );
  FLIP_FLOP_D \registres_reg[10][22]  ( .D(n5453), .CK(clock), .Q(
        \registres[10][22] ) );
  FLIP_FLOP_D \registres_reg[10][21]  ( .D(n5452), .CK(clock), .Q(
        \registres[10][21] ) );
  FLIP_FLOP_D \registres_reg[10][20]  ( .D(n5451), .CK(clock), .Q(
        \registres[10][20] ) );
  FLIP_FLOP_D \registres_reg[10][19]  ( .D(n5450), .CK(clock), .Q(
        \registres[10][19] ) );
  FLIP_FLOP_D \registres_reg[10][18]  ( .D(n5449), .CK(clock), .Q(
        \registres[10][18] ) );
  FLIP_FLOP_D \registres_reg[10][17]  ( .D(n5448), .CK(clock), .Q(
        \registres[10][17] ) );
  FLIP_FLOP_D \registres_reg[10][16]  ( .D(n5447), .CK(clock), .Q(
        \registres[10][16] ) );
  FLIP_FLOP_D \registres_reg[10][15]  ( .D(n5446), .CK(clock), .Q(
        \registres[10][15] ) );
  FLIP_FLOP_D \registres_reg[10][14]  ( .D(n5445), .CK(clock), .Q(
        \registres[10][14] ) );
  FLIP_FLOP_D \registres_reg[10][13]  ( .D(n5444), .CK(clock), .Q(
        \registres[10][13] ) );
  FLIP_FLOP_D \registres_reg[10][12]  ( .D(n5443), .CK(clock), .Q(
        \registres[10][12] ) );
  FLIP_FLOP_D \registres_reg[10][11]  ( .D(n5442), .CK(clock), .Q(
        \registres[10][11] ) );
  FLIP_FLOP_D \registres_reg[10][10]  ( .D(n5441), .CK(clock), .Q(
        \registres[10][10] ) );
  FLIP_FLOP_D \registres_reg[10][9]  ( .D(n5440), .CK(clock), .Q(
        \registres[10][9] ) );
  FLIP_FLOP_D \registres_reg[10][8]  ( .D(n5439), .CK(clock), .Q(
        \registres[10][8] ) );
  FLIP_FLOP_D \registres_reg[10][7]  ( .D(n5438), .CK(clock), .Q(
        \registres[10][7] ) );
  FLIP_FLOP_D \registres_reg[10][6]  ( .D(n5437), .CK(clock), .Q(
        \registres[10][6] ) );
  FLIP_FLOP_D \registres_reg[10][5]  ( .D(n5436), .CK(clock), .Q(
        \registres[10][5] ) );
  FLIP_FLOP_D \registres_reg[10][4]  ( .D(n5435), .CK(clock), .Q(
        \registres[10][4] ) );
  FLIP_FLOP_D \registres_reg[10][3]  ( .D(n5434), .CK(clock), .Q(
        \registres[10][3] ) );
  FLIP_FLOP_D \registres_reg[10][2]  ( .D(n5433), .CK(clock), .Q(
        \registres[10][2] ) );
  FLIP_FLOP_D \registres_reg[10][1]  ( .D(n5432), .CK(clock), .Q(
        \registres[10][1] ) );
  FLIP_FLOP_D \registres_reg[10][0]  ( .D(n5431), .CK(clock), .Q(
        \registres[10][0] ) );
  FLIP_FLOP_D \registres_reg[11][31]  ( .D(n5430), .CK(clock), .Q(
        \registres[11][31] ) );
  FLIP_FLOP_D \registres_reg[11][30]  ( .D(n5429), .CK(clock), .Q(
        \registres[11][30] ) );
  FLIP_FLOP_D \registres_reg[11][29]  ( .D(n5428), .CK(clock), .Q(
        \registres[11][29] ) );
  FLIP_FLOP_D \registres_reg[11][28]  ( .D(n5427), .CK(clock), .Q(
        \registres[11][28] ) );
  FLIP_FLOP_D \registres_reg[11][27]  ( .D(n5426), .CK(clock), .Q(
        \registres[11][27] ) );
  FLIP_FLOP_D \registres_reg[11][26]  ( .D(n5425), .CK(clock), .Q(
        \registres[11][26] ) );
  FLIP_FLOP_D \registres_reg[11][25]  ( .D(n5424), .CK(clock), .Q(
        \registres[11][25] ) );
  FLIP_FLOP_D \registres_reg[11][24]  ( .D(n5423), .CK(clock), .Q(
        \registres[11][24] ) );
  FLIP_FLOP_D \registres_reg[11][23]  ( .D(n5422), .CK(clock), .Q(
        \registres[11][23] ) );
  FLIP_FLOP_D \registres_reg[11][22]  ( .D(n5421), .CK(clock), .Q(
        \registres[11][22] ) );
  FLIP_FLOP_D \registres_reg[11][21]  ( .D(n5420), .CK(clock), .Q(
        \registres[11][21] ) );
  FLIP_FLOP_D \registres_reg[11][20]  ( .D(n5419), .CK(clock), .Q(
        \registres[11][20] ) );
  FLIP_FLOP_D \registres_reg[11][19]  ( .D(n5418), .CK(clock), .Q(
        \registres[11][19] ) );
  FLIP_FLOP_D \registres_reg[11][18]  ( .D(n5417), .CK(clock), .Q(
        \registres[11][18] ) );
  FLIP_FLOP_D \registres_reg[11][17]  ( .D(n5416), .CK(clock), .Q(
        \registres[11][17] ) );
  FLIP_FLOP_D \registres_reg[11][16]  ( .D(n5415), .CK(clock), .Q(
        \registres[11][16] ) );
  FLIP_FLOP_D \registres_reg[11][15]  ( .D(n5414), .CK(clock), .Q(
        \registres[11][15] ) );
  FLIP_FLOP_D \registres_reg[11][14]  ( .D(n5413), .CK(clock), .Q(
        \registres[11][14] ) );
  FLIP_FLOP_D \registres_reg[11][13]  ( .D(n5412), .CK(clock), .Q(
        \registres[11][13] ) );
  FLIP_FLOP_D \registres_reg[11][12]  ( .D(n5411), .CK(clock), .Q(
        \registres[11][12] ) );
  FLIP_FLOP_D \registres_reg[11][11]  ( .D(n5410), .CK(clock), .Q(
        \registres[11][11] ) );
  FLIP_FLOP_D \registres_reg[11][10]  ( .D(n5409), .CK(clock), .Q(
        \registres[11][10] ) );
  FLIP_FLOP_D \registres_reg[11][9]  ( .D(n5408), .CK(clock), .Q(
        \registres[11][9] ) );
  FLIP_FLOP_D \registres_reg[11][8]  ( .D(n5407), .CK(clock), .Q(
        \registres[11][8] ) );
  FLIP_FLOP_D \registres_reg[11][7]  ( .D(n5406), .CK(clock), .Q(
        \registres[11][7] ) );
  FLIP_FLOP_D \registres_reg[11][6]  ( .D(n5405), .CK(clock), .Q(
        \registres[11][6] ) );
  FLIP_FLOP_D \registres_reg[11][5]  ( .D(n5404), .CK(clock), .Q(
        \registres[11][5] ) );
  FLIP_FLOP_D \registres_reg[11][4]  ( .D(n5403), .CK(clock), .Q(
        \registres[11][4] ) );
  FLIP_FLOP_D \registres_reg[11][3]  ( .D(n5402), .CK(clock), .Q(
        \registres[11][3] ) );
  FLIP_FLOP_D \registres_reg[11][2]  ( .D(n5401), .CK(clock), .Q(
        \registres[11][2] ) );
  FLIP_FLOP_D \registres_reg[11][1]  ( .D(n5400), .CK(clock), .Q(
        \registres[11][1] ) );
  FLIP_FLOP_D \registres_reg[11][0]  ( .D(n5399), .CK(clock), .Q(
        \registres[11][0] ) );
  FLIP_FLOP_D \registres_reg[12][31]  ( .D(n5398), .CK(clock), .Q(
        \registres[12][31] ) );
  FLIP_FLOP_D \registres_reg[12][30]  ( .D(n5397), .CK(clock), .Q(
        \registres[12][30] ) );
  FLIP_FLOP_D \registres_reg[12][29]  ( .D(n5396), .CK(clock), .Q(
        \registres[12][29] ) );
  FLIP_FLOP_D \registres_reg[12][28]  ( .D(n5395), .CK(clock), .Q(
        \registres[12][28] ) );
  FLIP_FLOP_D \registres_reg[12][27]  ( .D(n5394), .CK(clock), .Q(
        \registres[12][27] ) );
  FLIP_FLOP_D \registres_reg[12][26]  ( .D(n5393), .CK(clock), .Q(
        \registres[12][26] ) );
  FLIP_FLOP_D \registres_reg[12][25]  ( .D(n5392), .CK(clock), .Q(
        \registres[12][25] ) );
  FLIP_FLOP_D \registres_reg[12][24]  ( .D(n5391), .CK(clock), .Q(
        \registres[12][24] ) );
  FLIP_FLOP_D \registres_reg[12][23]  ( .D(n5390), .CK(clock), .Q(
        \registres[12][23] ) );
  FLIP_FLOP_D \registres_reg[12][22]  ( .D(n5389), .CK(clock), .Q(
        \registres[12][22] ) );
  FLIP_FLOP_D \registres_reg[12][21]  ( .D(n5388), .CK(clock), .Q(
        \registres[12][21] ) );
  FLIP_FLOP_D \registres_reg[12][20]  ( .D(n5387), .CK(clock), .Q(
        \registres[12][20] ) );
  FLIP_FLOP_D \registres_reg[12][19]  ( .D(n5386), .CK(clock), .Q(
        \registres[12][19] ) );
  FLIP_FLOP_D \registres_reg[12][18]  ( .D(n5385), .CK(clock), .Q(
        \registres[12][18] ) );
  FLIP_FLOP_D \registres_reg[12][17]  ( .D(n5384), .CK(clock), .Q(
        \registres[12][17] ) );
  FLIP_FLOP_D \registres_reg[12][16]  ( .D(n5383), .CK(clock), .Q(
        \registres[12][16] ) );
  FLIP_FLOP_D \registres_reg[12][15]  ( .D(n5382), .CK(clock), .Q(
        \registres[12][15] ) );
  FLIP_FLOP_D \registres_reg[12][14]  ( .D(n5381), .CK(clock), .Q(
        \registres[12][14] ) );
  FLIP_FLOP_D \registres_reg[12][13]  ( .D(n5380), .CK(clock), .Q(
        \registres[12][13] ) );
  FLIP_FLOP_D \registres_reg[12][12]  ( .D(n5379), .CK(clock), .Q(
        \registres[12][12] ) );
  FLIP_FLOP_D \registres_reg[12][11]  ( .D(n5378), .CK(clock), .Q(
        \registres[12][11] ) );
  FLIP_FLOP_D \registres_reg[12][10]  ( .D(n5377), .CK(clock), .Q(
        \registres[12][10] ) );
  FLIP_FLOP_D \registres_reg[12][9]  ( .D(n5376), .CK(clock), .Q(
        \registres[12][9] ) );
  FLIP_FLOP_D \registres_reg[12][8]  ( .D(n5375), .CK(clock), .Q(
        \registres[12][8] ) );
  FLIP_FLOP_D \registres_reg[12][7]  ( .D(n5374), .CK(clock), .Q(
        \registres[12][7] ) );
  FLIP_FLOP_D \registres_reg[12][6]  ( .D(n5373), .CK(clock), .Q(
        \registres[12][6] ) );
  FLIP_FLOP_D \registres_reg[12][5]  ( .D(n5372), .CK(clock), .Q(
        \registres[12][5] ) );
  FLIP_FLOP_D \registres_reg[12][4]  ( .D(n5371), .CK(clock), .Q(
        \registres[12][4] ) );
  FLIP_FLOP_D \registres_reg[12][3]  ( .D(n5370), .CK(clock), .Q(
        \registres[12][3] ) );
  FLIP_FLOP_D \registres_reg[12][2]  ( .D(n5369), .CK(clock), .Q(
        \registres[12][2] ) );
  FLIP_FLOP_D \registres_reg[12][1]  ( .D(n5368), .CK(clock), .Q(
        \registres[12][1] ) );
  FLIP_FLOP_D \registres_reg[12][0]  ( .D(n5367), .CK(clock), .Q(
        \registres[12][0] ) );
  FLIP_FLOP_D \registres_reg[13][31]  ( .D(n5366), .CK(clock), .Q(
        \registres[13][31] ) );
  FLIP_FLOP_D \registres_reg[13][30]  ( .D(n5365), .CK(clock), .Q(
        \registres[13][30] ) );
  FLIP_FLOP_D \registres_reg[13][29]  ( .D(n5364), .CK(clock), .Q(
        \registres[13][29] ) );
  FLIP_FLOP_D \registres_reg[13][28]  ( .D(n5363), .CK(clock), .Q(
        \registres[13][28] ) );
  FLIP_FLOP_D \registres_reg[13][27]  ( .D(n5362), .CK(clock), .Q(
        \registres[13][27] ) );
  FLIP_FLOP_D \registres_reg[13][26]  ( .D(n5361), .CK(clock), .Q(
        \registres[13][26] ) );
  FLIP_FLOP_D \registres_reg[13][25]  ( .D(n5360), .CK(clock), .Q(
        \registres[13][25] ) );
  FLIP_FLOP_D \registres_reg[13][24]  ( .D(n5359), .CK(clock), .Q(
        \registres[13][24] ) );
  FLIP_FLOP_D \registres_reg[13][23]  ( .D(n5358), .CK(clock), .Q(
        \registres[13][23] ) );
  FLIP_FLOP_D \registres_reg[13][22]  ( .D(n5357), .CK(clock), .Q(
        \registres[13][22] ) );
  FLIP_FLOP_D \registres_reg[13][21]  ( .D(n5356), .CK(clock), .Q(
        \registres[13][21] ) );
  FLIP_FLOP_D \registres_reg[13][20]  ( .D(n5355), .CK(clock), .Q(
        \registres[13][20] ) );
  FLIP_FLOP_D \registres_reg[13][19]  ( .D(n5354), .CK(clock), .Q(
        \registres[13][19] ) );
  FLIP_FLOP_D \registres_reg[13][18]  ( .D(n5353), .CK(clock), .Q(
        \registres[13][18] ) );
  FLIP_FLOP_D \registres_reg[13][17]  ( .D(n5352), .CK(clock), .Q(
        \registres[13][17] ) );
  FLIP_FLOP_D \registres_reg[13][16]  ( .D(n5351), .CK(clock), .Q(
        \registres[13][16] ) );
  FLIP_FLOP_D \registres_reg[13][15]  ( .D(n5350), .CK(clock), .Q(
        \registres[13][15] ) );
  FLIP_FLOP_D \registres_reg[13][14]  ( .D(n5349), .CK(clock), .Q(
        \registres[13][14] ) );
  FLIP_FLOP_D \registres_reg[13][13]  ( .D(n5348), .CK(clock), .Q(
        \registres[13][13] ) );
  FLIP_FLOP_D \registres_reg[13][12]  ( .D(n5347), .CK(clock), .Q(
        \registres[13][12] ) );
  FLIP_FLOP_D \registres_reg[13][11]  ( .D(n5346), .CK(clock), .Q(
        \registres[13][11] ) );
  FLIP_FLOP_D \registres_reg[13][10]  ( .D(n5345), .CK(clock), .Q(
        \registres[13][10] ) );
  FLIP_FLOP_D \registres_reg[13][9]  ( .D(n5344), .CK(clock), .Q(
        \registres[13][9] ) );
  FLIP_FLOP_D \registres_reg[13][8]  ( .D(n5343), .CK(clock), .Q(
        \registres[13][8] ) );
  FLIP_FLOP_D \registres_reg[13][7]  ( .D(n5342), .CK(clock), .Q(
        \registres[13][7] ) );
  FLIP_FLOP_D \registres_reg[13][6]  ( .D(n5341), .CK(clock), .Q(
        \registres[13][6] ) );
  FLIP_FLOP_D \registres_reg[13][5]  ( .D(n5340), .CK(clock), .Q(
        \registres[13][5] ) );
  FLIP_FLOP_D \registres_reg[13][4]  ( .D(n5339), .CK(clock), .Q(
        \registres[13][4] ) );
  FLIP_FLOP_D \registres_reg[13][3]  ( .D(n5338), .CK(clock), .Q(
        \registres[13][3] ) );
  FLIP_FLOP_D \registres_reg[13][2]  ( .D(n5337), .CK(clock), .Q(
        \registres[13][2] ) );
  FLIP_FLOP_D \registres_reg[13][1]  ( .D(n5336), .CK(clock), .Q(
        \registres[13][1] ) );
  FLIP_FLOP_D \registres_reg[13][0]  ( .D(n5335), .CK(clock), .Q(
        \registres[13][0] ) );
  FLIP_FLOP_D \registres_reg[14][31]  ( .D(n5334), .CK(clock), .Q(
        \registres[14][31] ) );
  FLIP_FLOP_D \registres_reg[14][30]  ( .D(n5333), .CK(clock), .Q(
        \registres[14][30] ) );
  FLIP_FLOP_D \registres_reg[14][29]  ( .D(n5332), .CK(clock), .Q(
        \registres[14][29] ) );
  FLIP_FLOP_D \registres_reg[14][28]  ( .D(n5331), .CK(clock), .Q(
        \registres[14][28] ) );
  FLIP_FLOP_D \registres_reg[14][27]  ( .D(n5330), .CK(clock), .Q(
        \registres[14][27] ) );
  FLIP_FLOP_D \registres_reg[14][26]  ( .D(n5329), .CK(clock), .Q(
        \registres[14][26] ) );
  FLIP_FLOP_D \registres_reg[14][25]  ( .D(n5328), .CK(clock), .Q(
        \registres[14][25] ) );
  FLIP_FLOP_D \registres_reg[14][24]  ( .D(n5327), .CK(clock), .Q(
        \registres[14][24] ) );
  FLIP_FLOP_D \registres_reg[14][23]  ( .D(n5326), .CK(clock), .Q(
        \registres[14][23] ) );
  FLIP_FLOP_D \registres_reg[14][22]  ( .D(n5325), .CK(clock), .Q(
        \registres[14][22] ) );
  FLIP_FLOP_D \registres_reg[14][21]  ( .D(n5324), .CK(clock), .Q(
        \registres[14][21] ) );
  FLIP_FLOP_D \registres_reg[14][20]  ( .D(n5323), .CK(clock), .Q(
        \registres[14][20] ) );
  FLIP_FLOP_D \registres_reg[14][19]  ( .D(n5322), .CK(clock), .Q(
        \registres[14][19] ) );
  FLIP_FLOP_D \registres_reg[14][18]  ( .D(n5321), .CK(clock), .Q(
        \registres[14][18] ) );
  FLIP_FLOP_D \registres_reg[14][17]  ( .D(n5320), .CK(clock), .Q(
        \registres[14][17] ) );
  FLIP_FLOP_D \registres_reg[14][16]  ( .D(n5319), .CK(clock), .Q(
        \registres[14][16] ) );
  FLIP_FLOP_D \registres_reg[14][15]  ( .D(n5318), .CK(clock), .Q(
        \registres[14][15] ) );
  FLIP_FLOP_D \registres_reg[14][14]  ( .D(n5317), .CK(clock), .Q(
        \registres[14][14] ) );
  FLIP_FLOP_D \registres_reg[14][13]  ( .D(n5316), .CK(clock), .Q(
        \registres[14][13] ) );
  FLIP_FLOP_D \registres_reg[14][12]  ( .D(n5315), .CK(clock), .Q(
        \registres[14][12] ) );
  FLIP_FLOP_D \registres_reg[14][11]  ( .D(n5314), .CK(clock), .Q(
        \registres[14][11] ) );
  FLIP_FLOP_D \registres_reg[14][10]  ( .D(n5313), .CK(clock), .Q(
        \registres[14][10] ) );
  FLIP_FLOP_D \registres_reg[14][9]  ( .D(n5312), .CK(clock), .Q(
        \registres[14][9] ) );
  FLIP_FLOP_D \registres_reg[14][8]  ( .D(n5311), .CK(clock), .Q(
        \registres[14][8] ) );
  FLIP_FLOP_D \registres_reg[14][7]  ( .D(n5310), .CK(clock), .Q(
        \registres[14][7] ) );
  FLIP_FLOP_D \registres_reg[14][6]  ( .D(n5309), .CK(clock), .Q(
        \registres[14][6] ) );
  FLIP_FLOP_D \registres_reg[14][5]  ( .D(n5308), .CK(clock), .Q(
        \registres[14][5] ) );
  FLIP_FLOP_D \registres_reg[14][4]  ( .D(n5307), .CK(clock), .Q(
        \registres[14][4] ) );
  FLIP_FLOP_D \registres_reg[14][3]  ( .D(n5306), .CK(clock), .Q(
        \registres[14][3] ) );
  FLIP_FLOP_D \registres_reg[14][2]  ( .D(n5305), .CK(clock), .Q(
        \registres[14][2] ) );
  FLIP_FLOP_D \registres_reg[14][1]  ( .D(n5304), .CK(clock), .Q(
        \registres[14][1] ) );
  FLIP_FLOP_D \registres_reg[14][0]  ( .D(n5303), .CK(clock), .Q(
        \registres[14][0] ) );
  FLIP_FLOP_D \registres_reg[15][31]  ( .D(n5302), .CK(clock), .Q(
        \registres[15][31] ) );
  FLIP_FLOP_D \registres_reg[15][30]  ( .D(n5301), .CK(clock), .Q(
        \registres[15][30] ) );
  FLIP_FLOP_D \registres_reg[15][29]  ( .D(n5300), .CK(clock), .Q(
        \registres[15][29] ) );
  FLIP_FLOP_D \registres_reg[15][28]  ( .D(n5299), .CK(clock), .Q(
        \registres[15][28] ) );
  FLIP_FLOP_D \registres_reg[15][27]  ( .D(n5298), .CK(clock), .Q(
        \registres[15][27] ) );
  FLIP_FLOP_D \registres_reg[15][26]  ( .D(n5297), .CK(clock), .Q(
        \registres[15][26] ) );
  FLIP_FLOP_D \registres_reg[15][25]  ( .D(n5296), .CK(clock), .Q(
        \registres[15][25] ) );
  FLIP_FLOP_D \registres_reg[15][24]  ( .D(n5295), .CK(clock), .Q(
        \registres[15][24] ) );
  FLIP_FLOP_D \registres_reg[15][23]  ( .D(n5294), .CK(clock), .Q(
        \registres[15][23] ) );
  FLIP_FLOP_D \registres_reg[15][22]  ( .D(n5293), .CK(clock), .Q(
        \registres[15][22] ) );
  FLIP_FLOP_D \registres_reg[15][21]  ( .D(n5292), .CK(clock), .Q(
        \registres[15][21] ) );
  FLIP_FLOP_D \registres_reg[15][20]  ( .D(n5291), .CK(clock), .Q(
        \registres[15][20] ) );
  FLIP_FLOP_D \registres_reg[15][19]  ( .D(n5290), .CK(clock), .Q(
        \registres[15][19] ) );
  FLIP_FLOP_D \registres_reg[15][18]  ( .D(n5289), .CK(clock), .Q(
        \registres[15][18] ) );
  FLIP_FLOP_D \registres_reg[15][17]  ( .D(n5288), .CK(clock), .Q(
        \registres[15][17] ) );
  FLIP_FLOP_D \registres_reg[15][16]  ( .D(n5287), .CK(clock), .Q(
        \registres[15][16] ) );
  FLIP_FLOP_D \registres_reg[15][15]  ( .D(n5286), .CK(clock), .Q(
        \registres[15][15] ) );
  FLIP_FLOP_D \registres_reg[15][14]  ( .D(n5285), .CK(clock), .Q(
        \registres[15][14] ) );
  FLIP_FLOP_D \registres_reg[15][13]  ( .D(n5284), .CK(clock), .Q(
        \registres[15][13] ) );
  FLIP_FLOP_D \registres_reg[15][12]  ( .D(n5283), .CK(clock), .Q(
        \registres[15][12] ) );
  FLIP_FLOP_D \registres_reg[15][11]  ( .D(n5282), .CK(clock), .Q(
        \registres[15][11] ) );
  FLIP_FLOP_D \registres_reg[15][10]  ( .D(n5281), .CK(clock), .Q(
        \registres[15][10] ) );
  FLIP_FLOP_D \registres_reg[15][9]  ( .D(n5280), .CK(clock), .Q(
        \registres[15][9] ) );
  FLIP_FLOP_D \registres_reg[15][8]  ( .D(n5279), .CK(clock), .Q(
        \registres[15][8] ) );
  FLIP_FLOP_D \registres_reg[15][7]  ( .D(n5278), .CK(clock), .Q(
        \registres[15][7] ) );
  FLIP_FLOP_D \registres_reg[15][6]  ( .D(n5277), .CK(clock), .Q(
        \registres[15][6] ) );
  FLIP_FLOP_D \registres_reg[15][5]  ( .D(n5276), .CK(clock), .Q(
        \registres[15][5] ) );
  FLIP_FLOP_D \registres_reg[15][4]  ( .D(n5275), .CK(clock), .Q(
        \registres[15][4] ) );
  FLIP_FLOP_D \registres_reg[15][3]  ( .D(n5274), .CK(clock), .Q(
        \registres[15][3] ) );
  FLIP_FLOP_D \registres_reg[15][2]  ( .D(n5273), .CK(clock), .Q(
        \registres[15][2] ) );
  FLIP_FLOP_D \registres_reg[15][1]  ( .D(n5272), .CK(clock), .Q(
        \registres[15][1] ) );
  FLIP_FLOP_D \registres_reg[15][0]  ( .D(n5271), .CK(clock), .Q(
        \registres[15][0] ) );
  FLIP_FLOP_D \registres_reg[16][31]  ( .D(n5270), .CK(clock), .Q(
        \registres[16][31] ) );
  FLIP_FLOP_D \registres_reg[16][30]  ( .D(n5269), .CK(clock), .Q(
        \registres[16][30] ) );
  FLIP_FLOP_D \registres_reg[16][29]  ( .D(n5268), .CK(clock), .Q(
        \registres[16][29] ) );
  FLIP_FLOP_D \registres_reg[16][28]  ( .D(n5267), .CK(clock), .Q(
        \registres[16][28] ) );
  FLIP_FLOP_D \registres_reg[16][27]  ( .D(n5266), .CK(clock), .Q(
        \registres[16][27] ) );
  FLIP_FLOP_D \registres_reg[16][26]  ( .D(n5265), .CK(clock), .Q(
        \registres[16][26] ) );
  FLIP_FLOP_D \registres_reg[16][25]  ( .D(n5264), .CK(clock), .Q(
        \registres[16][25] ) );
  FLIP_FLOP_D \registres_reg[16][24]  ( .D(n5263), .CK(clock), .Q(
        \registres[16][24] ) );
  FLIP_FLOP_D \registres_reg[16][23]  ( .D(n5262), .CK(clock), .Q(
        \registres[16][23] ) );
  FLIP_FLOP_D \registres_reg[16][22]  ( .D(n5261), .CK(clock), .Q(
        \registres[16][22] ) );
  FLIP_FLOP_D \registres_reg[16][21]  ( .D(n5260), .CK(clock), .Q(
        \registres[16][21] ) );
  FLIP_FLOP_D \registres_reg[16][20]  ( .D(n5259), .CK(clock), .Q(
        \registres[16][20] ) );
  FLIP_FLOP_D \registres_reg[16][19]  ( .D(n5258), .CK(clock), .Q(
        \registres[16][19] ) );
  FLIP_FLOP_D \registres_reg[16][18]  ( .D(n5257), .CK(clock), .Q(
        \registres[16][18] ) );
  FLIP_FLOP_D \registres_reg[16][17]  ( .D(n5256), .CK(clock), .Q(
        \registres[16][17] ) );
  FLIP_FLOP_D \registres_reg[16][16]  ( .D(n5255), .CK(clock), .Q(
        \registres[16][16] ) );
  FLIP_FLOP_D \registres_reg[16][15]  ( .D(n5254), .CK(clock), .Q(
        \registres[16][15] ) );
  FLIP_FLOP_D \registres_reg[16][14]  ( .D(n5253), .CK(clock), .Q(
        \registres[16][14] ) );
  FLIP_FLOP_D \registres_reg[16][13]  ( .D(n5252), .CK(clock), .Q(
        \registres[16][13] ) );
  FLIP_FLOP_D \registres_reg[16][12]  ( .D(n5251), .CK(clock), .Q(
        \registres[16][12] ) );
  FLIP_FLOP_D \registres_reg[16][11]  ( .D(n5250), .CK(clock), .Q(
        \registres[16][11] ) );
  FLIP_FLOP_D \registres_reg[16][10]  ( .D(n5249), .CK(clock), .Q(
        \registres[16][10] ) );
  FLIP_FLOP_D \registres_reg[16][9]  ( .D(n5248), .CK(clock), .Q(
        \registres[16][9] ) );
  FLIP_FLOP_D \registres_reg[16][8]  ( .D(n5247), .CK(clock), .Q(
        \registres[16][8] ) );
  FLIP_FLOP_D \registres_reg[16][7]  ( .D(n5246), .CK(clock), .Q(
        \registres[16][7] ) );
  FLIP_FLOP_D \registres_reg[16][6]  ( .D(n5245), .CK(clock), .Q(
        \registres[16][6] ) );
  FLIP_FLOP_D \registres_reg[16][5]  ( .D(n5244), .CK(clock), .Q(
        \registres[16][5] ) );
  FLIP_FLOP_D \registres_reg[16][4]  ( .D(n5243), .CK(clock), .Q(
        \registres[16][4] ) );
  FLIP_FLOP_D \registres_reg[16][3]  ( .D(n5242), .CK(clock), .Q(
        \registres[16][3] ) );
  FLIP_FLOP_D \registres_reg[16][2]  ( .D(n5241), .CK(clock), .Q(
        \registres[16][2] ) );
  FLIP_FLOP_D \registres_reg[16][1]  ( .D(n5240), .CK(clock), .Q(
        \registres[16][1] ) );
  FLIP_FLOP_D \registres_reg[16][0]  ( .D(n5239), .CK(clock), .Q(
        \registres[16][0] ) );
  FLIP_FLOP_D \registres_reg[17][31]  ( .D(n5238), .CK(clock), .Q(
        \registres[17][31] ) );
  FLIP_FLOP_D \registres_reg[17][30]  ( .D(n5237), .CK(clock), .Q(
        \registres[17][30] ) );
  FLIP_FLOP_D \registres_reg[17][29]  ( .D(n5236), .CK(clock), .Q(
        \registres[17][29] ) );
  FLIP_FLOP_D \registres_reg[17][28]  ( .D(n5235), .CK(clock), .Q(
        \registres[17][28] ) );
  FLIP_FLOP_D \registres_reg[17][27]  ( .D(n5234), .CK(clock), .Q(
        \registres[17][27] ) );
  FLIP_FLOP_D \registres_reg[17][26]  ( .D(n5233), .CK(clock), .Q(
        \registres[17][26] ) );
  FLIP_FLOP_D \registres_reg[17][25]  ( .D(n5232), .CK(clock), .Q(
        \registres[17][25] ) );
  FLIP_FLOP_D \registres_reg[17][24]  ( .D(n5231), .CK(clock), .Q(
        \registres[17][24] ) );
  FLIP_FLOP_D \registres_reg[17][23]  ( .D(n5230), .CK(clock), .Q(
        \registres[17][23] ) );
  FLIP_FLOP_D \registres_reg[17][22]  ( .D(n5229), .CK(clock), .Q(
        \registres[17][22] ) );
  FLIP_FLOP_D \registres_reg[17][21]  ( .D(n5228), .CK(clock), .Q(
        \registres[17][21] ) );
  FLIP_FLOP_D \registres_reg[17][20]  ( .D(n5227), .CK(clock), .Q(
        \registres[17][20] ) );
  FLIP_FLOP_D \registres_reg[17][19]  ( .D(n5226), .CK(clock), .Q(
        \registres[17][19] ) );
  FLIP_FLOP_D \registres_reg[17][18]  ( .D(n5225), .CK(clock), .Q(
        \registres[17][18] ) );
  FLIP_FLOP_D \registres_reg[17][17]  ( .D(n5224), .CK(clock), .Q(
        \registres[17][17] ) );
  FLIP_FLOP_D \registres_reg[17][16]  ( .D(n5223), .CK(clock), .Q(
        \registres[17][16] ) );
  FLIP_FLOP_D \registres_reg[17][15]  ( .D(n5222), .CK(clock), .Q(
        \registres[17][15] ) );
  FLIP_FLOP_D \registres_reg[17][14]  ( .D(n5221), .CK(clock), .Q(
        \registres[17][14] ) );
  FLIP_FLOP_D \registres_reg[17][13]  ( .D(n5220), .CK(clock), .Q(
        \registres[17][13] ) );
  FLIP_FLOP_D \registres_reg[17][12]  ( .D(n5219), .CK(clock), .Q(
        \registres[17][12] ) );
  FLIP_FLOP_D \registres_reg[17][11]  ( .D(n5218), .CK(clock), .Q(
        \registres[17][11] ) );
  FLIP_FLOP_D \registres_reg[17][10]  ( .D(n5217), .CK(clock), .Q(
        \registres[17][10] ) );
  FLIP_FLOP_D \registres_reg[17][9]  ( .D(n5216), .CK(clock), .Q(
        \registres[17][9] ) );
  FLIP_FLOP_D \registres_reg[17][8]  ( .D(n5215), .CK(clock), .Q(
        \registres[17][8] ) );
  FLIP_FLOP_D \registres_reg[17][7]  ( .D(n5214), .CK(clock), .Q(
        \registres[17][7] ) );
  FLIP_FLOP_D \registres_reg[17][6]  ( .D(n5213), .CK(clock), .Q(
        \registres[17][6] ) );
  FLIP_FLOP_D \registres_reg[17][5]  ( .D(n5212), .CK(clock), .Q(
        \registres[17][5] ) );
  FLIP_FLOP_D \registres_reg[17][4]  ( .D(n5211), .CK(clock), .Q(
        \registres[17][4] ) );
  FLIP_FLOP_D \registres_reg[17][3]  ( .D(n5210), .CK(clock), .Q(
        \registres[17][3] ) );
  FLIP_FLOP_D \registres_reg[17][2]  ( .D(n5209), .CK(clock), .Q(
        \registres[17][2] ) );
  FLIP_FLOP_D \registres_reg[17][1]  ( .D(n5208), .CK(clock), .Q(
        \registres[17][1] ) );
  FLIP_FLOP_D \registres_reg[17][0]  ( .D(n5207), .CK(clock), .Q(
        \registres[17][0] ) );
  FLIP_FLOP_D \registres_reg[18][31]  ( .D(n5206), .CK(clock), .Q(
        \registres[18][31] ) );
  FLIP_FLOP_D \registres_reg[18][30]  ( .D(n5205), .CK(clock), .Q(
        \registres[18][30] ) );
  FLIP_FLOP_D \registres_reg[18][29]  ( .D(n5204), .CK(clock), .Q(
        \registres[18][29] ) );
  FLIP_FLOP_D \registres_reg[18][28]  ( .D(n5203), .CK(clock), .Q(
        \registres[18][28] ) );
  FLIP_FLOP_D \registres_reg[18][27]  ( .D(n5202), .CK(clock), .Q(
        \registres[18][27] ) );
  FLIP_FLOP_D \registres_reg[18][26]  ( .D(n5201), .CK(clock), .Q(
        \registres[18][26] ) );
  FLIP_FLOP_D \registres_reg[18][25]  ( .D(n5200), .CK(clock), .Q(
        \registres[18][25] ) );
  FLIP_FLOP_D \registres_reg[18][24]  ( .D(n5199), .CK(clock), .Q(
        \registres[18][24] ) );
  FLIP_FLOP_D \registres_reg[18][23]  ( .D(n5198), .CK(clock), .Q(
        \registres[18][23] ) );
  FLIP_FLOP_D \registres_reg[18][22]  ( .D(n5197), .CK(clock), .Q(
        \registres[18][22] ) );
  FLIP_FLOP_D \registres_reg[18][21]  ( .D(n5196), .CK(clock), .Q(
        \registres[18][21] ) );
  FLIP_FLOP_D \registres_reg[18][20]  ( .D(n5195), .CK(clock), .Q(
        \registres[18][20] ) );
  FLIP_FLOP_D \registres_reg[18][19]  ( .D(n5194), .CK(clock), .Q(
        \registres[18][19] ) );
  FLIP_FLOP_D \registres_reg[18][18]  ( .D(n5193), .CK(clock), .Q(
        \registres[18][18] ) );
  FLIP_FLOP_D \registres_reg[18][17]  ( .D(n5192), .CK(clock), .Q(
        \registres[18][17] ) );
  FLIP_FLOP_D \registres_reg[18][16]  ( .D(n5191), .CK(clock), .Q(
        \registres[18][16] ) );
  FLIP_FLOP_D \registres_reg[18][15]  ( .D(n5190), .CK(clock), .Q(
        \registres[18][15] ) );
  FLIP_FLOP_D \registres_reg[18][14]  ( .D(n5189), .CK(clock), .Q(
        \registres[18][14] ) );
  FLIP_FLOP_D \registres_reg[18][13]  ( .D(n5188), .CK(clock), .Q(
        \registres[18][13] ) );
  FLIP_FLOP_D \registres_reg[18][12]  ( .D(n5187), .CK(clock), .Q(
        \registres[18][12] ) );
  FLIP_FLOP_D \registres_reg[18][11]  ( .D(n5186), .CK(clock), .Q(
        \registres[18][11] ) );
  FLIP_FLOP_D \registres_reg[18][10]  ( .D(n5185), .CK(clock), .Q(
        \registres[18][10] ) );
  FLIP_FLOP_D \registres_reg[18][9]  ( .D(n5184), .CK(clock), .Q(
        \registres[18][9] ) );
  FLIP_FLOP_D \registres_reg[18][8]  ( .D(n5183), .CK(clock), .Q(
        \registres[18][8] ) );
  FLIP_FLOP_D \registres_reg[18][7]  ( .D(n5182), .CK(clock), .Q(
        \registres[18][7] ) );
  FLIP_FLOP_D \registres_reg[18][6]  ( .D(n5181), .CK(clock), .Q(
        \registres[18][6] ) );
  FLIP_FLOP_D \registres_reg[18][5]  ( .D(n5180), .CK(clock), .Q(
        \registres[18][5] ) );
  FLIP_FLOP_D \registres_reg[18][4]  ( .D(n5179), .CK(clock), .Q(
        \registres[18][4] ) );
  FLIP_FLOP_D \registres_reg[18][3]  ( .D(n5178), .CK(clock), .Q(
        \registres[18][3] ) );
  FLIP_FLOP_D \registres_reg[18][2]  ( .D(n5177), .CK(clock), .Q(
        \registres[18][2] ) );
  FLIP_FLOP_D \registres_reg[18][1]  ( .D(n5176), .CK(clock), .Q(
        \registres[18][1] ) );
  FLIP_FLOP_D \registres_reg[18][0]  ( .D(n5175), .CK(clock), .Q(
        \registres[18][0] ) );
  FLIP_FLOP_D \registres_reg[19][31]  ( .D(n5174), .CK(clock), .Q(
        \registres[19][31] ) );
  FLIP_FLOP_D \registres_reg[19][30]  ( .D(n5173), .CK(clock), .Q(
        \registres[19][30] ) );
  FLIP_FLOP_D \registres_reg[19][29]  ( .D(n5172), .CK(clock), .Q(
        \registres[19][29] ) );
  FLIP_FLOP_D \registres_reg[19][28]  ( .D(n5171), .CK(clock), .Q(
        \registres[19][28] ) );
  FLIP_FLOP_D \registres_reg[19][27]  ( .D(n5170), .CK(clock), .Q(
        \registres[19][27] ) );
  FLIP_FLOP_D \registres_reg[19][26]  ( .D(n5169), .CK(clock), .Q(
        \registres[19][26] ) );
  FLIP_FLOP_D \registres_reg[19][25]  ( .D(n5168), .CK(clock), .Q(
        \registres[19][25] ) );
  FLIP_FLOP_D \registres_reg[19][24]  ( .D(n5167), .CK(clock), .Q(
        \registres[19][24] ) );
  FLIP_FLOP_D \registres_reg[19][23]  ( .D(n5166), .CK(clock), .Q(
        \registres[19][23] ) );
  FLIP_FLOP_D \registres_reg[19][22]  ( .D(n5165), .CK(clock), .Q(
        \registres[19][22] ) );
  FLIP_FLOP_D \registres_reg[19][21]  ( .D(n5164), .CK(clock), .Q(
        \registres[19][21] ) );
  FLIP_FLOP_D \registres_reg[19][20]  ( .D(n5163), .CK(clock), .Q(
        \registres[19][20] ) );
  FLIP_FLOP_D \registres_reg[19][19]  ( .D(n5162), .CK(clock), .Q(
        \registres[19][19] ) );
  FLIP_FLOP_D \registres_reg[19][18]  ( .D(n5161), .CK(clock), .Q(
        \registres[19][18] ) );
  FLIP_FLOP_D \registres_reg[19][17]  ( .D(n5160), .CK(clock), .Q(
        \registres[19][17] ) );
  FLIP_FLOP_D \registres_reg[19][16]  ( .D(n5159), .CK(clock), .Q(
        \registres[19][16] ) );
  FLIP_FLOP_D \registres_reg[19][15]  ( .D(n5158), .CK(clock), .Q(
        \registres[19][15] ) );
  FLIP_FLOP_D \registres_reg[19][14]  ( .D(n5157), .CK(clock), .Q(
        \registres[19][14] ) );
  FLIP_FLOP_D \registres_reg[19][13]  ( .D(n5156), .CK(clock), .Q(
        \registres[19][13] ) );
  FLIP_FLOP_D \registres_reg[19][12]  ( .D(n5155), .CK(clock), .Q(
        \registres[19][12] ) );
  FLIP_FLOP_D \registres_reg[19][11]  ( .D(n5154), .CK(clock), .Q(
        \registres[19][11] ) );
  FLIP_FLOP_D \registres_reg[19][10]  ( .D(n5153), .CK(clock), .Q(
        \registres[19][10] ) );
  FLIP_FLOP_D \registres_reg[19][9]  ( .D(n5152), .CK(clock), .Q(
        \registres[19][9] ) );
  FLIP_FLOP_D \registres_reg[19][8]  ( .D(n5151), .CK(clock), .Q(
        \registres[19][8] ) );
  FLIP_FLOP_D \registres_reg[19][7]  ( .D(n5150), .CK(clock), .Q(
        \registres[19][7] ) );
  FLIP_FLOP_D \registres_reg[19][6]  ( .D(n5149), .CK(clock), .Q(
        \registres[19][6] ) );
  FLIP_FLOP_D \registres_reg[19][5]  ( .D(n5148), .CK(clock), .Q(
        \registres[19][5] ) );
  FLIP_FLOP_D \registres_reg[19][4]  ( .D(n5147), .CK(clock), .Q(
        \registres[19][4] ) );
  FLIP_FLOP_D \registres_reg[19][3]  ( .D(n5146), .CK(clock), .Q(
        \registres[19][3] ) );
  FLIP_FLOP_D \registres_reg[19][2]  ( .D(n5145), .CK(clock), .Q(
        \registres[19][2] ) );
  FLIP_FLOP_D \registres_reg[19][1]  ( .D(n5144), .CK(clock), .Q(
        \registres[19][1] ) );
  FLIP_FLOP_D \registres_reg[19][0]  ( .D(n5143), .CK(clock), .Q(
        \registres[19][0] ) );
  FLIP_FLOP_D \registres_reg[20][31]  ( .D(n5142), .CK(clock), .Q(
        \registres[20][31] ) );
  FLIP_FLOP_D \registres_reg[20][30]  ( .D(n5141), .CK(clock), .Q(
        \registres[20][30] ) );
  FLIP_FLOP_D \registres_reg[20][29]  ( .D(n5140), .CK(clock), .Q(
        \registres[20][29] ) );
  FLIP_FLOP_D \registres_reg[20][28]  ( .D(n5139), .CK(clock), .Q(
        \registres[20][28] ) );
  FLIP_FLOP_D \registres_reg[20][27]  ( .D(n5138), .CK(clock), .Q(
        \registres[20][27] ) );
  FLIP_FLOP_D \registres_reg[20][26]  ( .D(n5137), .CK(clock), .Q(
        \registres[20][26] ) );
  FLIP_FLOP_D \registres_reg[20][25]  ( .D(n5136), .CK(clock), .Q(
        \registres[20][25] ) );
  FLIP_FLOP_D \registres_reg[20][24]  ( .D(n5135), .CK(clock), .Q(
        \registres[20][24] ) );
  FLIP_FLOP_D \registres_reg[20][23]  ( .D(n5134), .CK(clock), .Q(
        \registres[20][23] ) );
  FLIP_FLOP_D \registres_reg[20][22]  ( .D(n5133), .CK(clock), .Q(
        \registres[20][22] ) );
  FLIP_FLOP_D \registres_reg[20][21]  ( .D(n5132), .CK(clock), .Q(
        \registres[20][21] ) );
  FLIP_FLOP_D \registres_reg[20][20]  ( .D(n5131), .CK(clock), .Q(
        \registres[20][20] ) );
  FLIP_FLOP_D \registres_reg[20][19]  ( .D(n5130), .CK(clock), .Q(
        \registres[20][19] ) );
  FLIP_FLOP_D \registres_reg[20][18]  ( .D(n5129), .CK(clock), .Q(
        \registres[20][18] ) );
  FLIP_FLOP_D \registres_reg[20][17]  ( .D(n5128), .CK(clock), .Q(
        \registres[20][17] ) );
  FLIP_FLOP_D \registres_reg[20][16]  ( .D(n5127), .CK(clock), .Q(
        \registres[20][16] ) );
  FLIP_FLOP_D \registres_reg[20][15]  ( .D(n5126), .CK(clock), .Q(
        \registres[20][15] ) );
  FLIP_FLOP_D \registres_reg[20][14]  ( .D(n5125), .CK(clock), .Q(
        \registres[20][14] ) );
  FLIP_FLOP_D \registres_reg[20][13]  ( .D(n5124), .CK(clock), .Q(
        \registres[20][13] ) );
  FLIP_FLOP_D \registres_reg[20][12]  ( .D(n5123), .CK(clock), .Q(
        \registres[20][12] ) );
  FLIP_FLOP_D \registres_reg[20][11]  ( .D(n5122), .CK(clock), .Q(
        \registres[20][11] ) );
  FLIP_FLOP_D \registres_reg[20][10]  ( .D(n5121), .CK(clock), .Q(
        \registres[20][10] ) );
  FLIP_FLOP_D \registres_reg[20][9]  ( .D(n5120), .CK(clock), .Q(
        \registres[20][9] ) );
  FLIP_FLOP_D \registres_reg[20][8]  ( .D(n5119), .CK(clock), .Q(
        \registres[20][8] ) );
  FLIP_FLOP_D \registres_reg[20][7]  ( .D(n5118), .CK(clock), .Q(
        \registres[20][7] ) );
  FLIP_FLOP_D \registres_reg[20][6]  ( .D(n5117), .CK(clock), .Q(
        \registres[20][6] ) );
  FLIP_FLOP_D \registres_reg[20][5]  ( .D(n5116), .CK(clock), .Q(
        \registres[20][5] ) );
  FLIP_FLOP_D \registres_reg[20][4]  ( .D(n5115), .CK(clock), .Q(
        \registres[20][4] ) );
  FLIP_FLOP_D \registres_reg[20][3]  ( .D(n5114), .CK(clock), .Q(
        \registres[20][3] ) );
  FLIP_FLOP_D \registres_reg[20][2]  ( .D(n5113), .CK(clock), .Q(
        \registres[20][2] ) );
  FLIP_FLOP_D \registres_reg[20][1]  ( .D(n5112), .CK(clock), .Q(
        \registres[20][1] ) );
  FLIP_FLOP_D \registres_reg[20][0]  ( .D(n5111), .CK(clock), .Q(
        \registres[20][0] ) );
  FLIP_FLOP_D \registres_reg[21][31]  ( .D(n5110), .CK(clock), .Q(
        \registres[21][31] ) );
  FLIP_FLOP_D \registres_reg[21][30]  ( .D(n5109), .CK(clock), .Q(
        \registres[21][30] ) );
  FLIP_FLOP_D \registres_reg[21][29]  ( .D(n5108), .CK(clock), .Q(
        \registres[21][29] ) );
  FLIP_FLOP_D \registres_reg[21][28]  ( .D(n5107), .CK(clock), .Q(
        \registres[21][28] ) );
  FLIP_FLOP_D \registres_reg[21][27]  ( .D(n5106), .CK(clock), .Q(
        \registres[21][27] ) );
  FLIP_FLOP_D \registres_reg[21][26]  ( .D(n5105), .CK(clock), .Q(
        \registres[21][26] ) );
  FLIP_FLOP_D \registres_reg[21][25]  ( .D(n5104), .CK(clock), .Q(
        \registres[21][25] ) );
  FLIP_FLOP_D \registres_reg[21][24]  ( .D(n5103), .CK(clock), .Q(
        \registres[21][24] ) );
  FLIP_FLOP_D \registres_reg[21][23]  ( .D(n5102), .CK(clock), .Q(
        \registres[21][23] ) );
  FLIP_FLOP_D \registres_reg[21][22]  ( .D(n5101), .CK(clock), .Q(
        \registres[21][22] ) );
  FLIP_FLOP_D \registres_reg[21][21]  ( .D(n5100), .CK(clock), .Q(
        \registres[21][21] ) );
  FLIP_FLOP_D \registres_reg[21][20]  ( .D(n5099), .CK(clock), .Q(
        \registres[21][20] ) );
  FLIP_FLOP_D \registres_reg[21][19]  ( .D(n5098), .CK(clock), .Q(
        \registres[21][19] ) );
  FLIP_FLOP_D \registres_reg[21][18]  ( .D(n5097), .CK(clock), .Q(
        \registres[21][18] ) );
  FLIP_FLOP_D \registres_reg[21][17]  ( .D(n5096), .CK(clock), .Q(
        \registres[21][17] ) );
  FLIP_FLOP_D \registres_reg[21][16]  ( .D(n5095), .CK(clock), .Q(
        \registres[21][16] ) );
  FLIP_FLOP_D \registres_reg[21][15]  ( .D(n5094), .CK(clock), .Q(
        \registres[21][15] ) );
  FLIP_FLOP_D \registres_reg[21][14]  ( .D(n5093), .CK(clock), .Q(
        \registres[21][14] ) );
  FLIP_FLOP_D \registres_reg[21][13]  ( .D(n5092), .CK(clock), .Q(
        \registres[21][13] ) );
  FLIP_FLOP_D \registres_reg[21][12]  ( .D(n5091), .CK(clock), .Q(
        \registres[21][12] ) );
  FLIP_FLOP_D \registres_reg[21][11]  ( .D(n5090), .CK(clock), .Q(
        \registres[21][11] ) );
  FLIP_FLOP_D \registres_reg[21][10]  ( .D(n5089), .CK(clock), .Q(
        \registres[21][10] ) );
  FLIP_FLOP_D \registres_reg[21][9]  ( .D(n5088), .CK(clock), .Q(
        \registres[21][9] ) );
  FLIP_FLOP_D \registres_reg[21][8]  ( .D(n5087), .CK(clock), .Q(
        \registres[21][8] ) );
  FLIP_FLOP_D \registres_reg[21][7]  ( .D(n5086), .CK(clock), .Q(
        \registres[21][7] ) );
  FLIP_FLOP_D \registres_reg[21][6]  ( .D(n5085), .CK(clock), .Q(
        \registres[21][6] ) );
  FLIP_FLOP_D \registres_reg[21][5]  ( .D(n5084), .CK(clock), .Q(
        \registres[21][5] ) );
  FLIP_FLOP_D \registres_reg[21][4]  ( .D(n5083), .CK(clock), .Q(
        \registres[21][4] ) );
  FLIP_FLOP_D \registres_reg[21][3]  ( .D(n5082), .CK(clock), .Q(
        \registres[21][3] ) );
  FLIP_FLOP_D \registres_reg[21][2]  ( .D(n5081), .CK(clock), .Q(
        \registres[21][2] ) );
  FLIP_FLOP_D \registres_reg[21][1]  ( .D(n5080), .CK(clock), .Q(
        \registres[21][1] ) );
  FLIP_FLOP_D \registres_reg[21][0]  ( .D(n5079), .CK(clock), .Q(
        \registres[21][0] ) );
  FLIP_FLOP_D \registres_reg[22][31]  ( .D(n5078), .CK(clock), .Q(
        \registres[22][31] ) );
  FLIP_FLOP_D \registres_reg[22][30]  ( .D(n5077), .CK(clock), .Q(
        \registres[22][30] ) );
  FLIP_FLOP_D \registres_reg[22][29]  ( .D(n5076), .CK(clock), .Q(
        \registres[22][29] ) );
  FLIP_FLOP_D \registres_reg[22][28]  ( .D(n5075), .CK(clock), .Q(
        \registres[22][28] ) );
  FLIP_FLOP_D \registres_reg[22][27]  ( .D(n5074), .CK(clock), .Q(
        \registres[22][27] ) );
  FLIP_FLOP_D \registres_reg[22][26]  ( .D(n5073), .CK(clock), .Q(
        \registres[22][26] ) );
  FLIP_FLOP_D \registres_reg[22][25]  ( .D(n5072), .CK(clock), .Q(
        \registres[22][25] ) );
  FLIP_FLOP_D \registres_reg[22][24]  ( .D(n5071), .CK(clock), .Q(
        \registres[22][24] ) );
  FLIP_FLOP_D \registres_reg[22][23]  ( .D(n5070), .CK(clock), .Q(
        \registres[22][23] ) );
  FLIP_FLOP_D \registres_reg[22][22]  ( .D(n5069), .CK(clock), .Q(
        \registres[22][22] ) );
  FLIP_FLOP_D \registres_reg[22][21]  ( .D(n5068), .CK(clock), .Q(
        \registres[22][21] ) );
  FLIP_FLOP_D \registres_reg[22][20]  ( .D(n5067), .CK(clock), .Q(
        \registres[22][20] ) );
  FLIP_FLOP_D \registres_reg[22][19]  ( .D(n5066), .CK(clock), .Q(
        \registres[22][19] ) );
  FLIP_FLOP_D \registres_reg[22][18]  ( .D(n5065), .CK(clock), .Q(
        \registres[22][18] ) );
  FLIP_FLOP_D \registres_reg[22][17]  ( .D(n5064), .CK(clock), .Q(
        \registres[22][17] ) );
  FLIP_FLOP_D \registres_reg[22][16]  ( .D(n5063), .CK(clock), .Q(
        \registres[22][16] ) );
  FLIP_FLOP_D \registres_reg[22][15]  ( .D(n5062), .CK(clock), .Q(
        \registres[22][15] ) );
  FLIP_FLOP_D \registres_reg[22][14]  ( .D(n5061), .CK(clock), .Q(
        \registres[22][14] ) );
  FLIP_FLOP_D \registres_reg[22][13]  ( .D(n5060), .CK(clock), .Q(
        \registres[22][13] ) );
  FLIP_FLOP_D \registres_reg[22][12]  ( .D(n5059), .CK(clock), .Q(
        \registres[22][12] ) );
  FLIP_FLOP_D \registres_reg[22][11]  ( .D(n5058), .CK(clock), .Q(
        \registres[22][11] ) );
  FLIP_FLOP_D \registres_reg[22][10]  ( .D(n5057), .CK(clock), .Q(
        \registres[22][10] ) );
  FLIP_FLOP_D \registres_reg[22][9]  ( .D(n5056), .CK(clock), .Q(
        \registres[22][9] ) );
  FLIP_FLOP_D \registres_reg[22][8]  ( .D(n5055), .CK(clock), .Q(
        \registres[22][8] ) );
  FLIP_FLOP_D \registres_reg[22][7]  ( .D(n5054), .CK(clock), .Q(
        \registres[22][7] ) );
  FLIP_FLOP_D \registres_reg[22][6]  ( .D(n5053), .CK(clock), .Q(
        \registres[22][6] ) );
  FLIP_FLOP_D \registres_reg[22][5]  ( .D(n5052), .CK(clock), .Q(
        \registres[22][5] ) );
  FLIP_FLOP_D \registres_reg[22][4]  ( .D(n5051), .CK(clock), .Q(
        \registres[22][4] ) );
  FLIP_FLOP_D \registres_reg[22][3]  ( .D(n5050), .CK(clock), .Q(
        \registres[22][3] ) );
  FLIP_FLOP_D \registres_reg[22][2]  ( .D(n5049), .CK(clock), .Q(
        \registres[22][2] ) );
  FLIP_FLOP_D \registres_reg[22][1]  ( .D(n5048), .CK(clock), .Q(
        \registres[22][1] ) );
  FLIP_FLOP_D \registres_reg[22][0]  ( .D(n5047), .CK(clock), .Q(
        \registres[22][0] ) );
  FLIP_FLOP_D \registres_reg[23][31]  ( .D(n5046), .CK(clock), .Q(
        \registres[23][31] ) );
  FLIP_FLOP_D \registres_reg[23][30]  ( .D(n5045), .CK(clock), .Q(
        \registres[23][30] ) );
  FLIP_FLOP_D \registres_reg[23][29]  ( .D(n5044), .CK(clock), .Q(
        \registres[23][29] ) );
  FLIP_FLOP_D \registres_reg[23][28]  ( .D(n5043), .CK(clock), .Q(
        \registres[23][28] ) );
  FLIP_FLOP_D \registres_reg[23][27]  ( .D(n5042), .CK(clock), .Q(
        \registres[23][27] ) );
  FLIP_FLOP_D \registres_reg[23][26]  ( .D(n5041), .CK(clock), .Q(
        \registres[23][26] ) );
  FLIP_FLOP_D \registres_reg[23][25]  ( .D(n5040), .CK(clock), .Q(
        \registres[23][25] ) );
  FLIP_FLOP_D \registres_reg[23][24]  ( .D(n5039), .CK(clock), .Q(
        \registres[23][24] ) );
  FLIP_FLOP_D \registres_reg[23][23]  ( .D(n5038), .CK(clock), .Q(
        \registres[23][23] ) );
  FLIP_FLOP_D \registres_reg[23][22]  ( .D(n5037), .CK(clock), .Q(
        \registres[23][22] ) );
  FLIP_FLOP_D \registres_reg[23][21]  ( .D(n5036), .CK(clock), .Q(
        \registres[23][21] ) );
  FLIP_FLOP_D \registres_reg[23][20]  ( .D(n5035), .CK(clock), .Q(
        \registres[23][20] ) );
  FLIP_FLOP_D \registres_reg[23][19]  ( .D(n5034), .CK(clock), .Q(
        \registres[23][19] ) );
  FLIP_FLOP_D \registres_reg[23][18]  ( .D(n5033), .CK(clock), .Q(
        \registres[23][18] ) );
  FLIP_FLOP_D \registres_reg[23][17]  ( .D(n5032), .CK(clock), .Q(
        \registres[23][17] ) );
  FLIP_FLOP_D \registres_reg[23][16]  ( .D(n5031), .CK(clock), .Q(
        \registres[23][16] ) );
  FLIP_FLOP_D \registres_reg[23][15]  ( .D(n5030), .CK(clock), .Q(
        \registres[23][15] ) );
  FLIP_FLOP_D \registres_reg[23][14]  ( .D(n5029), .CK(clock), .Q(
        \registres[23][14] ) );
  FLIP_FLOP_D \registres_reg[23][13]  ( .D(n5028), .CK(clock), .Q(
        \registres[23][13] ) );
  FLIP_FLOP_D \registres_reg[23][12]  ( .D(n5027), .CK(clock), .Q(
        \registres[23][12] ) );
  FLIP_FLOP_D \registres_reg[23][11]  ( .D(n5026), .CK(clock), .Q(
        \registres[23][11] ) );
  FLIP_FLOP_D \registres_reg[23][10]  ( .D(n5025), .CK(clock), .Q(
        \registres[23][10] ) );
  FLIP_FLOP_D \registres_reg[23][9]  ( .D(n5024), .CK(clock), .Q(
        \registres[23][9] ) );
  FLIP_FLOP_D \registres_reg[23][8]  ( .D(n5023), .CK(clock), .Q(
        \registres[23][8] ) );
  FLIP_FLOP_D \registres_reg[23][7]  ( .D(n5022), .CK(clock), .Q(
        \registres[23][7] ) );
  FLIP_FLOP_D \registres_reg[23][6]  ( .D(n5021), .CK(clock), .Q(
        \registres[23][6] ) );
  FLIP_FLOP_D \registres_reg[23][5]  ( .D(n5020), .CK(clock), .Q(
        \registres[23][5] ) );
  FLIP_FLOP_D \registres_reg[23][4]  ( .D(n5019), .CK(clock), .Q(
        \registres[23][4] ) );
  FLIP_FLOP_D \registres_reg[23][3]  ( .D(n5018), .CK(clock), .Q(
        \registres[23][3] ) );
  FLIP_FLOP_D \registres_reg[23][2]  ( .D(n5017), .CK(clock), .Q(
        \registres[23][2] ) );
  FLIP_FLOP_D \registres_reg[23][1]  ( .D(n5016), .CK(clock), .Q(
        \registres[23][1] ) );
  FLIP_FLOP_D \registres_reg[23][0]  ( .D(n5015), .CK(clock), .Q(
        \registres[23][0] ) );
  FLIP_FLOP_D \registres_reg[24][31]  ( .D(n5014), .CK(clock), .Q(
        \registres[24][31] ) );
  FLIP_FLOP_D \registres_reg[24][30]  ( .D(n5013), .CK(clock), .Q(
        \registres[24][30] ) );
  FLIP_FLOP_D \registres_reg[24][29]  ( .D(n5012), .CK(clock), .Q(
        \registres[24][29] ) );
  FLIP_FLOP_D \registres_reg[24][28]  ( .D(n5011), .CK(clock), .Q(
        \registres[24][28] ) );
  FLIP_FLOP_D \registres_reg[24][27]  ( .D(n5010), .CK(clock), .Q(
        \registres[24][27] ) );
  FLIP_FLOP_D \registres_reg[24][26]  ( .D(n5009), .CK(clock), .Q(
        \registres[24][26] ) );
  FLIP_FLOP_D \registres_reg[24][25]  ( .D(n5008), .CK(clock), .Q(
        \registres[24][25] ) );
  FLIP_FLOP_D \registres_reg[24][24]  ( .D(n5007), .CK(clock), .Q(
        \registres[24][24] ) );
  FLIP_FLOP_D \registres_reg[24][23]  ( .D(n5006), .CK(clock), .Q(
        \registres[24][23] ) );
  FLIP_FLOP_D \registres_reg[24][22]  ( .D(n5005), .CK(clock), .Q(
        \registres[24][22] ) );
  FLIP_FLOP_D \registres_reg[24][21]  ( .D(n5004), .CK(clock), .Q(
        \registres[24][21] ) );
  FLIP_FLOP_D \registres_reg[24][20]  ( .D(n5003), .CK(clock), .Q(
        \registres[24][20] ) );
  FLIP_FLOP_D \registres_reg[24][19]  ( .D(n5002), .CK(clock), .Q(
        \registres[24][19] ) );
  FLIP_FLOP_D \registres_reg[24][18]  ( .D(n5001), .CK(clock), .Q(
        \registres[24][18] ) );
  FLIP_FLOP_D \registres_reg[24][17]  ( .D(n5000), .CK(clock), .Q(
        \registres[24][17] ) );
  FLIP_FLOP_D \registres_reg[24][16]  ( .D(n4999), .CK(clock), .Q(
        \registres[24][16] ) );
  FLIP_FLOP_D \registres_reg[24][15]  ( .D(n4998), .CK(clock), .Q(
        \registres[24][15] ) );
  FLIP_FLOP_D \registres_reg[24][14]  ( .D(n4997), .CK(clock), .Q(
        \registres[24][14] ) );
  FLIP_FLOP_D \registres_reg[24][13]  ( .D(n4996), .CK(clock), .Q(
        \registres[24][13] ) );
  FLIP_FLOP_D \registres_reg[24][12]  ( .D(n4995), .CK(clock), .Q(
        \registres[24][12] ) );
  FLIP_FLOP_D \registres_reg[24][11]  ( .D(n4994), .CK(clock), .Q(
        \registres[24][11] ) );
  FLIP_FLOP_D \registres_reg[24][10]  ( .D(n4993), .CK(clock), .Q(
        \registres[24][10] ) );
  FLIP_FLOP_D \registres_reg[24][9]  ( .D(n4992), .CK(clock), .Q(
        \registres[24][9] ) );
  FLIP_FLOP_D \registres_reg[24][8]  ( .D(n4991), .CK(clock), .Q(
        \registres[24][8] ) );
  FLIP_FLOP_D \registres_reg[24][7]  ( .D(n4990), .CK(clock), .Q(
        \registres[24][7] ) );
  FLIP_FLOP_D \registres_reg[24][6]  ( .D(n4989), .CK(clock), .Q(
        \registres[24][6] ) );
  FLIP_FLOP_D \registres_reg[24][5]  ( .D(n4988), .CK(clock), .Q(
        \registres[24][5] ) );
  FLIP_FLOP_D \registres_reg[24][4]  ( .D(n4987), .CK(clock), .Q(
        \registres[24][4] ) );
  FLIP_FLOP_D \registres_reg[24][3]  ( .D(n4986), .CK(clock), .Q(
        \registres[24][3] ) );
  FLIP_FLOP_D \registres_reg[24][2]  ( .D(n4985), .CK(clock), .Q(
        \registres[24][2] ) );
  FLIP_FLOP_D \registres_reg[24][1]  ( .D(n4984), .CK(clock), .Q(
        \registres[24][1] ) );
  FLIP_FLOP_D \registres_reg[24][0]  ( .D(n4983), .CK(clock), .Q(
        \registres[24][0] ) );
  FLIP_FLOP_D \registres_reg[25][31]  ( .D(n4982), .CK(clock), .Q(
        \registres[25][31] ) );
  FLIP_FLOP_D \registres_reg[25][30]  ( .D(n4981), .CK(clock), .Q(
        \registres[25][30] ) );
  FLIP_FLOP_D \registres_reg[25][29]  ( .D(n4980), .CK(clock), .Q(
        \registres[25][29] ) );
  FLIP_FLOP_D \registres_reg[25][28]  ( .D(n4979), .CK(clock), .Q(
        \registres[25][28] ) );
  FLIP_FLOP_D \registres_reg[25][27]  ( .D(n4978), .CK(clock), .Q(
        \registres[25][27] ) );
  FLIP_FLOP_D \registres_reg[25][26]  ( .D(n4977), .CK(clock), .Q(
        \registres[25][26] ) );
  FLIP_FLOP_D \registres_reg[25][25]  ( .D(n4976), .CK(clock), .Q(
        \registres[25][25] ) );
  FLIP_FLOP_D \registres_reg[25][24]  ( .D(n4975), .CK(clock), .Q(
        \registres[25][24] ) );
  FLIP_FLOP_D \registres_reg[25][23]  ( .D(n4974), .CK(clock), .Q(
        \registres[25][23] ) );
  FLIP_FLOP_D \registres_reg[25][22]  ( .D(n4973), .CK(clock), .Q(
        \registres[25][22] ) );
  FLIP_FLOP_D \registres_reg[25][21]  ( .D(n4972), .CK(clock), .Q(
        \registres[25][21] ) );
  FLIP_FLOP_D \registres_reg[25][20]  ( .D(n4971), .CK(clock), .Q(
        \registres[25][20] ) );
  FLIP_FLOP_D \registres_reg[25][19]  ( .D(n4970), .CK(clock), .Q(
        \registres[25][19] ) );
  FLIP_FLOP_D \registres_reg[25][18]  ( .D(n4969), .CK(clock), .Q(
        \registres[25][18] ) );
  FLIP_FLOP_D \registres_reg[25][17]  ( .D(n4968), .CK(clock), .Q(
        \registres[25][17] ) );
  FLIP_FLOP_D \registres_reg[25][16]  ( .D(n4967), .CK(clock), .Q(
        \registres[25][16] ) );
  FLIP_FLOP_D \registres_reg[25][15]  ( .D(n4966), .CK(clock), .Q(
        \registres[25][15] ) );
  FLIP_FLOP_D \registres_reg[25][14]  ( .D(n4965), .CK(clock), .Q(
        \registres[25][14] ) );
  FLIP_FLOP_D \registres_reg[25][13]  ( .D(n4964), .CK(clock), .Q(
        \registres[25][13] ) );
  FLIP_FLOP_D \registres_reg[25][12]  ( .D(n4963), .CK(clock), .Q(
        \registres[25][12] ) );
  FLIP_FLOP_D \registres_reg[25][11]  ( .D(n4962), .CK(clock), .Q(
        \registres[25][11] ) );
  FLIP_FLOP_D \registres_reg[25][10]  ( .D(n4961), .CK(clock), .Q(
        \registres[25][10] ) );
  FLIP_FLOP_D \registres_reg[25][9]  ( .D(n4960), .CK(clock), .Q(
        \registres[25][9] ) );
  FLIP_FLOP_D \registres_reg[25][8]  ( .D(n4959), .CK(clock), .Q(
        \registres[25][8] ) );
  FLIP_FLOP_D \registres_reg[25][7]  ( .D(n4958), .CK(clock), .Q(
        \registres[25][7] ) );
  FLIP_FLOP_D \registres_reg[25][6]  ( .D(n4957), .CK(clock), .Q(
        \registres[25][6] ) );
  FLIP_FLOP_D \registres_reg[25][5]  ( .D(n4956), .CK(clock), .Q(
        \registres[25][5] ) );
  FLIP_FLOP_D \registres_reg[25][4]  ( .D(n4955), .CK(clock), .Q(
        \registres[25][4] ) );
  FLIP_FLOP_D \registres_reg[25][3]  ( .D(n4954), .CK(clock), .Q(
        \registres[25][3] ) );
  FLIP_FLOP_D \registres_reg[25][2]  ( .D(n4953), .CK(clock), .Q(
        \registres[25][2] ) );
  FLIP_FLOP_D \registres_reg[25][1]  ( .D(n4952), .CK(clock), .Q(
        \registres[25][1] ) );
  FLIP_FLOP_D \registres_reg[25][0]  ( .D(n4951), .CK(clock), .Q(
        \registres[25][0] ) );
  FLIP_FLOP_D \registres_reg[26][31]  ( .D(n4950), .CK(clock), .Q(
        \registres[26][31] ) );
  FLIP_FLOP_D \registres_reg[26][30]  ( .D(n4949), .CK(clock), .Q(
        \registres[26][30] ) );
  FLIP_FLOP_D \registres_reg[26][29]  ( .D(n4948), .CK(clock), .Q(
        \registres[26][29] ) );
  FLIP_FLOP_D \registres_reg[26][28]  ( .D(n4947), .CK(clock), .Q(
        \registres[26][28] ) );
  FLIP_FLOP_D \registres_reg[26][27]  ( .D(n4946), .CK(clock), .Q(
        \registres[26][27] ) );
  FLIP_FLOP_D \registres_reg[26][26]  ( .D(n4945), .CK(clock), .Q(
        \registres[26][26] ) );
  FLIP_FLOP_D \registres_reg[26][25]  ( .D(n4944), .CK(clock), .Q(
        \registres[26][25] ) );
  FLIP_FLOP_D \registres_reg[26][24]  ( .D(n4943), .CK(clock), .Q(
        \registres[26][24] ) );
  FLIP_FLOP_D \registres_reg[26][23]  ( .D(n4942), .CK(clock), .Q(
        \registres[26][23] ) );
  FLIP_FLOP_D \registres_reg[26][22]  ( .D(n4941), .CK(clock), .Q(
        \registres[26][22] ) );
  FLIP_FLOP_D \registres_reg[26][21]  ( .D(n4940), .CK(clock), .Q(
        \registres[26][21] ) );
  FLIP_FLOP_D \registres_reg[26][20]  ( .D(n4939), .CK(clock), .Q(
        \registres[26][20] ) );
  FLIP_FLOP_D \registres_reg[26][19]  ( .D(n4938), .CK(clock), .Q(
        \registres[26][19] ) );
  FLIP_FLOP_D \registres_reg[26][18]  ( .D(n4937), .CK(clock), .Q(
        \registres[26][18] ) );
  FLIP_FLOP_D \registres_reg[26][17]  ( .D(n4936), .CK(clock), .Q(
        \registres[26][17] ) );
  FLIP_FLOP_D \registres_reg[26][16]  ( .D(n4935), .CK(clock), .Q(
        \registres[26][16] ) );
  FLIP_FLOP_D \registres_reg[26][15]  ( .D(n4934), .CK(clock), .Q(
        \registres[26][15] ) );
  FLIP_FLOP_D \registres_reg[26][14]  ( .D(n4933), .CK(clock), .Q(
        \registres[26][14] ) );
  FLIP_FLOP_D \registres_reg[26][13]  ( .D(n4932), .CK(clock), .Q(
        \registres[26][13] ) );
  FLIP_FLOP_D \registres_reg[26][12]  ( .D(n4931), .CK(clock), .Q(
        \registres[26][12] ) );
  FLIP_FLOP_D \registres_reg[26][11]  ( .D(n4930), .CK(clock), .Q(
        \registres[26][11] ) );
  FLIP_FLOP_D \registres_reg[26][10]  ( .D(n4929), .CK(clock), .Q(
        \registres[26][10] ) );
  FLIP_FLOP_D \registres_reg[26][9]  ( .D(n4928), .CK(clock), .Q(
        \registres[26][9] ) );
  FLIP_FLOP_D \registres_reg[26][8]  ( .D(n4927), .CK(clock), .Q(
        \registres[26][8] ) );
  FLIP_FLOP_D \registres_reg[26][7]  ( .D(n4926), .CK(clock), .Q(
        \registres[26][7] ) );
  FLIP_FLOP_D \registres_reg[26][6]  ( .D(n4925), .CK(clock), .Q(
        \registres[26][6] ) );
  FLIP_FLOP_D \registres_reg[26][5]  ( .D(n4924), .CK(clock), .Q(
        \registres[26][5] ) );
  FLIP_FLOP_D \registres_reg[26][4]  ( .D(n4923), .CK(clock), .Q(
        \registres[26][4] ) );
  FLIP_FLOP_D \registres_reg[26][3]  ( .D(n4922), .CK(clock), .Q(
        \registres[26][3] ) );
  FLIP_FLOP_D \registres_reg[26][2]  ( .D(n4921), .CK(clock), .Q(
        \registres[26][2] ) );
  FLIP_FLOP_D \registres_reg[26][1]  ( .D(n4920), .CK(clock), .Q(
        \registres[26][1] ) );
  FLIP_FLOP_D \registres_reg[26][0]  ( .D(n4919), .CK(clock), .Q(
        \registres[26][0] ) );
  FLIP_FLOP_D \registres_reg[27][31]  ( .D(n4918), .CK(clock), .Q(
        \registres[27][31] ) );
  FLIP_FLOP_D \registres_reg[27][30]  ( .D(n4917), .CK(clock), .Q(
        \registres[27][30] ) );
  FLIP_FLOP_D \registres_reg[27][29]  ( .D(n4916), .CK(clock), .Q(
        \registres[27][29] ) );
  FLIP_FLOP_D \registres_reg[27][28]  ( .D(n4915), .CK(clock), .Q(
        \registres[27][28] ) );
  FLIP_FLOP_D \registres_reg[27][27]  ( .D(n4914), .CK(clock), .Q(
        \registres[27][27] ) );
  FLIP_FLOP_D \registres_reg[27][26]  ( .D(n4913), .CK(clock), .Q(
        \registres[27][26] ) );
  FLIP_FLOP_D \registres_reg[27][25]  ( .D(n4912), .CK(clock), .Q(
        \registres[27][25] ) );
  FLIP_FLOP_D \registres_reg[27][24]  ( .D(n4911), .CK(clock), .Q(
        \registres[27][24] ) );
  FLIP_FLOP_D \registres_reg[27][23]  ( .D(n4910), .CK(clock), .Q(
        \registres[27][23] ) );
  FLIP_FLOP_D \registres_reg[27][22]  ( .D(n4909), .CK(clock), .Q(
        \registres[27][22] ) );
  FLIP_FLOP_D \registres_reg[27][21]  ( .D(n4908), .CK(clock), .Q(
        \registres[27][21] ) );
  FLIP_FLOP_D \registres_reg[27][20]  ( .D(n4907), .CK(clock), .Q(
        \registres[27][20] ) );
  FLIP_FLOP_D \registres_reg[27][19]  ( .D(n4906), .CK(clock), .Q(
        \registres[27][19] ) );
  FLIP_FLOP_D \registres_reg[27][18]  ( .D(n4905), .CK(clock), .Q(
        \registres[27][18] ) );
  FLIP_FLOP_D \registres_reg[27][17]  ( .D(n4904), .CK(clock), .Q(
        \registres[27][17] ) );
  FLIP_FLOP_D \registres_reg[27][16]  ( .D(n4903), .CK(clock), .Q(
        \registres[27][16] ) );
  FLIP_FLOP_D \registres_reg[27][15]  ( .D(n4902), .CK(clock), .Q(
        \registres[27][15] ) );
  FLIP_FLOP_D \registres_reg[27][14]  ( .D(n4901), .CK(clock), .Q(
        \registres[27][14] ) );
  FLIP_FLOP_D \registres_reg[27][13]  ( .D(n4900), .CK(clock), .Q(
        \registres[27][13] ) );
  FLIP_FLOP_D \registres_reg[27][12]  ( .D(n4899), .CK(clock), .Q(
        \registres[27][12] ) );
  FLIP_FLOP_D \registres_reg[27][11]  ( .D(n4898), .CK(clock), .Q(
        \registres[27][11] ) );
  FLIP_FLOP_D \registres_reg[27][10]  ( .D(n4897), .CK(clock), .Q(
        \registres[27][10] ) );
  FLIP_FLOP_D \registres_reg[27][9]  ( .D(n4896), .CK(clock), .Q(
        \registres[27][9] ) );
  FLIP_FLOP_D \registres_reg[27][8]  ( .D(n4895), .CK(clock), .Q(
        \registres[27][8] ) );
  FLIP_FLOP_D \registres_reg[27][7]  ( .D(n4894), .CK(clock), .Q(
        \registres[27][7] ) );
  FLIP_FLOP_D \registres_reg[27][6]  ( .D(n4893), .CK(clock), .Q(
        \registres[27][6] ) );
  FLIP_FLOP_D \registres_reg[27][5]  ( .D(n4892), .CK(clock), .Q(
        \registres[27][5] ) );
  FLIP_FLOP_D \registres_reg[27][4]  ( .D(n4891), .CK(clock), .Q(
        \registres[27][4] ) );
  FLIP_FLOP_D \registres_reg[27][3]  ( .D(n4890), .CK(clock), .Q(
        \registres[27][3] ) );
  FLIP_FLOP_D \registres_reg[27][2]  ( .D(n4889), .CK(clock), .Q(
        \registres[27][2] ) );
  FLIP_FLOP_D \registres_reg[27][1]  ( .D(n4888), .CK(clock), .Q(
        \registres[27][1] ) );
  FLIP_FLOP_D \registres_reg[27][0]  ( .D(n4887), .CK(clock), .Q(
        \registres[27][0] ) );
  FLIP_FLOP_D \registres_reg[28][31]  ( .D(n4886), .CK(clock), .Q(
        \registres[28][31] ) );
  FLIP_FLOP_D \registres_reg[28][30]  ( .D(n4885), .CK(clock), .Q(
        \registres[28][30] ) );
  FLIP_FLOP_D \registres_reg[28][29]  ( .D(n4884), .CK(clock), .Q(
        \registres[28][29] ) );
  FLIP_FLOP_D \registres_reg[28][28]  ( .D(n4883), .CK(clock), .Q(
        \registres[28][28] ) );
  FLIP_FLOP_D \registres_reg[28][27]  ( .D(n4882), .CK(clock), .Q(
        \registres[28][27] ) );
  FLIP_FLOP_D \registres_reg[28][26]  ( .D(n4881), .CK(clock), .Q(
        \registres[28][26] ) );
  FLIP_FLOP_D \registres_reg[28][25]  ( .D(n4880), .CK(clock), .Q(
        \registres[28][25] ) );
  FLIP_FLOP_D \registres_reg[28][24]  ( .D(n4879), .CK(clock), .Q(
        \registres[28][24] ) );
  FLIP_FLOP_D \registres_reg[28][23]  ( .D(n4878), .CK(clock), .Q(
        \registres[28][23] ) );
  FLIP_FLOP_D \registres_reg[28][22]  ( .D(n4877), .CK(clock), .Q(
        \registres[28][22] ) );
  FLIP_FLOP_D \registres_reg[28][21]  ( .D(n4876), .CK(clock), .Q(
        \registres[28][21] ) );
  FLIP_FLOP_D \registres_reg[28][20]  ( .D(n4875), .CK(clock), .Q(
        \registres[28][20] ) );
  FLIP_FLOP_D \registres_reg[28][19]  ( .D(n4874), .CK(clock), .Q(
        \registres[28][19] ) );
  FLIP_FLOP_D \registres_reg[28][18]  ( .D(n4873), .CK(clock), .Q(
        \registres[28][18] ) );
  FLIP_FLOP_D \registres_reg[28][17]  ( .D(n4872), .CK(clock), .Q(
        \registres[28][17] ) );
  FLIP_FLOP_D \registres_reg[28][16]  ( .D(n4871), .CK(clock), .Q(
        \registres[28][16] ) );
  FLIP_FLOP_D \registres_reg[28][15]  ( .D(n4870), .CK(clock), .Q(
        \registres[28][15] ) );
  FLIP_FLOP_D \registres_reg[28][14]  ( .D(n4869), .CK(clock), .Q(
        \registres[28][14] ) );
  FLIP_FLOP_D \registres_reg[28][13]  ( .D(n4868), .CK(clock), .Q(
        \registres[28][13] ) );
  FLIP_FLOP_D \registres_reg[28][12]  ( .D(n4867), .CK(clock), .Q(
        \registres[28][12] ) );
  FLIP_FLOP_D \registres_reg[28][11]  ( .D(n4866), .CK(clock), .Q(
        \registres[28][11] ) );
  FLIP_FLOP_D \registres_reg[28][10]  ( .D(n4865), .CK(clock), .Q(
        \registres[28][10] ) );
  FLIP_FLOP_D \registres_reg[28][9]  ( .D(n4864), .CK(clock), .Q(
        \registres[28][9] ) );
  FLIP_FLOP_D \registres_reg[28][8]  ( .D(n4863), .CK(clock), .Q(
        \registres[28][8] ) );
  FLIP_FLOP_D \registres_reg[28][7]  ( .D(n4862), .CK(clock), .Q(
        \registres[28][7] ) );
  FLIP_FLOP_D \registres_reg[28][6]  ( .D(n4861), .CK(clock), .Q(
        \registres[28][6] ) );
  FLIP_FLOP_D \registres_reg[28][5]  ( .D(n4860), .CK(clock), .Q(
        \registres[28][5] ) );
  FLIP_FLOP_D \registres_reg[28][4]  ( .D(n4859), .CK(clock), .Q(
        \registres[28][4] ) );
  FLIP_FLOP_D \registres_reg[28][3]  ( .D(n4858), .CK(clock), .Q(
        \registres[28][3] ) );
  FLIP_FLOP_D \registres_reg[28][2]  ( .D(n4857), .CK(clock), .Q(
        \registres[28][2] ) );
  FLIP_FLOP_D \registres_reg[28][1]  ( .D(n4856), .CK(clock), .Q(
        \registres[28][1] ) );
  FLIP_FLOP_D \registres_reg[28][0]  ( .D(n4855), .CK(clock), .Q(
        \registres[28][0] ) );
  FLIP_FLOP_D \registres_reg[29][31]  ( .D(n4854), .CK(clock), .Q(
        \registres[29][31] ) );
  FLIP_FLOP_D \registres_reg[29][30]  ( .D(n4853), .CK(clock), .Q(
        \registres[29][30] ) );
  FLIP_FLOP_D \registres_reg[29][29]  ( .D(n4852), .CK(clock), .Q(
        \registres[29][29] ) );
  FLIP_FLOP_D \registres_reg[29][28]  ( .D(n4851), .CK(clock), .Q(
        \registres[29][28] ) );
  FLIP_FLOP_D \registres_reg[29][27]  ( .D(n4850), .CK(clock), .Q(
        \registres[29][27] ) );
  FLIP_FLOP_D \registres_reg[29][26]  ( .D(n4849), .CK(clock), .Q(
        \registres[29][26] ) );
  FLIP_FLOP_D \registres_reg[29][25]  ( .D(n4848), .CK(clock), .Q(
        \registres[29][25] ) );
  FLIP_FLOP_D \registres_reg[29][24]  ( .D(n4847), .CK(clock), .Q(
        \registres[29][24] ) );
  FLIP_FLOP_D \registres_reg[29][23]  ( .D(n4846), .CK(clock), .Q(
        \registres[29][23] ) );
  FLIP_FLOP_D \registres_reg[29][22]  ( .D(n4845), .CK(clock), .Q(
        \registres[29][22] ) );
  FLIP_FLOP_D \registres_reg[29][21]  ( .D(n4844), .CK(clock), .Q(
        \registres[29][21] ) );
  FLIP_FLOP_D \registres_reg[29][20]  ( .D(n4843), .CK(clock), .Q(
        \registres[29][20] ) );
  FLIP_FLOP_D \registres_reg[29][19]  ( .D(n4842), .CK(clock), .Q(
        \registres[29][19] ) );
  FLIP_FLOP_D \registres_reg[29][18]  ( .D(n4841), .CK(clock), .Q(
        \registres[29][18] ) );
  FLIP_FLOP_D \registres_reg[29][17]  ( .D(n4840), .CK(clock), .Q(
        \registres[29][17] ) );
  FLIP_FLOP_D \registres_reg[29][16]  ( .D(n4839), .CK(clock), .Q(
        \registres[29][16] ) );
  FLIP_FLOP_D \registres_reg[29][15]  ( .D(n4838), .CK(clock), .Q(
        \registres[29][15] ) );
  FLIP_FLOP_D \registres_reg[29][14]  ( .D(n4837), .CK(clock), .Q(
        \registres[29][14] ) );
  FLIP_FLOP_D \registres_reg[29][13]  ( .D(n4836), .CK(clock), .Q(
        \registres[29][13] ) );
  FLIP_FLOP_D \registres_reg[29][12]  ( .D(n4835), .CK(clock), .Q(
        \registres[29][12] ) );
  FLIP_FLOP_D \registres_reg[29][11]  ( .D(n4834), .CK(clock), .Q(
        \registres[29][11] ) );
  FLIP_FLOP_D \registres_reg[29][10]  ( .D(n4833), .CK(clock), .Q(
        \registres[29][10] ) );
  FLIP_FLOP_D \registres_reg[29][9]  ( .D(n4832), .CK(clock), .Q(
        \registres[29][9] ) );
  FLIP_FLOP_D \registres_reg[29][8]  ( .D(n4831), .CK(clock), .Q(
        \registres[29][8] ) );
  FLIP_FLOP_D \registres_reg[29][7]  ( .D(n4830), .CK(clock), .Q(
        \registres[29][7] ) );
  FLIP_FLOP_D \registres_reg[29][6]  ( .D(n4829), .CK(clock), .Q(
        \registres[29][6] ) );
  FLIP_FLOP_D \registres_reg[29][5]  ( .D(n4828), .CK(clock), .Q(
        \registres[29][5] ) );
  FLIP_FLOP_D \registres_reg[29][4]  ( .D(n4827), .CK(clock), .Q(
        \registres[29][4] ) );
  FLIP_FLOP_D \registres_reg[29][3]  ( .D(n4826), .CK(clock), .Q(
        \registres[29][3] ) );
  FLIP_FLOP_D \registres_reg[29][2]  ( .D(n4825), .CK(clock), .Q(
        \registres[29][2] ) );
  FLIP_FLOP_D \registres_reg[29][1]  ( .D(n4824), .CK(clock), .Q(
        \registres[29][1] ) );
  FLIP_FLOP_D \registres_reg[29][0]  ( .D(n4823), .CK(clock), .Q(
        \registres[29][0] ) );
  FLIP_FLOP_D \registres_reg[30][31]  ( .D(n4822), .CK(clock), .Q(
        \registres[30][31] ) );
  FLIP_FLOP_D \registres_reg[30][30]  ( .D(n4821), .CK(clock), .Q(
        \registres[30][30] ) );
  FLIP_FLOP_D \registres_reg[30][29]  ( .D(n4820), .CK(clock), .Q(
        \registres[30][29] ) );
  FLIP_FLOP_D \registres_reg[30][28]  ( .D(n4819), .CK(clock), .Q(
        \registres[30][28] ) );
  FLIP_FLOP_D \registres_reg[30][27]  ( .D(n4818), .CK(clock), .Q(
        \registres[30][27] ) );
  FLIP_FLOP_D \registres_reg[30][26]  ( .D(n4817), .CK(clock), .Q(
        \registres[30][26] ) );
  FLIP_FLOP_D \registres_reg[30][25]  ( .D(n4816), .CK(clock), .Q(
        \registres[30][25] ) );
  FLIP_FLOP_D \registres_reg[30][24]  ( .D(n4815), .CK(clock), .Q(
        \registres[30][24] ) );
  FLIP_FLOP_D \registres_reg[30][23]  ( .D(n4814), .CK(clock), .Q(
        \registres[30][23] ) );
  FLIP_FLOP_D \registres_reg[30][22]  ( .D(n4813), .CK(clock), .Q(
        \registres[30][22] ) );
  FLIP_FLOP_D \registres_reg[30][21]  ( .D(n4812), .CK(clock), .Q(
        \registres[30][21] ) );
  FLIP_FLOP_D \registres_reg[30][20]  ( .D(n4811), .CK(clock), .Q(
        \registres[30][20] ) );
  FLIP_FLOP_D \registres_reg[30][19]  ( .D(n4810), .CK(clock), .Q(
        \registres[30][19] ) );
  FLIP_FLOP_D \registres_reg[30][18]  ( .D(n4809), .CK(clock), .Q(
        \registres[30][18] ) );
  FLIP_FLOP_D \registres_reg[30][17]  ( .D(n4808), .CK(clock), .Q(
        \registres[30][17] ) );
  FLIP_FLOP_D \registres_reg[30][16]  ( .D(n4807), .CK(clock), .Q(
        \registres[30][16] ) );
  FLIP_FLOP_D \registres_reg[30][15]  ( .D(n4806), .CK(clock), .Q(
        \registres[30][15] ) );
  FLIP_FLOP_D \registres_reg[30][14]  ( .D(n4805), .CK(clock), .Q(
        \registres[30][14] ) );
  FLIP_FLOP_D \registres_reg[30][13]  ( .D(n4804), .CK(clock), .Q(
        \registres[30][13] ) );
  FLIP_FLOP_D \registres_reg[30][12]  ( .D(n4803), .CK(clock), .Q(
        \registres[30][12] ) );
  FLIP_FLOP_D \registres_reg[30][11]  ( .D(n4802), .CK(clock), .Q(
        \registres[30][11] ) );
  FLIP_FLOP_D \registres_reg[30][10]  ( .D(n4801), .CK(clock), .Q(
        \registres[30][10] ) );
  FLIP_FLOP_D \registres_reg[30][9]  ( .D(n4800), .CK(clock), .Q(
        \registres[30][9] ) );
  FLIP_FLOP_D \registres_reg[30][8]  ( .D(n4799), .CK(clock), .Q(
        \registres[30][8] ) );
  FLIP_FLOP_D \registres_reg[30][7]  ( .D(n4798), .CK(clock), .Q(
        \registres[30][7] ) );
  FLIP_FLOP_D \registres_reg[30][6]  ( .D(n4797), .CK(clock), .Q(
        \registres[30][6] ) );
  FLIP_FLOP_D \registres_reg[30][5]  ( .D(n4796), .CK(clock), .Q(
        \registres[30][5] ) );
  FLIP_FLOP_D \registres_reg[30][4]  ( .D(n4795), .CK(clock), .Q(
        \registres[30][4] ) );
  FLIP_FLOP_D \registres_reg[30][3]  ( .D(n4794), .CK(clock), .Q(
        \registres[30][3] ) );
  FLIP_FLOP_D \registres_reg[30][2]  ( .D(n4793), .CK(clock), .Q(
        \registres[30][2] ) );
  FLIP_FLOP_D \registres_reg[30][1]  ( .D(n4792), .CK(clock), .Q(
        \registres[30][1] ) );
  FLIP_FLOP_D \registres_reg[30][0]  ( .D(n4791), .CK(clock), .Q(
        \registres[30][0] ) );
  FLIP_FLOP_D \registres_reg[31][31]  ( .D(n4790), .CK(clock), .Q(
        \registres[31][31] ) );
  FLIP_FLOP_D \registres_reg[31][30]  ( .D(n4789), .CK(clock), .Q(
        \registres[31][30] ) );
  FLIP_FLOP_D \registres_reg[31][29]  ( .D(n4788), .CK(clock), .Q(
        \registres[31][29] ) );
  FLIP_FLOP_D \registres_reg[31][28]  ( .D(n4787), .CK(clock), .Q(
        \registres[31][28] ) );
  FLIP_FLOP_D \registres_reg[31][27]  ( .D(n4786), .CK(clock), .Q(
        \registres[31][27] ) );
  FLIP_FLOP_D \registres_reg[31][26]  ( .D(n4785), .CK(clock), .Q(
        \registres[31][26] ) );
  FLIP_FLOP_D \registres_reg[31][25]  ( .D(n4784), .CK(clock), .Q(
        \registres[31][25] ) );
  FLIP_FLOP_D \registres_reg[31][24]  ( .D(n4783), .CK(clock), .Q(
        \registres[31][24] ) );
  FLIP_FLOP_D \registres_reg[31][23]  ( .D(n4782), .CK(clock), .Q(
        \registres[31][23] ) );
  FLIP_FLOP_D \registres_reg[31][22]  ( .D(n4781), .CK(clock), .Q(
        \registres[31][22] ) );
  FLIP_FLOP_D \registres_reg[31][21]  ( .D(n4780), .CK(clock), .Q(
        \registres[31][21] ) );
  FLIP_FLOP_D \registres_reg[31][20]  ( .D(n4779), .CK(clock), .Q(
        \registres[31][20] ) );
  FLIP_FLOP_D \registres_reg[31][19]  ( .D(n4778), .CK(clock), .Q(
        \registres[31][19] ) );
  FLIP_FLOP_D \registres_reg[31][18]  ( .D(n4777), .CK(clock), .Q(
        \registres[31][18] ) );
  FLIP_FLOP_D \registres_reg[31][17]  ( .D(n4776), .CK(clock), .Q(
        \registres[31][17] ) );
  FLIP_FLOP_D \registres_reg[31][16]  ( .D(n4775), .CK(clock), .Q(
        \registres[31][16] ) );
  FLIP_FLOP_D \registres_reg[31][15]  ( .D(n4774), .CK(clock), .Q(
        \registres[31][15] ) );
  FLIP_FLOP_D \registres_reg[31][14]  ( .D(n4773), .CK(clock), .Q(
        \registres[31][14] ) );
  FLIP_FLOP_D \registres_reg[31][13]  ( .D(n4772), .CK(clock), .Q(
        \registres[31][13] ) );
  FLIP_FLOP_D \registres_reg[31][12]  ( .D(n4771), .CK(clock), .Q(
        \registres[31][12] ) );
  FLIP_FLOP_D \registres_reg[31][11]  ( .D(n4770), .CK(clock), .Q(
        \registres[31][11] ) );
  FLIP_FLOP_D \registres_reg[31][10]  ( .D(n4769), .CK(clock), .Q(
        \registres[31][10] ) );
  FLIP_FLOP_D \registres_reg[31][9]  ( .D(n4768), .CK(clock), .Q(
        \registres[31][9] ) );
  FLIP_FLOP_D \registres_reg[31][8]  ( .D(n4767), .CK(clock), .Q(
        \registres[31][8] ) );
  FLIP_FLOP_D \registres_reg[31][7]  ( .D(n4766), .CK(clock), .Q(
        \registres[31][7] ) );
  FLIP_FLOP_D \registres_reg[31][6]  ( .D(n4765), .CK(clock), .Q(
        \registres[31][6] ) );
  FLIP_FLOP_D \registres_reg[31][5]  ( .D(n4764), .CK(clock), .Q(
        \registres[31][5] ) );
  FLIP_FLOP_D \registres_reg[31][4]  ( .D(n4763), .CK(clock), .Q(
        \registres[31][4] ) );
  FLIP_FLOP_D \registres_reg[31][3]  ( .D(n4762), .CK(clock), .Q(
        \registres[31][3] ) );
  FLIP_FLOP_D \registres_reg[31][2]  ( .D(n4761), .CK(clock), .Q(
        \registres[31][2] ) );
  FLIP_FLOP_D \registres_reg[31][1]  ( .D(n4760), .CK(clock), .Q(
        \registres[31][1] ) );
  FLIP_FLOP_D \registres_reg[31][0]  ( .D(n4759), .CK(clock), .Q(
        \registres[31][0] ) );
  NAND_GATE U17 ( .I1(n16), .I2(n17), .O(n4759) );
  NAND_GATE U18 ( .I1(donnee[0]), .I2(n18), .O(n17) );
  NAND_GATE U19 ( .I1(\registres[31][0] ), .I2(n19), .O(n16) );
  NAND_GATE U20 ( .I1(n20), .I2(n21), .O(n4760) );
  NAND_GATE U21 ( .I1(donnee[1]), .I2(n18), .O(n21) );
  NAND_GATE U22 ( .I1(\registres[31][1] ), .I2(n19), .O(n20) );
  NAND_GATE U23 ( .I1(n22), .I2(n23), .O(n4761) );
  NAND_GATE U24 ( .I1(donnee[2]), .I2(n18), .O(n23) );
  NAND_GATE U25 ( .I1(\registres[31][2] ), .I2(n19), .O(n22) );
  NAND_GATE U26 ( .I1(n24), .I2(n25), .O(n4762) );
  NAND_GATE U27 ( .I1(donnee[3]), .I2(n18), .O(n25) );
  NAND_GATE U28 ( .I1(\registres[31][3] ), .I2(n19), .O(n24) );
  NAND_GATE U29 ( .I1(n26), .I2(n27), .O(n4763) );
  NAND_GATE U30 ( .I1(donnee[4]), .I2(n18), .O(n27) );
  NAND_GATE U31 ( .I1(\registres[31][4] ), .I2(n19), .O(n26) );
  NAND_GATE U32 ( .I1(n28), .I2(n29), .O(n4764) );
  NAND_GATE U33 ( .I1(donnee[5]), .I2(n18), .O(n29) );
  NAND_GATE U34 ( .I1(\registres[31][5] ), .I2(n19), .O(n28) );
  NAND_GATE U35 ( .I1(n30), .I2(n31), .O(n4765) );
  NAND_GATE U36 ( .I1(donnee[6]), .I2(n18), .O(n31) );
  NAND_GATE U37 ( .I1(\registres[31][6] ), .I2(n19), .O(n30) );
  NAND_GATE U38 ( .I1(n32), .I2(n33), .O(n4766) );
  NAND_GATE U39 ( .I1(donnee[7]), .I2(n18), .O(n33) );
  NAND_GATE U40 ( .I1(\registres[31][7] ), .I2(n19), .O(n32) );
  NAND_GATE U41 ( .I1(n34), .I2(n35), .O(n4767) );
  NAND_GATE U42 ( .I1(donnee[8]), .I2(n18), .O(n35) );
  NAND_GATE U43 ( .I1(\registres[31][8] ), .I2(n19), .O(n34) );
  NAND_GATE U44 ( .I1(n36), .I2(n37), .O(n4768) );
  NAND_GATE U45 ( .I1(donnee[9]), .I2(n18), .O(n37) );
  NAND_GATE U46 ( .I1(\registres[31][9] ), .I2(n19), .O(n36) );
  NAND_GATE U47 ( .I1(n38), .I2(n39), .O(n4769) );
  NAND_GATE U48 ( .I1(donnee[10]), .I2(n18), .O(n39) );
  NAND_GATE U49 ( .I1(\registres[31][10] ), .I2(n19), .O(n38) );
  NAND_GATE U50 ( .I1(n40), .I2(n41), .O(n4770) );
  NAND_GATE U51 ( .I1(donnee[11]), .I2(n18), .O(n41) );
  NAND_GATE U52 ( .I1(\registres[31][11] ), .I2(n19), .O(n40) );
  NAND_GATE U53 ( .I1(n42), .I2(n43), .O(n4771) );
  NAND_GATE U54 ( .I1(donnee[12]), .I2(n18), .O(n43) );
  NAND_GATE U55 ( .I1(\registres[31][12] ), .I2(n19), .O(n42) );
  NAND_GATE U56 ( .I1(n44), .I2(n45), .O(n4772) );
  NAND_GATE U57 ( .I1(donnee[13]), .I2(n18), .O(n45) );
  NAND_GATE U58 ( .I1(\registres[31][13] ), .I2(n19), .O(n44) );
  NAND_GATE U59 ( .I1(n46), .I2(n47), .O(n4773) );
  NAND_GATE U60 ( .I1(donnee[14]), .I2(n18), .O(n47) );
  NAND_GATE U61 ( .I1(\registres[31][14] ), .I2(n19), .O(n46) );
  NAND_GATE U62 ( .I1(n48), .I2(n49), .O(n4774) );
  NAND_GATE U63 ( .I1(donnee[15]), .I2(n18), .O(n49) );
  NAND_GATE U64 ( .I1(\registres[31][15] ), .I2(n19), .O(n48) );
  NAND_GATE U65 ( .I1(n50), .I2(n51), .O(n4775) );
  NAND_GATE U66 ( .I1(donnee[16]), .I2(n18), .O(n51) );
  NAND_GATE U67 ( .I1(\registres[31][16] ), .I2(n19), .O(n50) );
  NAND_GATE U68 ( .I1(n52), .I2(n53), .O(n4776) );
  NAND_GATE U69 ( .I1(donnee[17]), .I2(n18), .O(n53) );
  NAND_GATE U70 ( .I1(\registres[31][17] ), .I2(n19), .O(n52) );
  NAND_GATE U71 ( .I1(n54), .I2(n55), .O(n4777) );
  NAND_GATE U72 ( .I1(donnee[18]), .I2(n18), .O(n55) );
  NAND_GATE U73 ( .I1(\registres[31][18] ), .I2(n19), .O(n54) );
  NAND_GATE U74 ( .I1(n56), .I2(n57), .O(n4778) );
  NAND_GATE U75 ( .I1(donnee[19]), .I2(n18), .O(n57) );
  NAND_GATE U76 ( .I1(\registres[31][19] ), .I2(n19), .O(n56) );
  NAND_GATE U77 ( .I1(n58), .I2(n59), .O(n4779) );
  NAND_GATE U78 ( .I1(donnee[20]), .I2(n18), .O(n59) );
  NAND_GATE U79 ( .I1(\registres[31][20] ), .I2(n19), .O(n58) );
  NAND_GATE U80 ( .I1(n60), .I2(n61), .O(n4780) );
  NAND_GATE U81 ( .I1(donnee[21]), .I2(n18), .O(n61) );
  NAND_GATE U82 ( .I1(\registres[31][21] ), .I2(n19), .O(n60) );
  NAND_GATE U83 ( .I1(n62), .I2(n63), .O(n4781) );
  NAND_GATE U84 ( .I1(donnee[22]), .I2(n18), .O(n63) );
  NAND_GATE U85 ( .I1(\registres[31][22] ), .I2(n19), .O(n62) );
  NAND_GATE U86 ( .I1(n64), .I2(n65), .O(n4782) );
  NAND_GATE U87 ( .I1(donnee[23]), .I2(n18), .O(n65) );
  NAND_GATE U88 ( .I1(\registres[31][23] ), .I2(n19), .O(n64) );
  NAND_GATE U89 ( .I1(n66), .I2(n67), .O(n4783) );
  NAND_GATE U90 ( .I1(donnee[24]), .I2(n18), .O(n67) );
  NAND_GATE U91 ( .I1(\registres[31][24] ), .I2(n19), .O(n66) );
  NAND_GATE U92 ( .I1(n68), .I2(n69), .O(n4784) );
  NAND_GATE U93 ( .I1(donnee[25]), .I2(n18), .O(n69) );
  NAND_GATE U94 ( .I1(\registres[31][25] ), .I2(n19), .O(n68) );
  NAND_GATE U95 ( .I1(n70), .I2(n71), .O(n4785) );
  NAND_GATE U96 ( .I1(donnee[26]), .I2(n18), .O(n71) );
  NAND_GATE U97 ( .I1(\registres[31][26] ), .I2(n19), .O(n70) );
  NAND_GATE U98 ( .I1(n72), .I2(n73), .O(n4786) );
  NAND_GATE U99 ( .I1(donnee[27]), .I2(n18), .O(n73) );
  NAND_GATE U100 ( .I1(\registres[31][27] ), .I2(n19), .O(n72) );
  NAND_GATE U101 ( .I1(n74), .I2(n75), .O(n4787) );
  NAND_GATE U102 ( .I1(donnee[28]), .I2(n18), .O(n75) );
  NAND_GATE U103 ( .I1(\registres[31][28] ), .I2(n19), .O(n74) );
  NAND_GATE U104 ( .I1(n76), .I2(n77), .O(n4788) );
  NAND_GATE U105 ( .I1(donnee[29]), .I2(n18), .O(n77) );
  NAND_GATE U106 ( .I1(\registres[31][29] ), .I2(n19), .O(n76) );
  NAND_GATE U107 ( .I1(n78), .I2(n79), .O(n4789) );
  NAND_GATE U108 ( .I1(donnee[30]), .I2(n18), .O(n79) );
  NAND_GATE U109 ( .I1(\registres[31][30] ), .I2(n19), .O(n78) );
  NAND_GATE U110 ( .I1(n80), .I2(n81), .O(n4790) );
  NAND_GATE U111 ( .I1(donnee[31]), .I2(n18), .O(n81) );
  AND_GATE U112 ( .I1(n82), .I2(n1), .O(n18) );
  NAND_GATE U113 ( .I1(\registres[31][31] ), .I2(n19), .O(n80) );
  NOR_GATE U114 ( .I1(n82), .I2(reset), .O(n19) );
  AND3_GATE U115 ( .I1(n83), .I2(cmd_ecr), .I3(n84), .O(n82) );
  NAND_GATE U116 ( .I1(n85), .I2(n86), .O(n4791) );
  NAND_GATE U117 ( .I1(n87), .I2(donnee[0]), .O(n86) );
  NAND_GATE U118 ( .I1(\registres[30][0] ), .I2(n88), .O(n85) );
  NAND_GATE U119 ( .I1(n89), .I2(n90), .O(n4792) );
  NAND_GATE U120 ( .I1(n87), .I2(donnee[1]), .O(n90) );
  NAND_GATE U121 ( .I1(\registres[30][1] ), .I2(n88), .O(n89) );
  NAND_GATE U122 ( .I1(n91), .I2(n92), .O(n4793) );
  NAND_GATE U123 ( .I1(n87), .I2(donnee[2]), .O(n92) );
  NAND_GATE U124 ( .I1(\registres[30][2] ), .I2(n88), .O(n91) );
  NAND_GATE U125 ( .I1(n93), .I2(n94), .O(n4794) );
  NAND_GATE U126 ( .I1(n87), .I2(donnee[3]), .O(n94) );
  NAND_GATE U127 ( .I1(\registres[30][3] ), .I2(n88), .O(n93) );
  NAND_GATE U128 ( .I1(n95), .I2(n96), .O(n4795) );
  NAND_GATE U129 ( .I1(n87), .I2(donnee[4]), .O(n96) );
  NAND_GATE U130 ( .I1(\registres[30][4] ), .I2(n88), .O(n95) );
  NAND_GATE U131 ( .I1(n97), .I2(n98), .O(n4796) );
  NAND_GATE U132 ( .I1(n87), .I2(donnee[5]), .O(n98) );
  NAND_GATE U133 ( .I1(\registres[30][5] ), .I2(n88), .O(n97) );
  NAND_GATE U134 ( .I1(n99), .I2(n100), .O(n4797) );
  NAND_GATE U135 ( .I1(n87), .I2(donnee[6]), .O(n100) );
  NAND_GATE U136 ( .I1(\registres[30][6] ), .I2(n88), .O(n99) );
  NAND_GATE U137 ( .I1(n101), .I2(n102), .O(n4798) );
  NAND_GATE U138 ( .I1(n87), .I2(donnee[7]), .O(n102) );
  NAND_GATE U139 ( .I1(\registres[30][7] ), .I2(n88), .O(n101) );
  NAND_GATE U140 ( .I1(n103), .I2(n104), .O(n4799) );
  NAND_GATE U141 ( .I1(n87), .I2(donnee[8]), .O(n104) );
  NAND_GATE U142 ( .I1(\registres[30][8] ), .I2(n88), .O(n103) );
  NAND_GATE U143 ( .I1(n105), .I2(n106), .O(n4800) );
  NAND_GATE U144 ( .I1(n87), .I2(donnee[9]), .O(n106) );
  NAND_GATE U145 ( .I1(\registres[30][9] ), .I2(n88), .O(n105) );
  NAND_GATE U146 ( .I1(n107), .I2(n108), .O(n4801) );
  NAND_GATE U147 ( .I1(n87), .I2(donnee[10]), .O(n108) );
  NAND_GATE U148 ( .I1(\registres[30][10] ), .I2(n88), .O(n107) );
  NAND_GATE U149 ( .I1(n109), .I2(n110), .O(n4802) );
  NAND_GATE U150 ( .I1(n87), .I2(donnee[11]), .O(n110) );
  NAND_GATE U151 ( .I1(\registres[30][11] ), .I2(n88), .O(n109) );
  NAND_GATE U152 ( .I1(n111), .I2(n112), .O(n4803) );
  NAND_GATE U153 ( .I1(n87), .I2(donnee[12]), .O(n112) );
  NAND_GATE U154 ( .I1(\registres[30][12] ), .I2(n88), .O(n111) );
  NAND_GATE U155 ( .I1(n113), .I2(n114), .O(n4804) );
  NAND_GATE U156 ( .I1(n87), .I2(donnee[13]), .O(n114) );
  NAND_GATE U157 ( .I1(\registres[30][13] ), .I2(n88), .O(n113) );
  NAND_GATE U158 ( .I1(n115), .I2(n116), .O(n4805) );
  NAND_GATE U159 ( .I1(n87), .I2(donnee[14]), .O(n116) );
  NAND_GATE U160 ( .I1(\registres[30][14] ), .I2(n88), .O(n115) );
  NAND_GATE U161 ( .I1(n117), .I2(n118), .O(n4806) );
  NAND_GATE U162 ( .I1(n87), .I2(donnee[15]), .O(n118) );
  NAND_GATE U163 ( .I1(\registres[30][15] ), .I2(n88), .O(n117) );
  NAND_GATE U164 ( .I1(n119), .I2(n120), .O(n4807) );
  NAND_GATE U165 ( .I1(n87), .I2(donnee[16]), .O(n120) );
  NAND_GATE U166 ( .I1(\registres[30][16] ), .I2(n88), .O(n119) );
  NAND_GATE U167 ( .I1(n121), .I2(n122), .O(n4808) );
  NAND_GATE U168 ( .I1(n87), .I2(donnee[17]), .O(n122) );
  NAND_GATE U169 ( .I1(\registres[30][17] ), .I2(n88), .O(n121) );
  NAND_GATE U170 ( .I1(n123), .I2(n124), .O(n4809) );
  NAND_GATE U171 ( .I1(n87), .I2(donnee[18]), .O(n124) );
  NAND_GATE U172 ( .I1(\registres[30][18] ), .I2(n88), .O(n123) );
  NAND_GATE U173 ( .I1(n125), .I2(n126), .O(n4810) );
  NAND_GATE U174 ( .I1(n87), .I2(donnee[19]), .O(n126) );
  NAND_GATE U175 ( .I1(\registres[30][19] ), .I2(n88), .O(n125) );
  NAND_GATE U176 ( .I1(n127), .I2(n128), .O(n4811) );
  NAND_GATE U177 ( .I1(n87), .I2(donnee[20]), .O(n128) );
  NAND_GATE U178 ( .I1(\registres[30][20] ), .I2(n88), .O(n127) );
  NAND_GATE U179 ( .I1(n129), .I2(n130), .O(n4812) );
  NAND_GATE U180 ( .I1(n87), .I2(donnee[21]), .O(n130) );
  NAND_GATE U181 ( .I1(\registres[30][21] ), .I2(n88), .O(n129) );
  NAND_GATE U182 ( .I1(n131), .I2(n132), .O(n4813) );
  NAND_GATE U183 ( .I1(n87), .I2(donnee[22]), .O(n132) );
  NAND_GATE U184 ( .I1(\registres[30][22] ), .I2(n88), .O(n131) );
  NAND_GATE U185 ( .I1(n133), .I2(n134), .O(n4814) );
  NAND_GATE U186 ( .I1(n87), .I2(donnee[23]), .O(n134) );
  NAND_GATE U187 ( .I1(\registres[30][23] ), .I2(n88), .O(n133) );
  NAND_GATE U188 ( .I1(n135), .I2(n136), .O(n4815) );
  NAND_GATE U189 ( .I1(n87), .I2(donnee[24]), .O(n136) );
  NAND_GATE U190 ( .I1(\registres[30][24] ), .I2(n88), .O(n135) );
  NAND_GATE U191 ( .I1(n137), .I2(n138), .O(n4816) );
  NAND_GATE U192 ( .I1(n87), .I2(donnee[25]), .O(n138) );
  NAND_GATE U193 ( .I1(\registres[30][25] ), .I2(n88), .O(n137) );
  NAND_GATE U194 ( .I1(n139), .I2(n140), .O(n4817) );
  NAND_GATE U195 ( .I1(n87), .I2(donnee[26]), .O(n140) );
  NAND_GATE U196 ( .I1(\registres[30][26] ), .I2(n88), .O(n139) );
  NAND_GATE U197 ( .I1(n141), .I2(n142), .O(n4818) );
  NAND_GATE U198 ( .I1(n87), .I2(donnee[27]), .O(n142) );
  NAND_GATE U199 ( .I1(\registres[30][27] ), .I2(n88), .O(n141) );
  NAND_GATE U200 ( .I1(n143), .I2(n144), .O(n4819) );
  NAND_GATE U201 ( .I1(n87), .I2(donnee[28]), .O(n144) );
  NAND_GATE U202 ( .I1(\registres[30][28] ), .I2(n88), .O(n143) );
  NAND_GATE U203 ( .I1(n145), .I2(n146), .O(n4820) );
  NAND_GATE U204 ( .I1(n87), .I2(donnee[29]), .O(n146) );
  NAND_GATE U205 ( .I1(\registres[30][29] ), .I2(n88), .O(n145) );
  NAND_GATE U206 ( .I1(n147), .I2(n148), .O(n4821) );
  NAND_GATE U207 ( .I1(n87), .I2(donnee[30]), .O(n148) );
  NAND_GATE U208 ( .I1(\registres[30][30] ), .I2(n88), .O(n147) );
  NAND_GATE U209 ( .I1(n149), .I2(n150), .O(n4822) );
  NAND_GATE U210 ( .I1(n87), .I2(donnee[31]), .O(n150) );
  AND_GATE U211 ( .I1(n151), .I2(n1), .O(n87) );
  NAND_GATE U212 ( .I1(\registres[30][31] ), .I2(n88), .O(n149) );
  NOR_GATE U213 ( .I1(n151), .I2(reset), .O(n88) );
  AND3_GATE U214 ( .I1(n83), .I2(cmd_ecr), .I3(n152), .O(n151) );
  NAND_GATE U215 ( .I1(n153), .I2(n154), .O(n4823) );
  NAND_GATE U216 ( .I1(n155), .I2(donnee[0]), .O(n154) );
  NAND_GATE U217 ( .I1(\registres[29][0] ), .I2(n156), .O(n153) );
  NAND_GATE U218 ( .I1(n157), .I2(n158), .O(n4824) );
  NAND_GATE U219 ( .I1(n155), .I2(donnee[1]), .O(n158) );
  NAND_GATE U220 ( .I1(\registres[29][1] ), .I2(n156), .O(n157) );
  NAND_GATE U221 ( .I1(n159), .I2(n160), .O(n4825) );
  NAND_GATE U222 ( .I1(n155), .I2(donnee[2]), .O(n160) );
  NAND_GATE U223 ( .I1(\registres[29][2] ), .I2(n156), .O(n159) );
  NAND_GATE U224 ( .I1(n161), .I2(n162), .O(n4826) );
  NAND_GATE U225 ( .I1(n155), .I2(donnee[3]), .O(n162) );
  NAND_GATE U226 ( .I1(\registres[29][3] ), .I2(n156), .O(n161) );
  NAND_GATE U227 ( .I1(n163), .I2(n164), .O(n4827) );
  NAND_GATE U228 ( .I1(n155), .I2(donnee[4]), .O(n164) );
  NAND_GATE U229 ( .I1(\registres[29][4] ), .I2(n156), .O(n163) );
  NAND_GATE U230 ( .I1(n165), .I2(n166), .O(n4828) );
  NAND_GATE U231 ( .I1(n155), .I2(donnee[5]), .O(n166) );
  NAND_GATE U232 ( .I1(\registres[29][5] ), .I2(n156), .O(n165) );
  NAND_GATE U233 ( .I1(n167), .I2(n168), .O(n4829) );
  NAND_GATE U234 ( .I1(n155), .I2(donnee[6]), .O(n168) );
  NAND_GATE U235 ( .I1(\registres[29][6] ), .I2(n156), .O(n167) );
  NAND_GATE U236 ( .I1(n169), .I2(n170), .O(n4830) );
  NAND_GATE U237 ( .I1(n155), .I2(donnee[7]), .O(n170) );
  NAND_GATE U238 ( .I1(\registres[29][7] ), .I2(n156), .O(n169) );
  NAND_GATE U239 ( .I1(n171), .I2(n172), .O(n4831) );
  NAND_GATE U240 ( .I1(n155), .I2(donnee[8]), .O(n172) );
  NAND_GATE U241 ( .I1(\registres[29][8] ), .I2(n156), .O(n171) );
  NAND_GATE U242 ( .I1(n173), .I2(n174), .O(n4832) );
  NAND_GATE U243 ( .I1(n155), .I2(donnee[9]), .O(n174) );
  NAND_GATE U244 ( .I1(\registres[29][9] ), .I2(n156), .O(n173) );
  NAND_GATE U245 ( .I1(n175), .I2(n176), .O(n4833) );
  NAND_GATE U246 ( .I1(n155), .I2(donnee[10]), .O(n176) );
  NAND_GATE U247 ( .I1(\registres[29][10] ), .I2(n156), .O(n175) );
  NAND_GATE U248 ( .I1(n177), .I2(n178), .O(n4834) );
  NAND_GATE U249 ( .I1(n155), .I2(donnee[11]), .O(n178) );
  NAND_GATE U250 ( .I1(\registres[29][11] ), .I2(n156), .O(n177) );
  NAND_GATE U251 ( .I1(n179), .I2(n180), .O(n4835) );
  NAND_GATE U252 ( .I1(n155), .I2(donnee[12]), .O(n180) );
  NAND_GATE U253 ( .I1(\registres[29][12] ), .I2(n156), .O(n179) );
  NAND_GATE U254 ( .I1(n181), .I2(n182), .O(n4836) );
  NAND_GATE U255 ( .I1(n155), .I2(donnee[13]), .O(n182) );
  NAND_GATE U256 ( .I1(\registres[29][13] ), .I2(n156), .O(n181) );
  NAND_GATE U257 ( .I1(n183), .I2(n184), .O(n4837) );
  NAND_GATE U258 ( .I1(n155), .I2(donnee[14]), .O(n184) );
  NAND_GATE U259 ( .I1(\registres[29][14] ), .I2(n156), .O(n183) );
  NAND_GATE U260 ( .I1(n185), .I2(n186), .O(n4838) );
  NAND_GATE U261 ( .I1(n155), .I2(donnee[15]), .O(n186) );
  NAND_GATE U262 ( .I1(\registres[29][15] ), .I2(n156), .O(n185) );
  NAND_GATE U263 ( .I1(n187), .I2(n188), .O(n4839) );
  NAND_GATE U264 ( .I1(n155), .I2(donnee[16]), .O(n188) );
  NAND_GATE U265 ( .I1(\registres[29][16] ), .I2(n156), .O(n187) );
  NAND_GATE U266 ( .I1(n189), .I2(n190), .O(n4840) );
  NAND_GATE U267 ( .I1(n155), .I2(donnee[17]), .O(n190) );
  NAND_GATE U268 ( .I1(\registres[29][17] ), .I2(n156), .O(n189) );
  NAND_GATE U269 ( .I1(n191), .I2(n192), .O(n4841) );
  NAND_GATE U270 ( .I1(n155), .I2(donnee[18]), .O(n192) );
  NAND_GATE U271 ( .I1(\registres[29][18] ), .I2(n156), .O(n191) );
  NAND_GATE U272 ( .I1(n193), .I2(n194), .O(n4842) );
  NAND_GATE U273 ( .I1(n155), .I2(donnee[19]), .O(n194) );
  NAND_GATE U274 ( .I1(\registres[29][19] ), .I2(n156), .O(n193) );
  NAND_GATE U275 ( .I1(n195), .I2(n196), .O(n4843) );
  NAND_GATE U276 ( .I1(n155), .I2(donnee[20]), .O(n196) );
  NAND_GATE U277 ( .I1(\registres[29][20] ), .I2(n156), .O(n195) );
  NAND_GATE U278 ( .I1(n197), .I2(n198), .O(n4844) );
  NAND_GATE U279 ( .I1(n155), .I2(donnee[21]), .O(n198) );
  NAND_GATE U280 ( .I1(\registres[29][21] ), .I2(n156), .O(n197) );
  NAND_GATE U281 ( .I1(n199), .I2(n200), .O(n4845) );
  NAND_GATE U282 ( .I1(n155), .I2(donnee[22]), .O(n200) );
  NAND_GATE U283 ( .I1(\registres[29][22] ), .I2(n156), .O(n199) );
  NAND_GATE U284 ( .I1(n201), .I2(n202), .O(n4846) );
  NAND_GATE U285 ( .I1(n155), .I2(donnee[23]), .O(n202) );
  NAND_GATE U286 ( .I1(\registres[29][23] ), .I2(n156), .O(n201) );
  NAND_GATE U287 ( .I1(n203), .I2(n204), .O(n4847) );
  NAND_GATE U288 ( .I1(n155), .I2(donnee[24]), .O(n204) );
  NAND_GATE U289 ( .I1(\registres[29][24] ), .I2(n156), .O(n203) );
  NAND_GATE U290 ( .I1(n205), .I2(n206), .O(n4848) );
  NAND_GATE U291 ( .I1(n155), .I2(donnee[25]), .O(n206) );
  NAND_GATE U292 ( .I1(\registres[29][25] ), .I2(n156), .O(n205) );
  NAND_GATE U293 ( .I1(n207), .I2(n208), .O(n4849) );
  NAND_GATE U294 ( .I1(n155), .I2(donnee[26]), .O(n208) );
  NAND_GATE U295 ( .I1(\registres[29][26] ), .I2(n156), .O(n207) );
  NAND_GATE U296 ( .I1(n209), .I2(n210), .O(n4850) );
  NAND_GATE U297 ( .I1(n155), .I2(donnee[27]), .O(n210) );
  NAND_GATE U298 ( .I1(\registres[29][27] ), .I2(n156), .O(n209) );
  NAND_GATE U299 ( .I1(n211), .I2(n212), .O(n4851) );
  NAND_GATE U300 ( .I1(n155), .I2(donnee[28]), .O(n212) );
  NAND_GATE U301 ( .I1(\registres[29][28] ), .I2(n156), .O(n211) );
  NAND_GATE U302 ( .I1(n213), .I2(n214), .O(n4852) );
  NAND_GATE U303 ( .I1(n155), .I2(donnee[29]), .O(n214) );
  NAND_GATE U304 ( .I1(\registres[29][29] ), .I2(n156), .O(n213) );
  NAND_GATE U305 ( .I1(n215), .I2(n216), .O(n4853) );
  NAND_GATE U306 ( .I1(n155), .I2(donnee[30]), .O(n216) );
  NAND_GATE U307 ( .I1(\registres[29][30] ), .I2(n156), .O(n215) );
  NAND_GATE U308 ( .I1(n217), .I2(n218), .O(n4854) );
  NAND_GATE U309 ( .I1(n155), .I2(donnee[31]), .O(n218) );
  AND_GATE U310 ( .I1(n219), .I2(n1), .O(n155) );
  NAND_GATE U311 ( .I1(\registres[29][31] ), .I2(n156), .O(n217) );
  NOR_GATE U312 ( .I1(n219), .I2(reset), .O(n156) );
  AND3_GATE U313 ( .I1(n83), .I2(cmd_ecr), .I3(n220), .O(n219) );
  NAND_GATE U314 ( .I1(n221), .I2(n222), .O(n4855) );
  NAND_GATE U315 ( .I1(n223), .I2(donnee[0]), .O(n222) );
  NAND_GATE U316 ( .I1(\registres[28][0] ), .I2(n224), .O(n221) );
  NAND_GATE U317 ( .I1(n225), .I2(n226), .O(n4856) );
  NAND_GATE U318 ( .I1(n223), .I2(donnee[1]), .O(n226) );
  NAND_GATE U319 ( .I1(\registres[28][1] ), .I2(n224), .O(n225) );
  NAND_GATE U320 ( .I1(n227), .I2(n228), .O(n4857) );
  NAND_GATE U321 ( .I1(n223), .I2(donnee[2]), .O(n228) );
  NAND_GATE U322 ( .I1(\registres[28][2] ), .I2(n224), .O(n227) );
  NAND_GATE U323 ( .I1(n229), .I2(n230), .O(n4858) );
  NAND_GATE U324 ( .I1(n223), .I2(donnee[3]), .O(n230) );
  NAND_GATE U325 ( .I1(\registres[28][3] ), .I2(n224), .O(n229) );
  NAND_GATE U326 ( .I1(n231), .I2(n232), .O(n4859) );
  NAND_GATE U327 ( .I1(n223), .I2(donnee[4]), .O(n232) );
  NAND_GATE U328 ( .I1(\registres[28][4] ), .I2(n224), .O(n231) );
  NAND_GATE U329 ( .I1(n233), .I2(n234), .O(n4860) );
  NAND_GATE U330 ( .I1(n223), .I2(donnee[5]), .O(n234) );
  NAND_GATE U331 ( .I1(\registres[28][5] ), .I2(n224), .O(n233) );
  NAND_GATE U332 ( .I1(n235), .I2(n236), .O(n4861) );
  NAND_GATE U333 ( .I1(n223), .I2(donnee[6]), .O(n236) );
  NAND_GATE U334 ( .I1(\registres[28][6] ), .I2(n224), .O(n235) );
  NAND_GATE U335 ( .I1(n237), .I2(n238), .O(n4862) );
  NAND_GATE U336 ( .I1(n223), .I2(donnee[7]), .O(n238) );
  NAND_GATE U337 ( .I1(\registres[28][7] ), .I2(n224), .O(n237) );
  NAND_GATE U338 ( .I1(n239), .I2(n240), .O(n4863) );
  NAND_GATE U339 ( .I1(n223), .I2(donnee[8]), .O(n240) );
  NAND_GATE U340 ( .I1(\registres[28][8] ), .I2(n224), .O(n239) );
  NAND_GATE U341 ( .I1(n241), .I2(n242), .O(n4864) );
  NAND_GATE U342 ( .I1(n223), .I2(donnee[9]), .O(n242) );
  NAND_GATE U343 ( .I1(\registres[28][9] ), .I2(n224), .O(n241) );
  NAND_GATE U344 ( .I1(n243), .I2(n244), .O(n4865) );
  NAND_GATE U345 ( .I1(n223), .I2(donnee[10]), .O(n244) );
  NAND_GATE U346 ( .I1(\registres[28][10] ), .I2(n224), .O(n243) );
  NAND_GATE U347 ( .I1(n245), .I2(n246), .O(n4866) );
  NAND_GATE U348 ( .I1(n223), .I2(donnee[11]), .O(n246) );
  NAND_GATE U349 ( .I1(\registres[28][11] ), .I2(n224), .O(n245) );
  NAND_GATE U350 ( .I1(n247), .I2(n248), .O(n4867) );
  NAND_GATE U351 ( .I1(n223), .I2(donnee[12]), .O(n248) );
  NAND_GATE U352 ( .I1(\registres[28][12] ), .I2(n224), .O(n247) );
  NAND_GATE U353 ( .I1(n249), .I2(n250), .O(n4868) );
  NAND_GATE U354 ( .I1(n223), .I2(donnee[13]), .O(n250) );
  NAND_GATE U355 ( .I1(\registres[28][13] ), .I2(n224), .O(n249) );
  NAND_GATE U356 ( .I1(n251), .I2(n252), .O(n4869) );
  NAND_GATE U357 ( .I1(n223), .I2(donnee[14]), .O(n252) );
  NAND_GATE U358 ( .I1(\registres[28][14] ), .I2(n224), .O(n251) );
  NAND_GATE U359 ( .I1(n253), .I2(n254), .O(n4870) );
  NAND_GATE U360 ( .I1(n223), .I2(donnee[15]), .O(n254) );
  NAND_GATE U361 ( .I1(\registres[28][15] ), .I2(n224), .O(n253) );
  NAND_GATE U362 ( .I1(n255), .I2(n256), .O(n4871) );
  NAND_GATE U363 ( .I1(n223), .I2(donnee[16]), .O(n256) );
  NAND_GATE U364 ( .I1(\registres[28][16] ), .I2(n224), .O(n255) );
  NAND_GATE U365 ( .I1(n257), .I2(n258), .O(n4872) );
  NAND_GATE U366 ( .I1(n223), .I2(donnee[17]), .O(n258) );
  NAND_GATE U367 ( .I1(\registres[28][17] ), .I2(n224), .O(n257) );
  NAND_GATE U368 ( .I1(n259), .I2(n260), .O(n4873) );
  NAND_GATE U369 ( .I1(n223), .I2(donnee[18]), .O(n260) );
  NAND_GATE U370 ( .I1(\registres[28][18] ), .I2(n224), .O(n259) );
  NAND_GATE U371 ( .I1(n261), .I2(n262), .O(n4874) );
  NAND_GATE U372 ( .I1(n223), .I2(donnee[19]), .O(n262) );
  NAND_GATE U373 ( .I1(\registres[28][19] ), .I2(n224), .O(n261) );
  NAND_GATE U374 ( .I1(n263), .I2(n264), .O(n4875) );
  NAND_GATE U375 ( .I1(n223), .I2(donnee[20]), .O(n264) );
  NAND_GATE U376 ( .I1(\registres[28][20] ), .I2(n224), .O(n263) );
  NAND_GATE U377 ( .I1(n265), .I2(n266), .O(n4876) );
  NAND_GATE U378 ( .I1(n223), .I2(donnee[21]), .O(n266) );
  NAND_GATE U379 ( .I1(\registres[28][21] ), .I2(n224), .O(n265) );
  NAND_GATE U380 ( .I1(n267), .I2(n268), .O(n4877) );
  NAND_GATE U381 ( .I1(n223), .I2(donnee[22]), .O(n268) );
  NAND_GATE U382 ( .I1(\registres[28][22] ), .I2(n224), .O(n267) );
  NAND_GATE U383 ( .I1(n269), .I2(n270), .O(n4878) );
  NAND_GATE U384 ( .I1(n223), .I2(donnee[23]), .O(n270) );
  NAND_GATE U385 ( .I1(\registres[28][23] ), .I2(n224), .O(n269) );
  NAND_GATE U386 ( .I1(n271), .I2(n272), .O(n4879) );
  NAND_GATE U387 ( .I1(n223), .I2(donnee[24]), .O(n272) );
  NAND_GATE U388 ( .I1(\registres[28][24] ), .I2(n224), .O(n271) );
  NAND_GATE U389 ( .I1(n273), .I2(n274), .O(n4880) );
  NAND_GATE U390 ( .I1(n223), .I2(donnee[25]), .O(n274) );
  NAND_GATE U391 ( .I1(\registres[28][25] ), .I2(n224), .O(n273) );
  NAND_GATE U392 ( .I1(n275), .I2(n276), .O(n4881) );
  NAND_GATE U393 ( .I1(n223), .I2(donnee[26]), .O(n276) );
  NAND_GATE U394 ( .I1(\registres[28][26] ), .I2(n224), .O(n275) );
  NAND_GATE U395 ( .I1(n277), .I2(n278), .O(n4882) );
  NAND_GATE U396 ( .I1(n223), .I2(donnee[27]), .O(n278) );
  NAND_GATE U397 ( .I1(\registres[28][27] ), .I2(n224), .O(n277) );
  NAND_GATE U398 ( .I1(n279), .I2(n280), .O(n4883) );
  NAND_GATE U399 ( .I1(n223), .I2(donnee[28]), .O(n280) );
  NAND_GATE U400 ( .I1(\registres[28][28] ), .I2(n224), .O(n279) );
  NAND_GATE U401 ( .I1(n281), .I2(n282), .O(n4884) );
  NAND_GATE U402 ( .I1(n223), .I2(donnee[29]), .O(n282) );
  NAND_GATE U403 ( .I1(\registres[28][29] ), .I2(n224), .O(n281) );
  NAND_GATE U404 ( .I1(n283), .I2(n284), .O(n4885) );
  NAND_GATE U405 ( .I1(n223), .I2(donnee[30]), .O(n284) );
  NAND_GATE U406 ( .I1(\registres[28][30] ), .I2(n224), .O(n283) );
  NAND_GATE U407 ( .I1(n285), .I2(n286), .O(n4886) );
  NAND_GATE U408 ( .I1(n223), .I2(donnee[31]), .O(n286) );
  AND_GATE U409 ( .I1(n287), .I2(n1), .O(n223) );
  NAND_GATE U410 ( .I1(\registres[28][31] ), .I2(n224), .O(n285) );
  NOR_GATE U411 ( .I1(n287), .I2(reset), .O(n224) );
  AND3_GATE U412 ( .I1(n83), .I2(cmd_ecr), .I3(n288), .O(n287) );
  NAND_GATE U413 ( .I1(n289), .I2(n290), .O(n4887) );
  NAND_GATE U414 ( .I1(n291), .I2(donnee[0]), .O(n290) );
  NAND_GATE U415 ( .I1(\registres[27][0] ), .I2(n292), .O(n289) );
  NAND_GATE U416 ( .I1(n293), .I2(n294), .O(n4888) );
  NAND_GATE U417 ( .I1(n291), .I2(donnee[1]), .O(n294) );
  NAND_GATE U418 ( .I1(\registres[27][1] ), .I2(n292), .O(n293) );
  NAND_GATE U419 ( .I1(n295), .I2(n296), .O(n4889) );
  NAND_GATE U420 ( .I1(n291), .I2(donnee[2]), .O(n296) );
  NAND_GATE U421 ( .I1(\registres[27][2] ), .I2(n292), .O(n295) );
  NAND_GATE U422 ( .I1(n297), .I2(n298), .O(n4890) );
  NAND_GATE U423 ( .I1(n291), .I2(donnee[3]), .O(n298) );
  NAND_GATE U424 ( .I1(\registres[27][3] ), .I2(n292), .O(n297) );
  NAND_GATE U425 ( .I1(n299), .I2(n300), .O(n4891) );
  NAND_GATE U426 ( .I1(n291), .I2(donnee[4]), .O(n300) );
  NAND_GATE U427 ( .I1(\registres[27][4] ), .I2(n292), .O(n299) );
  NAND_GATE U428 ( .I1(n301), .I2(n302), .O(n4892) );
  NAND_GATE U429 ( .I1(n291), .I2(donnee[5]), .O(n302) );
  NAND_GATE U430 ( .I1(\registres[27][5] ), .I2(n292), .O(n301) );
  NAND_GATE U431 ( .I1(n303), .I2(n304), .O(n4893) );
  NAND_GATE U432 ( .I1(n291), .I2(donnee[6]), .O(n304) );
  NAND_GATE U433 ( .I1(\registres[27][6] ), .I2(n292), .O(n303) );
  NAND_GATE U434 ( .I1(n305), .I2(n306), .O(n4894) );
  NAND_GATE U435 ( .I1(n291), .I2(donnee[7]), .O(n306) );
  NAND_GATE U436 ( .I1(\registres[27][7] ), .I2(n292), .O(n305) );
  NAND_GATE U437 ( .I1(n307), .I2(n308), .O(n4895) );
  NAND_GATE U438 ( .I1(n291), .I2(donnee[8]), .O(n308) );
  NAND_GATE U439 ( .I1(\registres[27][8] ), .I2(n292), .O(n307) );
  NAND_GATE U440 ( .I1(n309), .I2(n310), .O(n4896) );
  NAND_GATE U441 ( .I1(n291), .I2(donnee[9]), .O(n310) );
  NAND_GATE U442 ( .I1(\registres[27][9] ), .I2(n292), .O(n309) );
  NAND_GATE U443 ( .I1(n311), .I2(n312), .O(n4897) );
  NAND_GATE U444 ( .I1(n291), .I2(donnee[10]), .O(n312) );
  NAND_GATE U445 ( .I1(\registres[27][10] ), .I2(n292), .O(n311) );
  NAND_GATE U446 ( .I1(n313), .I2(n314), .O(n4898) );
  NAND_GATE U447 ( .I1(n291), .I2(donnee[11]), .O(n314) );
  NAND_GATE U448 ( .I1(\registres[27][11] ), .I2(n292), .O(n313) );
  NAND_GATE U449 ( .I1(n315), .I2(n316), .O(n4899) );
  NAND_GATE U450 ( .I1(n291), .I2(donnee[12]), .O(n316) );
  NAND_GATE U451 ( .I1(\registres[27][12] ), .I2(n292), .O(n315) );
  NAND_GATE U452 ( .I1(n317), .I2(n318), .O(n4900) );
  NAND_GATE U453 ( .I1(n291), .I2(donnee[13]), .O(n318) );
  NAND_GATE U454 ( .I1(\registres[27][13] ), .I2(n292), .O(n317) );
  NAND_GATE U455 ( .I1(n319), .I2(n320), .O(n4901) );
  NAND_GATE U456 ( .I1(n291), .I2(donnee[14]), .O(n320) );
  NAND_GATE U457 ( .I1(\registres[27][14] ), .I2(n292), .O(n319) );
  NAND_GATE U458 ( .I1(n321), .I2(n322), .O(n4902) );
  NAND_GATE U459 ( .I1(n291), .I2(donnee[15]), .O(n322) );
  NAND_GATE U460 ( .I1(\registres[27][15] ), .I2(n292), .O(n321) );
  NAND_GATE U461 ( .I1(n323), .I2(n324), .O(n4903) );
  NAND_GATE U462 ( .I1(n291), .I2(donnee[16]), .O(n324) );
  NAND_GATE U463 ( .I1(\registres[27][16] ), .I2(n292), .O(n323) );
  NAND_GATE U464 ( .I1(n325), .I2(n326), .O(n4904) );
  NAND_GATE U465 ( .I1(n291), .I2(donnee[17]), .O(n326) );
  NAND_GATE U466 ( .I1(\registres[27][17] ), .I2(n292), .O(n325) );
  NAND_GATE U467 ( .I1(n327), .I2(n328), .O(n4905) );
  NAND_GATE U468 ( .I1(n291), .I2(donnee[18]), .O(n328) );
  NAND_GATE U469 ( .I1(\registres[27][18] ), .I2(n292), .O(n327) );
  NAND_GATE U470 ( .I1(n329), .I2(n330), .O(n4906) );
  NAND_GATE U471 ( .I1(n291), .I2(donnee[19]), .O(n330) );
  NAND_GATE U472 ( .I1(\registres[27][19] ), .I2(n292), .O(n329) );
  NAND_GATE U473 ( .I1(n331), .I2(n332), .O(n4907) );
  NAND_GATE U474 ( .I1(n291), .I2(donnee[20]), .O(n332) );
  NAND_GATE U475 ( .I1(\registres[27][20] ), .I2(n292), .O(n331) );
  NAND_GATE U476 ( .I1(n333), .I2(n334), .O(n4908) );
  NAND_GATE U477 ( .I1(n291), .I2(donnee[21]), .O(n334) );
  NAND_GATE U478 ( .I1(\registres[27][21] ), .I2(n292), .O(n333) );
  NAND_GATE U479 ( .I1(n335), .I2(n336), .O(n4909) );
  NAND_GATE U480 ( .I1(n291), .I2(donnee[22]), .O(n336) );
  NAND_GATE U481 ( .I1(\registres[27][22] ), .I2(n292), .O(n335) );
  NAND_GATE U482 ( .I1(n337), .I2(n338), .O(n4910) );
  NAND_GATE U483 ( .I1(n291), .I2(donnee[23]), .O(n338) );
  NAND_GATE U484 ( .I1(\registres[27][23] ), .I2(n292), .O(n337) );
  NAND_GATE U485 ( .I1(n339), .I2(n340), .O(n4911) );
  NAND_GATE U486 ( .I1(n291), .I2(donnee[24]), .O(n340) );
  NAND_GATE U487 ( .I1(\registres[27][24] ), .I2(n292), .O(n339) );
  NAND_GATE U488 ( .I1(n341), .I2(n342), .O(n4912) );
  NAND_GATE U489 ( .I1(n291), .I2(donnee[25]), .O(n342) );
  NAND_GATE U490 ( .I1(\registres[27][25] ), .I2(n292), .O(n341) );
  NAND_GATE U491 ( .I1(n343), .I2(n344), .O(n4913) );
  NAND_GATE U492 ( .I1(n291), .I2(donnee[26]), .O(n344) );
  NAND_GATE U493 ( .I1(\registres[27][26] ), .I2(n292), .O(n343) );
  NAND_GATE U494 ( .I1(n345), .I2(n346), .O(n4914) );
  NAND_GATE U495 ( .I1(n291), .I2(donnee[27]), .O(n346) );
  NAND_GATE U496 ( .I1(\registres[27][27] ), .I2(n292), .O(n345) );
  NAND_GATE U497 ( .I1(n347), .I2(n348), .O(n4915) );
  NAND_GATE U498 ( .I1(n291), .I2(donnee[28]), .O(n348) );
  NAND_GATE U499 ( .I1(\registres[27][28] ), .I2(n292), .O(n347) );
  NAND_GATE U500 ( .I1(n349), .I2(n350), .O(n4916) );
  NAND_GATE U501 ( .I1(n291), .I2(donnee[29]), .O(n350) );
  NAND_GATE U502 ( .I1(\registres[27][29] ), .I2(n292), .O(n349) );
  NAND_GATE U503 ( .I1(n351), .I2(n352), .O(n4917) );
  NAND_GATE U504 ( .I1(n291), .I2(donnee[30]), .O(n352) );
  NAND_GATE U505 ( .I1(\registres[27][30] ), .I2(n292), .O(n351) );
  NAND_GATE U506 ( .I1(n353), .I2(n354), .O(n4918) );
  NAND_GATE U507 ( .I1(n291), .I2(donnee[31]), .O(n354) );
  AND_GATE U508 ( .I1(n355), .I2(n1), .O(n291) );
  NAND_GATE U509 ( .I1(\registres[27][31] ), .I2(n292), .O(n353) );
  NOR_GATE U510 ( .I1(n355), .I2(reset), .O(n292) );
  AND3_GATE U511 ( .I1(n83), .I2(cmd_ecr), .I3(n356), .O(n355) );
  NAND_GATE U512 ( .I1(n357), .I2(n358), .O(n4919) );
  NAND_GATE U513 ( .I1(n359), .I2(donnee[0]), .O(n358) );
  NAND_GATE U514 ( .I1(\registres[26][0] ), .I2(n360), .O(n357) );
  NAND_GATE U515 ( .I1(n361), .I2(n362), .O(n4920) );
  NAND_GATE U516 ( .I1(n359), .I2(donnee[1]), .O(n362) );
  NAND_GATE U517 ( .I1(\registres[26][1] ), .I2(n360), .O(n361) );
  NAND_GATE U518 ( .I1(n363), .I2(n364), .O(n4921) );
  NAND_GATE U519 ( .I1(n359), .I2(donnee[2]), .O(n364) );
  NAND_GATE U520 ( .I1(\registres[26][2] ), .I2(n360), .O(n363) );
  NAND_GATE U521 ( .I1(n365), .I2(n366), .O(n4922) );
  NAND_GATE U522 ( .I1(n359), .I2(donnee[3]), .O(n366) );
  NAND_GATE U523 ( .I1(\registres[26][3] ), .I2(n360), .O(n365) );
  NAND_GATE U524 ( .I1(n367), .I2(n368), .O(n4923) );
  NAND_GATE U525 ( .I1(n359), .I2(donnee[4]), .O(n368) );
  NAND_GATE U526 ( .I1(\registres[26][4] ), .I2(n360), .O(n367) );
  NAND_GATE U527 ( .I1(n369), .I2(n370), .O(n4924) );
  NAND_GATE U528 ( .I1(n359), .I2(donnee[5]), .O(n370) );
  NAND_GATE U529 ( .I1(\registres[26][5] ), .I2(n360), .O(n369) );
  NAND_GATE U530 ( .I1(n371), .I2(n372), .O(n4925) );
  NAND_GATE U531 ( .I1(n359), .I2(donnee[6]), .O(n372) );
  NAND_GATE U532 ( .I1(\registres[26][6] ), .I2(n360), .O(n371) );
  NAND_GATE U533 ( .I1(n373), .I2(n374), .O(n4926) );
  NAND_GATE U534 ( .I1(n359), .I2(donnee[7]), .O(n374) );
  NAND_GATE U535 ( .I1(\registres[26][7] ), .I2(n360), .O(n373) );
  NAND_GATE U536 ( .I1(n375), .I2(n376), .O(n4927) );
  NAND_GATE U537 ( .I1(n359), .I2(donnee[8]), .O(n376) );
  NAND_GATE U538 ( .I1(\registres[26][8] ), .I2(n360), .O(n375) );
  NAND_GATE U539 ( .I1(n377), .I2(n378), .O(n4928) );
  NAND_GATE U540 ( .I1(n359), .I2(donnee[9]), .O(n378) );
  NAND_GATE U541 ( .I1(\registres[26][9] ), .I2(n360), .O(n377) );
  NAND_GATE U542 ( .I1(n379), .I2(n380), .O(n4929) );
  NAND_GATE U543 ( .I1(n359), .I2(donnee[10]), .O(n380) );
  NAND_GATE U544 ( .I1(\registres[26][10] ), .I2(n360), .O(n379) );
  NAND_GATE U545 ( .I1(n381), .I2(n382), .O(n4930) );
  NAND_GATE U546 ( .I1(n359), .I2(donnee[11]), .O(n382) );
  NAND_GATE U547 ( .I1(\registres[26][11] ), .I2(n360), .O(n381) );
  NAND_GATE U548 ( .I1(n383), .I2(n384), .O(n4931) );
  NAND_GATE U549 ( .I1(n359), .I2(donnee[12]), .O(n384) );
  NAND_GATE U550 ( .I1(\registres[26][12] ), .I2(n360), .O(n383) );
  NAND_GATE U551 ( .I1(n385), .I2(n386), .O(n4932) );
  NAND_GATE U552 ( .I1(n359), .I2(donnee[13]), .O(n386) );
  NAND_GATE U553 ( .I1(\registres[26][13] ), .I2(n360), .O(n385) );
  NAND_GATE U554 ( .I1(n387), .I2(n388), .O(n4933) );
  NAND_GATE U555 ( .I1(n359), .I2(donnee[14]), .O(n388) );
  NAND_GATE U556 ( .I1(\registres[26][14] ), .I2(n360), .O(n387) );
  NAND_GATE U557 ( .I1(n389), .I2(n390), .O(n4934) );
  NAND_GATE U558 ( .I1(n359), .I2(donnee[15]), .O(n390) );
  NAND_GATE U559 ( .I1(\registres[26][15] ), .I2(n360), .O(n389) );
  NAND_GATE U560 ( .I1(n391), .I2(n392), .O(n4935) );
  NAND_GATE U561 ( .I1(n359), .I2(donnee[16]), .O(n392) );
  NAND_GATE U562 ( .I1(\registres[26][16] ), .I2(n360), .O(n391) );
  NAND_GATE U563 ( .I1(n393), .I2(n394), .O(n4936) );
  NAND_GATE U564 ( .I1(n359), .I2(donnee[17]), .O(n394) );
  NAND_GATE U565 ( .I1(\registres[26][17] ), .I2(n360), .O(n393) );
  NAND_GATE U566 ( .I1(n395), .I2(n396), .O(n4937) );
  NAND_GATE U567 ( .I1(n359), .I2(donnee[18]), .O(n396) );
  NAND_GATE U568 ( .I1(\registres[26][18] ), .I2(n360), .O(n395) );
  NAND_GATE U569 ( .I1(n397), .I2(n398), .O(n4938) );
  NAND_GATE U570 ( .I1(n359), .I2(donnee[19]), .O(n398) );
  NAND_GATE U571 ( .I1(\registres[26][19] ), .I2(n360), .O(n397) );
  NAND_GATE U572 ( .I1(n399), .I2(n400), .O(n4939) );
  NAND_GATE U573 ( .I1(n359), .I2(donnee[20]), .O(n400) );
  NAND_GATE U574 ( .I1(\registres[26][20] ), .I2(n360), .O(n399) );
  NAND_GATE U575 ( .I1(n401), .I2(n402), .O(n4940) );
  NAND_GATE U576 ( .I1(n359), .I2(donnee[21]), .O(n402) );
  NAND_GATE U577 ( .I1(\registres[26][21] ), .I2(n360), .O(n401) );
  NAND_GATE U578 ( .I1(n403), .I2(n404), .O(n4941) );
  NAND_GATE U579 ( .I1(n359), .I2(donnee[22]), .O(n404) );
  NAND_GATE U580 ( .I1(\registres[26][22] ), .I2(n360), .O(n403) );
  NAND_GATE U581 ( .I1(n405), .I2(n406), .O(n4942) );
  NAND_GATE U582 ( .I1(n359), .I2(donnee[23]), .O(n406) );
  NAND_GATE U583 ( .I1(\registres[26][23] ), .I2(n360), .O(n405) );
  NAND_GATE U584 ( .I1(n407), .I2(n408), .O(n4943) );
  NAND_GATE U585 ( .I1(n359), .I2(donnee[24]), .O(n408) );
  NAND_GATE U586 ( .I1(\registres[26][24] ), .I2(n360), .O(n407) );
  NAND_GATE U587 ( .I1(n409), .I2(n410), .O(n4944) );
  NAND_GATE U588 ( .I1(n359), .I2(donnee[25]), .O(n410) );
  NAND_GATE U589 ( .I1(\registres[26][25] ), .I2(n360), .O(n409) );
  NAND_GATE U590 ( .I1(n411), .I2(n412), .O(n4945) );
  NAND_GATE U591 ( .I1(n359), .I2(donnee[26]), .O(n412) );
  NAND_GATE U592 ( .I1(\registres[26][26] ), .I2(n360), .O(n411) );
  NAND_GATE U593 ( .I1(n413), .I2(n414), .O(n4946) );
  NAND_GATE U594 ( .I1(n359), .I2(donnee[27]), .O(n414) );
  NAND_GATE U595 ( .I1(\registres[26][27] ), .I2(n360), .O(n413) );
  NAND_GATE U596 ( .I1(n415), .I2(n416), .O(n4947) );
  NAND_GATE U597 ( .I1(n359), .I2(donnee[28]), .O(n416) );
  NAND_GATE U598 ( .I1(\registres[26][28] ), .I2(n360), .O(n415) );
  NAND_GATE U599 ( .I1(n417), .I2(n418), .O(n4948) );
  NAND_GATE U600 ( .I1(n359), .I2(donnee[29]), .O(n418) );
  NAND_GATE U601 ( .I1(\registres[26][29] ), .I2(n360), .O(n417) );
  NAND_GATE U602 ( .I1(n419), .I2(n420), .O(n4949) );
  NAND_GATE U603 ( .I1(n359), .I2(donnee[30]), .O(n420) );
  NAND_GATE U604 ( .I1(\registres[26][30] ), .I2(n360), .O(n419) );
  NAND_GATE U605 ( .I1(n421), .I2(n422), .O(n4950) );
  NAND_GATE U606 ( .I1(n359), .I2(donnee[31]), .O(n422) );
  AND_GATE U607 ( .I1(n423), .I2(n1), .O(n359) );
  NAND_GATE U608 ( .I1(\registres[26][31] ), .I2(n360), .O(n421) );
  NOR_GATE U609 ( .I1(n423), .I2(reset), .O(n360) );
  AND3_GATE U610 ( .I1(n83), .I2(cmd_ecr), .I3(n424), .O(n423) );
  NAND_GATE U611 ( .I1(n425), .I2(n426), .O(n4951) );
  NAND_GATE U612 ( .I1(n427), .I2(donnee[0]), .O(n426) );
  NAND_GATE U613 ( .I1(\registres[25][0] ), .I2(n428), .O(n425) );
  NAND_GATE U614 ( .I1(n429), .I2(n430), .O(n4952) );
  NAND_GATE U615 ( .I1(n427), .I2(donnee[1]), .O(n430) );
  NAND_GATE U616 ( .I1(\registres[25][1] ), .I2(n428), .O(n429) );
  NAND_GATE U617 ( .I1(n431), .I2(n432), .O(n4953) );
  NAND_GATE U618 ( .I1(n427), .I2(donnee[2]), .O(n432) );
  NAND_GATE U619 ( .I1(\registres[25][2] ), .I2(n428), .O(n431) );
  NAND_GATE U620 ( .I1(n433), .I2(n434), .O(n4954) );
  NAND_GATE U621 ( .I1(n427), .I2(donnee[3]), .O(n434) );
  NAND_GATE U622 ( .I1(\registres[25][3] ), .I2(n428), .O(n433) );
  NAND_GATE U623 ( .I1(n435), .I2(n436), .O(n4955) );
  NAND_GATE U624 ( .I1(n427), .I2(donnee[4]), .O(n436) );
  NAND_GATE U625 ( .I1(\registres[25][4] ), .I2(n428), .O(n435) );
  NAND_GATE U626 ( .I1(n437), .I2(n438), .O(n4956) );
  NAND_GATE U627 ( .I1(n427), .I2(donnee[5]), .O(n438) );
  NAND_GATE U628 ( .I1(\registres[25][5] ), .I2(n428), .O(n437) );
  NAND_GATE U629 ( .I1(n439), .I2(n440), .O(n4957) );
  NAND_GATE U630 ( .I1(n427), .I2(donnee[6]), .O(n440) );
  NAND_GATE U631 ( .I1(\registres[25][6] ), .I2(n428), .O(n439) );
  NAND_GATE U632 ( .I1(n441), .I2(n442), .O(n4958) );
  NAND_GATE U633 ( .I1(n427), .I2(donnee[7]), .O(n442) );
  NAND_GATE U634 ( .I1(\registres[25][7] ), .I2(n428), .O(n441) );
  NAND_GATE U635 ( .I1(n443), .I2(n444), .O(n4959) );
  NAND_GATE U636 ( .I1(n427), .I2(donnee[8]), .O(n444) );
  NAND_GATE U637 ( .I1(\registres[25][8] ), .I2(n428), .O(n443) );
  NAND_GATE U638 ( .I1(n445), .I2(n446), .O(n4960) );
  NAND_GATE U639 ( .I1(n427), .I2(donnee[9]), .O(n446) );
  NAND_GATE U640 ( .I1(\registres[25][9] ), .I2(n428), .O(n445) );
  NAND_GATE U641 ( .I1(n447), .I2(n448), .O(n4961) );
  NAND_GATE U642 ( .I1(n427), .I2(donnee[10]), .O(n448) );
  NAND_GATE U643 ( .I1(\registres[25][10] ), .I2(n428), .O(n447) );
  NAND_GATE U644 ( .I1(n449), .I2(n450), .O(n4962) );
  NAND_GATE U645 ( .I1(n427), .I2(donnee[11]), .O(n450) );
  NAND_GATE U646 ( .I1(\registres[25][11] ), .I2(n428), .O(n449) );
  NAND_GATE U647 ( .I1(n451), .I2(n452), .O(n4963) );
  NAND_GATE U648 ( .I1(n427), .I2(donnee[12]), .O(n452) );
  NAND_GATE U649 ( .I1(\registres[25][12] ), .I2(n428), .O(n451) );
  NAND_GATE U650 ( .I1(n453), .I2(n454), .O(n4964) );
  NAND_GATE U651 ( .I1(n427), .I2(donnee[13]), .O(n454) );
  NAND_GATE U652 ( .I1(\registres[25][13] ), .I2(n428), .O(n453) );
  NAND_GATE U653 ( .I1(n455), .I2(n456), .O(n4965) );
  NAND_GATE U654 ( .I1(n427), .I2(donnee[14]), .O(n456) );
  NAND_GATE U655 ( .I1(\registres[25][14] ), .I2(n428), .O(n455) );
  NAND_GATE U656 ( .I1(n457), .I2(n458), .O(n4966) );
  NAND_GATE U657 ( .I1(n427), .I2(donnee[15]), .O(n458) );
  NAND_GATE U658 ( .I1(\registres[25][15] ), .I2(n428), .O(n457) );
  NAND_GATE U659 ( .I1(n459), .I2(n460), .O(n4967) );
  NAND_GATE U660 ( .I1(n427), .I2(donnee[16]), .O(n460) );
  NAND_GATE U661 ( .I1(\registres[25][16] ), .I2(n428), .O(n459) );
  NAND_GATE U662 ( .I1(n461), .I2(n462), .O(n4968) );
  NAND_GATE U663 ( .I1(n427), .I2(donnee[17]), .O(n462) );
  NAND_GATE U664 ( .I1(\registres[25][17] ), .I2(n428), .O(n461) );
  NAND_GATE U665 ( .I1(n463), .I2(n464), .O(n4969) );
  NAND_GATE U666 ( .I1(n427), .I2(donnee[18]), .O(n464) );
  NAND_GATE U667 ( .I1(\registres[25][18] ), .I2(n428), .O(n463) );
  NAND_GATE U668 ( .I1(n465), .I2(n466), .O(n4970) );
  NAND_GATE U669 ( .I1(n427), .I2(donnee[19]), .O(n466) );
  NAND_GATE U670 ( .I1(\registres[25][19] ), .I2(n428), .O(n465) );
  NAND_GATE U671 ( .I1(n467), .I2(n468), .O(n4971) );
  NAND_GATE U672 ( .I1(n427), .I2(donnee[20]), .O(n468) );
  NAND_GATE U673 ( .I1(\registres[25][20] ), .I2(n428), .O(n467) );
  NAND_GATE U674 ( .I1(n469), .I2(n470), .O(n4972) );
  NAND_GATE U675 ( .I1(n427), .I2(donnee[21]), .O(n470) );
  NAND_GATE U676 ( .I1(\registres[25][21] ), .I2(n428), .O(n469) );
  NAND_GATE U677 ( .I1(n471), .I2(n472), .O(n4973) );
  NAND_GATE U678 ( .I1(n427), .I2(donnee[22]), .O(n472) );
  NAND_GATE U679 ( .I1(\registres[25][22] ), .I2(n428), .O(n471) );
  NAND_GATE U680 ( .I1(n473), .I2(n474), .O(n4974) );
  NAND_GATE U681 ( .I1(n427), .I2(donnee[23]), .O(n474) );
  NAND_GATE U682 ( .I1(\registres[25][23] ), .I2(n428), .O(n473) );
  NAND_GATE U683 ( .I1(n475), .I2(n476), .O(n4975) );
  NAND_GATE U684 ( .I1(n427), .I2(donnee[24]), .O(n476) );
  NAND_GATE U685 ( .I1(\registres[25][24] ), .I2(n428), .O(n475) );
  NAND_GATE U686 ( .I1(n477), .I2(n478), .O(n4976) );
  NAND_GATE U687 ( .I1(n427), .I2(donnee[25]), .O(n478) );
  NAND_GATE U688 ( .I1(\registres[25][25] ), .I2(n428), .O(n477) );
  NAND_GATE U689 ( .I1(n479), .I2(n480), .O(n4977) );
  NAND_GATE U690 ( .I1(n427), .I2(donnee[26]), .O(n480) );
  NAND_GATE U691 ( .I1(\registres[25][26] ), .I2(n428), .O(n479) );
  NAND_GATE U692 ( .I1(n481), .I2(n482), .O(n4978) );
  NAND_GATE U693 ( .I1(n427), .I2(donnee[27]), .O(n482) );
  NAND_GATE U694 ( .I1(\registres[25][27] ), .I2(n428), .O(n481) );
  NAND_GATE U695 ( .I1(n483), .I2(n484), .O(n4979) );
  NAND_GATE U696 ( .I1(n427), .I2(donnee[28]), .O(n484) );
  NAND_GATE U697 ( .I1(\registres[25][28] ), .I2(n428), .O(n483) );
  NAND_GATE U698 ( .I1(n485), .I2(n486), .O(n4980) );
  NAND_GATE U699 ( .I1(n427), .I2(donnee[29]), .O(n486) );
  NAND_GATE U700 ( .I1(\registres[25][29] ), .I2(n428), .O(n485) );
  NAND_GATE U701 ( .I1(n487), .I2(n488), .O(n4981) );
  NAND_GATE U702 ( .I1(n427), .I2(donnee[30]), .O(n488) );
  NAND_GATE U703 ( .I1(\registres[25][30] ), .I2(n428), .O(n487) );
  NAND_GATE U704 ( .I1(n489), .I2(n490), .O(n4982) );
  NAND_GATE U705 ( .I1(n427), .I2(donnee[31]), .O(n490) );
  AND_GATE U706 ( .I1(n491), .I2(n1), .O(n427) );
  NAND_GATE U707 ( .I1(\registres[25][31] ), .I2(n428), .O(n489) );
  NOR_GATE U708 ( .I1(n491), .I2(reset), .O(n428) );
  AND3_GATE U709 ( .I1(n83), .I2(cmd_ecr), .I3(n492), .O(n491) );
  NAND_GATE U710 ( .I1(n493), .I2(n494), .O(n4983) );
  NAND_GATE U711 ( .I1(n495), .I2(donnee[0]), .O(n494) );
  NAND_GATE U712 ( .I1(\registres[24][0] ), .I2(n496), .O(n493) );
  NAND_GATE U713 ( .I1(n497), .I2(n498), .O(n4984) );
  NAND_GATE U714 ( .I1(n495), .I2(donnee[1]), .O(n498) );
  NAND_GATE U715 ( .I1(\registres[24][1] ), .I2(n496), .O(n497) );
  NAND_GATE U716 ( .I1(n499), .I2(n500), .O(n4985) );
  NAND_GATE U717 ( .I1(n495), .I2(donnee[2]), .O(n500) );
  NAND_GATE U718 ( .I1(\registres[24][2] ), .I2(n496), .O(n499) );
  NAND_GATE U719 ( .I1(n501), .I2(n502), .O(n4986) );
  NAND_GATE U720 ( .I1(n495), .I2(donnee[3]), .O(n502) );
  NAND_GATE U721 ( .I1(\registres[24][3] ), .I2(n496), .O(n501) );
  NAND_GATE U722 ( .I1(n503), .I2(n504), .O(n4987) );
  NAND_GATE U723 ( .I1(n495), .I2(donnee[4]), .O(n504) );
  NAND_GATE U724 ( .I1(\registres[24][4] ), .I2(n496), .O(n503) );
  NAND_GATE U725 ( .I1(n505), .I2(n506), .O(n4988) );
  NAND_GATE U726 ( .I1(n495), .I2(donnee[5]), .O(n506) );
  NAND_GATE U727 ( .I1(\registres[24][5] ), .I2(n496), .O(n505) );
  NAND_GATE U728 ( .I1(n507), .I2(n508), .O(n4989) );
  NAND_GATE U729 ( .I1(n495), .I2(donnee[6]), .O(n508) );
  NAND_GATE U730 ( .I1(\registres[24][6] ), .I2(n496), .O(n507) );
  NAND_GATE U731 ( .I1(n509), .I2(n510), .O(n4990) );
  NAND_GATE U732 ( .I1(n495), .I2(donnee[7]), .O(n510) );
  NAND_GATE U733 ( .I1(\registres[24][7] ), .I2(n496), .O(n509) );
  NAND_GATE U734 ( .I1(n511), .I2(n512), .O(n4991) );
  NAND_GATE U735 ( .I1(n495), .I2(donnee[8]), .O(n512) );
  NAND_GATE U736 ( .I1(\registres[24][8] ), .I2(n496), .O(n511) );
  NAND_GATE U737 ( .I1(n513), .I2(n514), .O(n4992) );
  NAND_GATE U738 ( .I1(n495), .I2(donnee[9]), .O(n514) );
  NAND_GATE U739 ( .I1(\registres[24][9] ), .I2(n496), .O(n513) );
  NAND_GATE U740 ( .I1(n515), .I2(n516), .O(n4993) );
  NAND_GATE U741 ( .I1(n495), .I2(donnee[10]), .O(n516) );
  NAND_GATE U742 ( .I1(\registres[24][10] ), .I2(n496), .O(n515) );
  NAND_GATE U743 ( .I1(n517), .I2(n518), .O(n4994) );
  NAND_GATE U744 ( .I1(n495), .I2(donnee[11]), .O(n518) );
  NAND_GATE U745 ( .I1(\registres[24][11] ), .I2(n496), .O(n517) );
  NAND_GATE U746 ( .I1(n519), .I2(n520), .O(n4995) );
  NAND_GATE U747 ( .I1(n495), .I2(donnee[12]), .O(n520) );
  NAND_GATE U748 ( .I1(\registres[24][12] ), .I2(n496), .O(n519) );
  NAND_GATE U749 ( .I1(n521), .I2(n522), .O(n4996) );
  NAND_GATE U750 ( .I1(n495), .I2(donnee[13]), .O(n522) );
  NAND_GATE U751 ( .I1(\registres[24][13] ), .I2(n496), .O(n521) );
  NAND_GATE U752 ( .I1(n523), .I2(n524), .O(n4997) );
  NAND_GATE U753 ( .I1(n495), .I2(donnee[14]), .O(n524) );
  NAND_GATE U754 ( .I1(\registres[24][14] ), .I2(n496), .O(n523) );
  NAND_GATE U755 ( .I1(n525), .I2(n526), .O(n4998) );
  NAND_GATE U756 ( .I1(n495), .I2(donnee[15]), .O(n526) );
  NAND_GATE U757 ( .I1(\registres[24][15] ), .I2(n496), .O(n525) );
  NAND_GATE U758 ( .I1(n527), .I2(n528), .O(n4999) );
  NAND_GATE U759 ( .I1(n495), .I2(donnee[16]), .O(n528) );
  NAND_GATE U760 ( .I1(\registres[24][16] ), .I2(n496), .O(n527) );
  NAND_GATE U761 ( .I1(n529), .I2(n530), .O(n5000) );
  NAND_GATE U762 ( .I1(n495), .I2(donnee[17]), .O(n530) );
  NAND_GATE U763 ( .I1(\registres[24][17] ), .I2(n496), .O(n529) );
  NAND_GATE U764 ( .I1(n531), .I2(n532), .O(n5001) );
  NAND_GATE U765 ( .I1(n495), .I2(donnee[18]), .O(n532) );
  NAND_GATE U766 ( .I1(\registres[24][18] ), .I2(n496), .O(n531) );
  NAND_GATE U767 ( .I1(n533), .I2(n534), .O(n5002) );
  NAND_GATE U768 ( .I1(n495), .I2(donnee[19]), .O(n534) );
  NAND_GATE U769 ( .I1(\registres[24][19] ), .I2(n496), .O(n533) );
  NAND_GATE U770 ( .I1(n535), .I2(n536), .O(n5003) );
  NAND_GATE U771 ( .I1(n495), .I2(donnee[20]), .O(n536) );
  NAND_GATE U772 ( .I1(\registres[24][20] ), .I2(n496), .O(n535) );
  NAND_GATE U773 ( .I1(n537), .I2(n538), .O(n5004) );
  NAND_GATE U774 ( .I1(n495), .I2(donnee[21]), .O(n538) );
  NAND_GATE U775 ( .I1(\registres[24][21] ), .I2(n496), .O(n537) );
  NAND_GATE U776 ( .I1(n539), .I2(n540), .O(n5005) );
  NAND_GATE U777 ( .I1(n495), .I2(donnee[22]), .O(n540) );
  NAND_GATE U778 ( .I1(\registres[24][22] ), .I2(n496), .O(n539) );
  NAND_GATE U779 ( .I1(n541), .I2(n542), .O(n5006) );
  NAND_GATE U780 ( .I1(n495), .I2(donnee[23]), .O(n542) );
  NAND_GATE U781 ( .I1(\registres[24][23] ), .I2(n496), .O(n541) );
  NAND_GATE U782 ( .I1(n543), .I2(n544), .O(n5007) );
  NAND_GATE U783 ( .I1(n495), .I2(donnee[24]), .O(n544) );
  NAND_GATE U784 ( .I1(\registres[24][24] ), .I2(n496), .O(n543) );
  NAND_GATE U785 ( .I1(n545), .I2(n546), .O(n5008) );
  NAND_GATE U786 ( .I1(n495), .I2(donnee[25]), .O(n546) );
  NAND_GATE U787 ( .I1(\registres[24][25] ), .I2(n496), .O(n545) );
  NAND_GATE U788 ( .I1(n547), .I2(n548), .O(n5009) );
  NAND_GATE U789 ( .I1(n495), .I2(donnee[26]), .O(n548) );
  NAND_GATE U790 ( .I1(\registres[24][26] ), .I2(n496), .O(n547) );
  NAND_GATE U791 ( .I1(n549), .I2(n550), .O(n5010) );
  NAND_GATE U792 ( .I1(n495), .I2(donnee[27]), .O(n550) );
  NAND_GATE U793 ( .I1(\registres[24][27] ), .I2(n496), .O(n549) );
  NAND_GATE U794 ( .I1(n551), .I2(n552), .O(n5011) );
  NAND_GATE U795 ( .I1(n495), .I2(donnee[28]), .O(n552) );
  NAND_GATE U796 ( .I1(\registres[24][28] ), .I2(n496), .O(n551) );
  NAND_GATE U797 ( .I1(n553), .I2(n554), .O(n5012) );
  NAND_GATE U798 ( .I1(n495), .I2(donnee[29]), .O(n554) );
  NAND_GATE U799 ( .I1(\registres[24][29] ), .I2(n496), .O(n553) );
  NAND_GATE U800 ( .I1(n555), .I2(n556), .O(n5013) );
  NAND_GATE U801 ( .I1(n495), .I2(donnee[30]), .O(n556) );
  NAND_GATE U802 ( .I1(\registres[24][30] ), .I2(n496), .O(n555) );
  NAND_GATE U803 ( .I1(n557), .I2(n558), .O(n5014) );
  NAND_GATE U804 ( .I1(n495), .I2(donnee[31]), .O(n558) );
  AND_GATE U805 ( .I1(n559), .I2(n1), .O(n495) );
  NAND_GATE U806 ( .I1(\registres[24][31] ), .I2(n496), .O(n557) );
  NOR_GATE U807 ( .I1(n559), .I2(reset), .O(n496) );
  AND3_GATE U808 ( .I1(n83), .I2(cmd_ecr), .I3(n560), .O(n559) );
  AND_GATE U809 ( .I1(reg_dest[4]), .I2(reg_dest[3]), .O(n83) );
  NAND_GATE U810 ( .I1(n561), .I2(n562), .O(n5015) );
  NAND_GATE U811 ( .I1(n563), .I2(donnee[0]), .O(n562) );
  NAND_GATE U812 ( .I1(\registres[23][0] ), .I2(n564), .O(n561) );
  NAND_GATE U813 ( .I1(n565), .I2(n566), .O(n5016) );
  NAND_GATE U814 ( .I1(n563), .I2(donnee[1]), .O(n566) );
  NAND_GATE U815 ( .I1(\registres[23][1] ), .I2(n564), .O(n565) );
  NAND_GATE U816 ( .I1(n567), .I2(n568), .O(n5017) );
  NAND_GATE U817 ( .I1(n563), .I2(donnee[2]), .O(n568) );
  NAND_GATE U818 ( .I1(\registres[23][2] ), .I2(n564), .O(n567) );
  NAND_GATE U819 ( .I1(n569), .I2(n570), .O(n5018) );
  NAND_GATE U820 ( .I1(n563), .I2(donnee[3]), .O(n570) );
  NAND_GATE U821 ( .I1(\registres[23][3] ), .I2(n564), .O(n569) );
  NAND_GATE U822 ( .I1(n571), .I2(n572), .O(n5019) );
  NAND_GATE U823 ( .I1(n563), .I2(donnee[4]), .O(n572) );
  NAND_GATE U824 ( .I1(\registres[23][4] ), .I2(n564), .O(n571) );
  NAND_GATE U825 ( .I1(n573), .I2(n574), .O(n5020) );
  NAND_GATE U826 ( .I1(n563), .I2(donnee[5]), .O(n574) );
  NAND_GATE U827 ( .I1(\registres[23][5] ), .I2(n564), .O(n573) );
  NAND_GATE U828 ( .I1(n575), .I2(n576), .O(n5021) );
  NAND_GATE U829 ( .I1(n563), .I2(donnee[6]), .O(n576) );
  NAND_GATE U830 ( .I1(\registres[23][6] ), .I2(n564), .O(n575) );
  NAND_GATE U831 ( .I1(n577), .I2(n578), .O(n5022) );
  NAND_GATE U832 ( .I1(n563), .I2(donnee[7]), .O(n578) );
  NAND_GATE U833 ( .I1(\registres[23][7] ), .I2(n564), .O(n577) );
  NAND_GATE U834 ( .I1(n579), .I2(n580), .O(n5023) );
  NAND_GATE U835 ( .I1(n563), .I2(donnee[8]), .O(n580) );
  NAND_GATE U836 ( .I1(\registres[23][8] ), .I2(n564), .O(n579) );
  NAND_GATE U837 ( .I1(n581), .I2(n582), .O(n5024) );
  NAND_GATE U838 ( .I1(n563), .I2(donnee[9]), .O(n582) );
  NAND_GATE U839 ( .I1(\registres[23][9] ), .I2(n564), .O(n581) );
  NAND_GATE U840 ( .I1(n583), .I2(n584), .O(n5025) );
  NAND_GATE U841 ( .I1(n563), .I2(donnee[10]), .O(n584) );
  NAND_GATE U842 ( .I1(\registres[23][10] ), .I2(n564), .O(n583) );
  NAND_GATE U843 ( .I1(n585), .I2(n586), .O(n5026) );
  NAND_GATE U844 ( .I1(n563), .I2(donnee[11]), .O(n586) );
  NAND_GATE U845 ( .I1(\registres[23][11] ), .I2(n564), .O(n585) );
  NAND_GATE U846 ( .I1(n587), .I2(n588), .O(n5027) );
  NAND_GATE U847 ( .I1(n563), .I2(donnee[12]), .O(n588) );
  NAND_GATE U848 ( .I1(\registres[23][12] ), .I2(n564), .O(n587) );
  NAND_GATE U849 ( .I1(n589), .I2(n590), .O(n5028) );
  NAND_GATE U850 ( .I1(n563), .I2(donnee[13]), .O(n590) );
  NAND_GATE U851 ( .I1(\registres[23][13] ), .I2(n564), .O(n589) );
  NAND_GATE U852 ( .I1(n591), .I2(n592), .O(n5029) );
  NAND_GATE U853 ( .I1(n563), .I2(donnee[14]), .O(n592) );
  NAND_GATE U854 ( .I1(\registres[23][14] ), .I2(n564), .O(n591) );
  NAND_GATE U855 ( .I1(n593), .I2(n594), .O(n5030) );
  NAND_GATE U856 ( .I1(n563), .I2(donnee[15]), .O(n594) );
  NAND_GATE U857 ( .I1(\registres[23][15] ), .I2(n564), .O(n593) );
  NAND_GATE U858 ( .I1(n595), .I2(n596), .O(n5031) );
  NAND_GATE U859 ( .I1(n563), .I2(donnee[16]), .O(n596) );
  NAND_GATE U860 ( .I1(\registres[23][16] ), .I2(n564), .O(n595) );
  NAND_GATE U861 ( .I1(n597), .I2(n598), .O(n5032) );
  NAND_GATE U862 ( .I1(n563), .I2(donnee[17]), .O(n598) );
  NAND_GATE U863 ( .I1(\registres[23][17] ), .I2(n564), .O(n597) );
  NAND_GATE U864 ( .I1(n599), .I2(n600), .O(n5033) );
  NAND_GATE U865 ( .I1(n563), .I2(donnee[18]), .O(n600) );
  NAND_GATE U866 ( .I1(\registres[23][18] ), .I2(n564), .O(n599) );
  NAND_GATE U867 ( .I1(n601), .I2(n602), .O(n5034) );
  NAND_GATE U868 ( .I1(n563), .I2(donnee[19]), .O(n602) );
  NAND_GATE U869 ( .I1(\registres[23][19] ), .I2(n564), .O(n601) );
  NAND_GATE U870 ( .I1(n603), .I2(n604), .O(n5035) );
  NAND_GATE U871 ( .I1(n563), .I2(donnee[20]), .O(n604) );
  NAND_GATE U872 ( .I1(\registres[23][20] ), .I2(n564), .O(n603) );
  NAND_GATE U873 ( .I1(n605), .I2(n606), .O(n5036) );
  NAND_GATE U874 ( .I1(n563), .I2(donnee[21]), .O(n606) );
  NAND_GATE U875 ( .I1(\registres[23][21] ), .I2(n564), .O(n605) );
  NAND_GATE U876 ( .I1(n607), .I2(n608), .O(n5037) );
  NAND_GATE U877 ( .I1(n563), .I2(donnee[22]), .O(n608) );
  NAND_GATE U878 ( .I1(\registres[23][22] ), .I2(n564), .O(n607) );
  NAND_GATE U879 ( .I1(n609), .I2(n610), .O(n5038) );
  NAND_GATE U880 ( .I1(n563), .I2(donnee[23]), .O(n610) );
  NAND_GATE U881 ( .I1(\registres[23][23] ), .I2(n564), .O(n609) );
  NAND_GATE U882 ( .I1(n611), .I2(n612), .O(n5039) );
  NAND_GATE U883 ( .I1(n563), .I2(donnee[24]), .O(n612) );
  NAND_GATE U884 ( .I1(\registres[23][24] ), .I2(n564), .O(n611) );
  NAND_GATE U885 ( .I1(n613), .I2(n614), .O(n5040) );
  NAND_GATE U886 ( .I1(n563), .I2(donnee[25]), .O(n614) );
  NAND_GATE U887 ( .I1(\registres[23][25] ), .I2(n564), .O(n613) );
  NAND_GATE U888 ( .I1(n615), .I2(n616), .O(n5041) );
  NAND_GATE U889 ( .I1(n563), .I2(donnee[26]), .O(n616) );
  NAND_GATE U890 ( .I1(\registres[23][26] ), .I2(n564), .O(n615) );
  NAND_GATE U891 ( .I1(n617), .I2(n618), .O(n5042) );
  NAND_GATE U892 ( .I1(n563), .I2(donnee[27]), .O(n618) );
  NAND_GATE U893 ( .I1(\registres[23][27] ), .I2(n564), .O(n617) );
  NAND_GATE U894 ( .I1(n619), .I2(n620), .O(n5043) );
  NAND_GATE U895 ( .I1(n563), .I2(donnee[28]), .O(n620) );
  NAND_GATE U896 ( .I1(\registres[23][28] ), .I2(n564), .O(n619) );
  NAND_GATE U897 ( .I1(n621), .I2(n622), .O(n5044) );
  NAND_GATE U898 ( .I1(n563), .I2(donnee[29]), .O(n622) );
  NAND_GATE U899 ( .I1(\registres[23][29] ), .I2(n564), .O(n621) );
  NAND_GATE U900 ( .I1(n623), .I2(n624), .O(n5045) );
  NAND_GATE U901 ( .I1(n563), .I2(donnee[30]), .O(n624) );
  NAND_GATE U902 ( .I1(\registres[23][30] ), .I2(n564), .O(n623) );
  NAND_GATE U903 ( .I1(n625), .I2(n626), .O(n5046) );
  NAND_GATE U904 ( .I1(n563), .I2(donnee[31]), .O(n626) );
  AND_GATE U905 ( .I1(n627), .I2(n1), .O(n563) );
  NAND_GATE U906 ( .I1(\registres[23][31] ), .I2(n564), .O(n625) );
  NOR_GATE U907 ( .I1(n627), .I2(reset), .O(n564) );
  AND3_GATE U908 ( .I1(n84), .I2(cmd_ecr), .I3(n628), .O(n627) );
  NAND_GATE U909 ( .I1(n629), .I2(n630), .O(n5047) );
  NAND_GATE U910 ( .I1(n631), .I2(donnee[0]), .O(n630) );
  NAND_GATE U911 ( .I1(\registres[22][0] ), .I2(n632), .O(n629) );
  NAND_GATE U912 ( .I1(n633), .I2(n634), .O(n5048) );
  NAND_GATE U913 ( .I1(n631), .I2(donnee[1]), .O(n634) );
  NAND_GATE U914 ( .I1(\registres[22][1] ), .I2(n632), .O(n633) );
  NAND_GATE U915 ( .I1(n635), .I2(n636), .O(n5049) );
  NAND_GATE U916 ( .I1(n631), .I2(donnee[2]), .O(n636) );
  NAND_GATE U917 ( .I1(\registres[22][2] ), .I2(n632), .O(n635) );
  NAND_GATE U918 ( .I1(n637), .I2(n638), .O(n5050) );
  NAND_GATE U919 ( .I1(n631), .I2(donnee[3]), .O(n638) );
  NAND_GATE U920 ( .I1(\registres[22][3] ), .I2(n632), .O(n637) );
  NAND_GATE U921 ( .I1(n639), .I2(n640), .O(n5051) );
  NAND_GATE U922 ( .I1(n631), .I2(donnee[4]), .O(n640) );
  NAND_GATE U923 ( .I1(\registres[22][4] ), .I2(n632), .O(n639) );
  NAND_GATE U924 ( .I1(n641), .I2(n642), .O(n5052) );
  NAND_GATE U925 ( .I1(n631), .I2(donnee[5]), .O(n642) );
  NAND_GATE U926 ( .I1(\registres[22][5] ), .I2(n632), .O(n641) );
  NAND_GATE U927 ( .I1(n643), .I2(n644), .O(n5053) );
  NAND_GATE U928 ( .I1(n631), .I2(donnee[6]), .O(n644) );
  NAND_GATE U929 ( .I1(\registres[22][6] ), .I2(n632), .O(n643) );
  NAND_GATE U930 ( .I1(n645), .I2(n646), .O(n5054) );
  NAND_GATE U931 ( .I1(n631), .I2(donnee[7]), .O(n646) );
  NAND_GATE U932 ( .I1(\registres[22][7] ), .I2(n632), .O(n645) );
  NAND_GATE U933 ( .I1(n647), .I2(n648), .O(n5055) );
  NAND_GATE U934 ( .I1(n631), .I2(donnee[8]), .O(n648) );
  NAND_GATE U935 ( .I1(\registres[22][8] ), .I2(n632), .O(n647) );
  NAND_GATE U936 ( .I1(n649), .I2(n650), .O(n5056) );
  NAND_GATE U937 ( .I1(n631), .I2(donnee[9]), .O(n650) );
  NAND_GATE U938 ( .I1(\registres[22][9] ), .I2(n632), .O(n649) );
  NAND_GATE U939 ( .I1(n651), .I2(n652), .O(n5057) );
  NAND_GATE U940 ( .I1(n631), .I2(donnee[10]), .O(n652) );
  NAND_GATE U941 ( .I1(\registres[22][10] ), .I2(n632), .O(n651) );
  NAND_GATE U942 ( .I1(n653), .I2(n654), .O(n5058) );
  NAND_GATE U943 ( .I1(n631), .I2(donnee[11]), .O(n654) );
  NAND_GATE U944 ( .I1(\registres[22][11] ), .I2(n632), .O(n653) );
  NAND_GATE U945 ( .I1(n655), .I2(n656), .O(n5059) );
  NAND_GATE U946 ( .I1(n631), .I2(donnee[12]), .O(n656) );
  NAND_GATE U947 ( .I1(\registres[22][12] ), .I2(n632), .O(n655) );
  NAND_GATE U948 ( .I1(n657), .I2(n658), .O(n5060) );
  NAND_GATE U949 ( .I1(n631), .I2(donnee[13]), .O(n658) );
  NAND_GATE U950 ( .I1(\registres[22][13] ), .I2(n632), .O(n657) );
  NAND_GATE U951 ( .I1(n659), .I2(n660), .O(n5061) );
  NAND_GATE U952 ( .I1(n631), .I2(donnee[14]), .O(n660) );
  NAND_GATE U953 ( .I1(\registres[22][14] ), .I2(n632), .O(n659) );
  NAND_GATE U954 ( .I1(n661), .I2(n662), .O(n5062) );
  NAND_GATE U955 ( .I1(n631), .I2(donnee[15]), .O(n662) );
  NAND_GATE U956 ( .I1(\registres[22][15] ), .I2(n632), .O(n661) );
  NAND_GATE U957 ( .I1(n663), .I2(n664), .O(n5063) );
  NAND_GATE U958 ( .I1(n631), .I2(donnee[16]), .O(n664) );
  NAND_GATE U959 ( .I1(\registres[22][16] ), .I2(n632), .O(n663) );
  NAND_GATE U960 ( .I1(n665), .I2(n666), .O(n5064) );
  NAND_GATE U961 ( .I1(n631), .I2(donnee[17]), .O(n666) );
  NAND_GATE U962 ( .I1(\registres[22][17] ), .I2(n632), .O(n665) );
  NAND_GATE U963 ( .I1(n667), .I2(n668), .O(n5065) );
  NAND_GATE U964 ( .I1(n631), .I2(donnee[18]), .O(n668) );
  NAND_GATE U965 ( .I1(\registres[22][18] ), .I2(n632), .O(n667) );
  NAND_GATE U966 ( .I1(n669), .I2(n670), .O(n5066) );
  NAND_GATE U967 ( .I1(n631), .I2(donnee[19]), .O(n670) );
  NAND_GATE U968 ( .I1(\registres[22][19] ), .I2(n632), .O(n669) );
  NAND_GATE U969 ( .I1(n671), .I2(n672), .O(n5067) );
  NAND_GATE U970 ( .I1(n631), .I2(donnee[20]), .O(n672) );
  NAND_GATE U971 ( .I1(\registres[22][20] ), .I2(n632), .O(n671) );
  NAND_GATE U972 ( .I1(n673), .I2(n674), .O(n5068) );
  NAND_GATE U973 ( .I1(n631), .I2(donnee[21]), .O(n674) );
  NAND_GATE U974 ( .I1(\registres[22][21] ), .I2(n632), .O(n673) );
  NAND_GATE U975 ( .I1(n675), .I2(n676), .O(n5069) );
  NAND_GATE U976 ( .I1(n631), .I2(donnee[22]), .O(n676) );
  NAND_GATE U977 ( .I1(\registres[22][22] ), .I2(n632), .O(n675) );
  NAND_GATE U978 ( .I1(n677), .I2(n678), .O(n5070) );
  NAND_GATE U979 ( .I1(n631), .I2(donnee[23]), .O(n678) );
  NAND_GATE U980 ( .I1(\registres[22][23] ), .I2(n632), .O(n677) );
  NAND_GATE U981 ( .I1(n679), .I2(n680), .O(n5071) );
  NAND_GATE U982 ( .I1(n631), .I2(donnee[24]), .O(n680) );
  NAND_GATE U983 ( .I1(\registres[22][24] ), .I2(n632), .O(n679) );
  NAND_GATE U984 ( .I1(n681), .I2(n682), .O(n5072) );
  NAND_GATE U985 ( .I1(n631), .I2(donnee[25]), .O(n682) );
  NAND_GATE U986 ( .I1(\registres[22][25] ), .I2(n632), .O(n681) );
  NAND_GATE U987 ( .I1(n683), .I2(n684), .O(n5073) );
  NAND_GATE U988 ( .I1(n631), .I2(donnee[26]), .O(n684) );
  NAND_GATE U989 ( .I1(\registres[22][26] ), .I2(n632), .O(n683) );
  NAND_GATE U990 ( .I1(n685), .I2(n686), .O(n5074) );
  NAND_GATE U991 ( .I1(n631), .I2(donnee[27]), .O(n686) );
  NAND_GATE U992 ( .I1(\registres[22][27] ), .I2(n632), .O(n685) );
  NAND_GATE U993 ( .I1(n687), .I2(n688), .O(n5075) );
  NAND_GATE U994 ( .I1(n631), .I2(donnee[28]), .O(n688) );
  NAND_GATE U995 ( .I1(\registres[22][28] ), .I2(n632), .O(n687) );
  NAND_GATE U996 ( .I1(n689), .I2(n690), .O(n5076) );
  NAND_GATE U997 ( .I1(n631), .I2(donnee[29]), .O(n690) );
  NAND_GATE U998 ( .I1(\registres[22][29] ), .I2(n632), .O(n689) );
  NAND_GATE U999 ( .I1(n691), .I2(n692), .O(n5077) );
  NAND_GATE U1000 ( .I1(n631), .I2(donnee[30]), .O(n692) );
  NAND_GATE U1001 ( .I1(\registres[22][30] ), .I2(n632), .O(n691) );
  NAND_GATE U1002 ( .I1(n693), .I2(n694), .O(n5078) );
  NAND_GATE U1003 ( .I1(n631), .I2(donnee[31]), .O(n694) );
  AND_GATE U1004 ( .I1(n695), .I2(n1), .O(n631) );
  NAND_GATE U1005 ( .I1(\registres[22][31] ), .I2(n632), .O(n693) );
  NOR_GATE U1006 ( .I1(n695), .I2(reset), .O(n632) );
  AND3_GATE U1007 ( .I1(n152), .I2(cmd_ecr), .I3(n628), .O(n695) );
  NAND_GATE U1008 ( .I1(n696), .I2(n697), .O(n5079) );
  NAND_GATE U1009 ( .I1(n698), .I2(donnee[0]), .O(n697) );
  NAND_GATE U1010 ( .I1(\registres[21][0] ), .I2(n699), .O(n696) );
  NAND_GATE U1011 ( .I1(n700), .I2(n701), .O(n5080) );
  NAND_GATE U1012 ( .I1(n698), .I2(donnee[1]), .O(n701) );
  NAND_GATE U1013 ( .I1(\registres[21][1] ), .I2(n699), .O(n700) );
  NAND_GATE U1014 ( .I1(n702), .I2(n703), .O(n5081) );
  NAND_GATE U1015 ( .I1(n698), .I2(donnee[2]), .O(n703) );
  NAND_GATE U1016 ( .I1(\registres[21][2] ), .I2(n699), .O(n702) );
  NAND_GATE U1017 ( .I1(n704), .I2(n705), .O(n5082) );
  NAND_GATE U1018 ( .I1(n698), .I2(donnee[3]), .O(n705) );
  NAND_GATE U1019 ( .I1(\registres[21][3] ), .I2(n699), .O(n704) );
  NAND_GATE U1020 ( .I1(n706), .I2(n707), .O(n5083) );
  NAND_GATE U1021 ( .I1(n698), .I2(donnee[4]), .O(n707) );
  NAND_GATE U1022 ( .I1(\registres[21][4] ), .I2(n699), .O(n706) );
  NAND_GATE U1023 ( .I1(n708), .I2(n709), .O(n5084) );
  NAND_GATE U1024 ( .I1(n698), .I2(donnee[5]), .O(n709) );
  NAND_GATE U1025 ( .I1(\registres[21][5] ), .I2(n699), .O(n708) );
  NAND_GATE U1026 ( .I1(n710), .I2(n711), .O(n5085) );
  NAND_GATE U1027 ( .I1(n698), .I2(donnee[6]), .O(n711) );
  NAND_GATE U1028 ( .I1(\registres[21][6] ), .I2(n699), .O(n710) );
  NAND_GATE U1029 ( .I1(n712), .I2(n713), .O(n5086) );
  NAND_GATE U1030 ( .I1(n698), .I2(donnee[7]), .O(n713) );
  NAND_GATE U1031 ( .I1(\registres[21][7] ), .I2(n699), .O(n712) );
  NAND_GATE U1032 ( .I1(n714), .I2(n715), .O(n5087) );
  NAND_GATE U1033 ( .I1(n698), .I2(donnee[8]), .O(n715) );
  NAND_GATE U1034 ( .I1(\registres[21][8] ), .I2(n699), .O(n714) );
  NAND_GATE U1035 ( .I1(n716), .I2(n717), .O(n5088) );
  NAND_GATE U1036 ( .I1(n698), .I2(donnee[9]), .O(n717) );
  NAND_GATE U1037 ( .I1(\registres[21][9] ), .I2(n699), .O(n716) );
  NAND_GATE U1038 ( .I1(n718), .I2(n719), .O(n5089) );
  NAND_GATE U1039 ( .I1(n698), .I2(donnee[10]), .O(n719) );
  NAND_GATE U1040 ( .I1(\registres[21][10] ), .I2(n699), .O(n718) );
  NAND_GATE U1041 ( .I1(n720), .I2(n721), .O(n5090) );
  NAND_GATE U1042 ( .I1(n698), .I2(donnee[11]), .O(n721) );
  NAND_GATE U1043 ( .I1(\registres[21][11] ), .I2(n699), .O(n720) );
  NAND_GATE U1044 ( .I1(n722), .I2(n723), .O(n5091) );
  NAND_GATE U1045 ( .I1(n698), .I2(donnee[12]), .O(n723) );
  NAND_GATE U1046 ( .I1(\registres[21][12] ), .I2(n699), .O(n722) );
  NAND_GATE U1047 ( .I1(n724), .I2(n725), .O(n5092) );
  NAND_GATE U1048 ( .I1(n698), .I2(donnee[13]), .O(n725) );
  NAND_GATE U1049 ( .I1(\registres[21][13] ), .I2(n699), .O(n724) );
  NAND_GATE U1050 ( .I1(n726), .I2(n727), .O(n5093) );
  NAND_GATE U1051 ( .I1(n698), .I2(donnee[14]), .O(n727) );
  NAND_GATE U1052 ( .I1(\registres[21][14] ), .I2(n699), .O(n726) );
  NAND_GATE U1053 ( .I1(n728), .I2(n729), .O(n5094) );
  NAND_GATE U1054 ( .I1(n698), .I2(donnee[15]), .O(n729) );
  NAND_GATE U1055 ( .I1(\registres[21][15] ), .I2(n699), .O(n728) );
  NAND_GATE U1056 ( .I1(n730), .I2(n731), .O(n5095) );
  NAND_GATE U1057 ( .I1(n698), .I2(donnee[16]), .O(n731) );
  NAND_GATE U1058 ( .I1(\registres[21][16] ), .I2(n699), .O(n730) );
  NAND_GATE U1059 ( .I1(n732), .I2(n733), .O(n5096) );
  NAND_GATE U1060 ( .I1(n698), .I2(donnee[17]), .O(n733) );
  NAND_GATE U1061 ( .I1(\registres[21][17] ), .I2(n699), .O(n732) );
  NAND_GATE U1062 ( .I1(n734), .I2(n735), .O(n5097) );
  NAND_GATE U1063 ( .I1(n698), .I2(donnee[18]), .O(n735) );
  NAND_GATE U1064 ( .I1(\registres[21][18] ), .I2(n699), .O(n734) );
  NAND_GATE U1065 ( .I1(n736), .I2(n737), .O(n5098) );
  NAND_GATE U1066 ( .I1(n698), .I2(donnee[19]), .O(n737) );
  NAND_GATE U1067 ( .I1(\registres[21][19] ), .I2(n699), .O(n736) );
  NAND_GATE U1068 ( .I1(n738), .I2(n739), .O(n5099) );
  NAND_GATE U1069 ( .I1(n698), .I2(donnee[20]), .O(n739) );
  NAND_GATE U1070 ( .I1(\registres[21][20] ), .I2(n699), .O(n738) );
  NAND_GATE U1071 ( .I1(n740), .I2(n741), .O(n5100) );
  NAND_GATE U1072 ( .I1(n698), .I2(donnee[21]), .O(n741) );
  NAND_GATE U1073 ( .I1(\registres[21][21] ), .I2(n699), .O(n740) );
  NAND_GATE U1074 ( .I1(n742), .I2(n743), .O(n5101) );
  NAND_GATE U1075 ( .I1(n698), .I2(donnee[22]), .O(n743) );
  NAND_GATE U1076 ( .I1(\registres[21][22] ), .I2(n699), .O(n742) );
  NAND_GATE U1077 ( .I1(n744), .I2(n745), .O(n5102) );
  NAND_GATE U1078 ( .I1(n698), .I2(donnee[23]), .O(n745) );
  NAND_GATE U1079 ( .I1(\registres[21][23] ), .I2(n699), .O(n744) );
  NAND_GATE U1080 ( .I1(n746), .I2(n747), .O(n5103) );
  NAND_GATE U1081 ( .I1(n698), .I2(donnee[24]), .O(n747) );
  NAND_GATE U1082 ( .I1(\registres[21][24] ), .I2(n699), .O(n746) );
  NAND_GATE U1083 ( .I1(n748), .I2(n749), .O(n5104) );
  NAND_GATE U1084 ( .I1(n698), .I2(donnee[25]), .O(n749) );
  NAND_GATE U1085 ( .I1(\registres[21][25] ), .I2(n699), .O(n748) );
  NAND_GATE U1086 ( .I1(n750), .I2(n751), .O(n5105) );
  NAND_GATE U1087 ( .I1(n698), .I2(donnee[26]), .O(n751) );
  NAND_GATE U1088 ( .I1(\registres[21][26] ), .I2(n699), .O(n750) );
  NAND_GATE U1089 ( .I1(n752), .I2(n753), .O(n5106) );
  NAND_GATE U1090 ( .I1(n698), .I2(donnee[27]), .O(n753) );
  NAND_GATE U1091 ( .I1(\registres[21][27] ), .I2(n699), .O(n752) );
  NAND_GATE U1092 ( .I1(n754), .I2(n755), .O(n5107) );
  NAND_GATE U1093 ( .I1(n698), .I2(donnee[28]), .O(n755) );
  NAND_GATE U1094 ( .I1(\registres[21][28] ), .I2(n699), .O(n754) );
  NAND_GATE U1095 ( .I1(n756), .I2(n757), .O(n5108) );
  NAND_GATE U1096 ( .I1(n698), .I2(donnee[29]), .O(n757) );
  NAND_GATE U1097 ( .I1(\registres[21][29] ), .I2(n699), .O(n756) );
  NAND_GATE U1098 ( .I1(n758), .I2(n759), .O(n5109) );
  NAND_GATE U1099 ( .I1(n698), .I2(donnee[30]), .O(n759) );
  NAND_GATE U1100 ( .I1(\registres[21][30] ), .I2(n699), .O(n758) );
  NAND_GATE U1101 ( .I1(n760), .I2(n761), .O(n5110) );
  NAND_GATE U1102 ( .I1(n698), .I2(donnee[31]), .O(n761) );
  AND_GATE U1103 ( .I1(n762), .I2(n1), .O(n698) );
  NAND_GATE U1104 ( .I1(\registres[21][31] ), .I2(n699), .O(n760) );
  NOR_GATE U1105 ( .I1(n762), .I2(reset), .O(n699) );
  AND3_GATE U1106 ( .I1(n220), .I2(cmd_ecr), .I3(n628), .O(n762) );
  NAND_GATE U1107 ( .I1(n763), .I2(n764), .O(n5111) );
  NAND_GATE U1108 ( .I1(n765), .I2(donnee[0]), .O(n764) );
  NAND_GATE U1109 ( .I1(\registres[20][0] ), .I2(n766), .O(n763) );
  NAND_GATE U1110 ( .I1(n767), .I2(n768), .O(n5112) );
  NAND_GATE U1111 ( .I1(n765), .I2(donnee[1]), .O(n768) );
  NAND_GATE U1112 ( .I1(\registres[20][1] ), .I2(n766), .O(n767) );
  NAND_GATE U1113 ( .I1(n769), .I2(n770), .O(n5113) );
  NAND_GATE U1114 ( .I1(n765), .I2(donnee[2]), .O(n770) );
  NAND_GATE U1115 ( .I1(\registres[20][2] ), .I2(n766), .O(n769) );
  NAND_GATE U1116 ( .I1(n771), .I2(n772), .O(n5114) );
  NAND_GATE U1117 ( .I1(n765), .I2(donnee[3]), .O(n772) );
  NAND_GATE U1118 ( .I1(\registres[20][3] ), .I2(n766), .O(n771) );
  NAND_GATE U1119 ( .I1(n773), .I2(n774), .O(n5115) );
  NAND_GATE U1120 ( .I1(n765), .I2(donnee[4]), .O(n774) );
  NAND_GATE U1121 ( .I1(\registres[20][4] ), .I2(n766), .O(n773) );
  NAND_GATE U1122 ( .I1(n775), .I2(n776), .O(n5116) );
  NAND_GATE U1123 ( .I1(n765), .I2(donnee[5]), .O(n776) );
  NAND_GATE U1124 ( .I1(\registres[20][5] ), .I2(n766), .O(n775) );
  NAND_GATE U1125 ( .I1(n777), .I2(n778), .O(n5117) );
  NAND_GATE U1126 ( .I1(n765), .I2(donnee[6]), .O(n778) );
  NAND_GATE U1127 ( .I1(\registres[20][6] ), .I2(n766), .O(n777) );
  NAND_GATE U1128 ( .I1(n779), .I2(n780), .O(n5118) );
  NAND_GATE U1129 ( .I1(n765), .I2(donnee[7]), .O(n780) );
  NAND_GATE U1130 ( .I1(\registres[20][7] ), .I2(n766), .O(n779) );
  NAND_GATE U1131 ( .I1(n781), .I2(n782), .O(n5119) );
  NAND_GATE U1132 ( .I1(n765), .I2(donnee[8]), .O(n782) );
  NAND_GATE U1133 ( .I1(\registres[20][8] ), .I2(n766), .O(n781) );
  NAND_GATE U1134 ( .I1(n783), .I2(n784), .O(n5120) );
  NAND_GATE U1135 ( .I1(n765), .I2(donnee[9]), .O(n784) );
  NAND_GATE U1136 ( .I1(\registres[20][9] ), .I2(n766), .O(n783) );
  NAND_GATE U1137 ( .I1(n785), .I2(n786), .O(n5121) );
  NAND_GATE U1138 ( .I1(n765), .I2(donnee[10]), .O(n786) );
  NAND_GATE U1139 ( .I1(\registres[20][10] ), .I2(n766), .O(n785) );
  NAND_GATE U1140 ( .I1(n787), .I2(n788), .O(n5122) );
  NAND_GATE U1141 ( .I1(n765), .I2(donnee[11]), .O(n788) );
  NAND_GATE U1142 ( .I1(\registres[20][11] ), .I2(n766), .O(n787) );
  NAND_GATE U1143 ( .I1(n789), .I2(n790), .O(n5123) );
  NAND_GATE U1144 ( .I1(n765), .I2(donnee[12]), .O(n790) );
  NAND_GATE U1145 ( .I1(\registres[20][12] ), .I2(n766), .O(n789) );
  NAND_GATE U1146 ( .I1(n791), .I2(n792), .O(n5124) );
  NAND_GATE U1147 ( .I1(n765), .I2(donnee[13]), .O(n792) );
  NAND_GATE U1148 ( .I1(\registres[20][13] ), .I2(n766), .O(n791) );
  NAND_GATE U1149 ( .I1(n793), .I2(n794), .O(n5125) );
  NAND_GATE U1150 ( .I1(n765), .I2(donnee[14]), .O(n794) );
  NAND_GATE U1151 ( .I1(\registres[20][14] ), .I2(n766), .O(n793) );
  NAND_GATE U1152 ( .I1(n795), .I2(n796), .O(n5126) );
  NAND_GATE U1153 ( .I1(n765), .I2(donnee[15]), .O(n796) );
  NAND_GATE U1154 ( .I1(\registres[20][15] ), .I2(n766), .O(n795) );
  NAND_GATE U1155 ( .I1(n797), .I2(n798), .O(n5127) );
  NAND_GATE U1156 ( .I1(n765), .I2(donnee[16]), .O(n798) );
  NAND_GATE U1157 ( .I1(\registres[20][16] ), .I2(n766), .O(n797) );
  NAND_GATE U1158 ( .I1(n799), .I2(n800), .O(n5128) );
  NAND_GATE U1159 ( .I1(n765), .I2(donnee[17]), .O(n800) );
  NAND_GATE U1160 ( .I1(\registres[20][17] ), .I2(n766), .O(n799) );
  NAND_GATE U1161 ( .I1(n801), .I2(n802), .O(n5129) );
  NAND_GATE U1162 ( .I1(n765), .I2(donnee[18]), .O(n802) );
  NAND_GATE U1163 ( .I1(\registres[20][18] ), .I2(n766), .O(n801) );
  NAND_GATE U1164 ( .I1(n803), .I2(n804), .O(n5130) );
  NAND_GATE U1165 ( .I1(n765), .I2(donnee[19]), .O(n804) );
  NAND_GATE U1166 ( .I1(\registres[20][19] ), .I2(n766), .O(n803) );
  NAND_GATE U1167 ( .I1(n805), .I2(n806), .O(n5131) );
  NAND_GATE U1168 ( .I1(n765), .I2(donnee[20]), .O(n806) );
  NAND_GATE U1169 ( .I1(\registres[20][20] ), .I2(n766), .O(n805) );
  NAND_GATE U1170 ( .I1(n807), .I2(n808), .O(n5132) );
  NAND_GATE U1171 ( .I1(n765), .I2(donnee[21]), .O(n808) );
  NAND_GATE U1172 ( .I1(\registres[20][21] ), .I2(n766), .O(n807) );
  NAND_GATE U1173 ( .I1(n809), .I2(n810), .O(n5133) );
  NAND_GATE U1174 ( .I1(n765), .I2(donnee[22]), .O(n810) );
  NAND_GATE U1175 ( .I1(\registres[20][22] ), .I2(n766), .O(n809) );
  NAND_GATE U1176 ( .I1(n811), .I2(n812), .O(n5134) );
  NAND_GATE U1177 ( .I1(n765), .I2(donnee[23]), .O(n812) );
  NAND_GATE U1178 ( .I1(\registres[20][23] ), .I2(n766), .O(n811) );
  NAND_GATE U1179 ( .I1(n813), .I2(n814), .O(n5135) );
  NAND_GATE U1180 ( .I1(n765), .I2(donnee[24]), .O(n814) );
  NAND_GATE U1181 ( .I1(\registres[20][24] ), .I2(n766), .O(n813) );
  NAND_GATE U1182 ( .I1(n815), .I2(n816), .O(n5136) );
  NAND_GATE U1183 ( .I1(n765), .I2(donnee[25]), .O(n816) );
  NAND_GATE U1184 ( .I1(\registres[20][25] ), .I2(n766), .O(n815) );
  NAND_GATE U1185 ( .I1(n817), .I2(n818), .O(n5137) );
  NAND_GATE U1186 ( .I1(n765), .I2(donnee[26]), .O(n818) );
  NAND_GATE U1187 ( .I1(\registres[20][26] ), .I2(n766), .O(n817) );
  NAND_GATE U1188 ( .I1(n819), .I2(n820), .O(n5138) );
  NAND_GATE U1189 ( .I1(n765), .I2(donnee[27]), .O(n820) );
  NAND_GATE U1190 ( .I1(\registres[20][27] ), .I2(n766), .O(n819) );
  NAND_GATE U1191 ( .I1(n821), .I2(n822), .O(n5139) );
  NAND_GATE U1192 ( .I1(n765), .I2(donnee[28]), .O(n822) );
  NAND_GATE U1193 ( .I1(\registres[20][28] ), .I2(n766), .O(n821) );
  NAND_GATE U1194 ( .I1(n823), .I2(n824), .O(n5140) );
  NAND_GATE U1195 ( .I1(n765), .I2(donnee[29]), .O(n824) );
  NAND_GATE U1196 ( .I1(\registres[20][29] ), .I2(n766), .O(n823) );
  NAND_GATE U1197 ( .I1(n825), .I2(n826), .O(n5141) );
  NAND_GATE U1198 ( .I1(n765), .I2(donnee[30]), .O(n826) );
  NAND_GATE U1199 ( .I1(\registres[20][30] ), .I2(n766), .O(n825) );
  NAND_GATE U1200 ( .I1(n827), .I2(n828), .O(n5142) );
  NAND_GATE U1201 ( .I1(n765), .I2(donnee[31]), .O(n828) );
  AND_GATE U1202 ( .I1(n829), .I2(n1), .O(n765) );
  NAND_GATE U1203 ( .I1(\registres[20][31] ), .I2(n766), .O(n827) );
  NOR_GATE U1204 ( .I1(n829), .I2(reset), .O(n766) );
  AND3_GATE U1205 ( .I1(n288), .I2(cmd_ecr), .I3(n628), .O(n829) );
  NAND_GATE U1206 ( .I1(n830), .I2(n831), .O(n5143) );
  NAND_GATE U1207 ( .I1(n832), .I2(donnee[0]), .O(n831) );
  NAND_GATE U1208 ( .I1(\registres[19][0] ), .I2(n833), .O(n830) );
  NAND_GATE U1209 ( .I1(n834), .I2(n835), .O(n5144) );
  NAND_GATE U1210 ( .I1(n832), .I2(donnee[1]), .O(n835) );
  NAND_GATE U1211 ( .I1(\registres[19][1] ), .I2(n833), .O(n834) );
  NAND_GATE U1212 ( .I1(n836), .I2(n837), .O(n5145) );
  NAND_GATE U1213 ( .I1(n832), .I2(donnee[2]), .O(n837) );
  NAND_GATE U1214 ( .I1(\registres[19][2] ), .I2(n833), .O(n836) );
  NAND_GATE U1215 ( .I1(n838), .I2(n839), .O(n5146) );
  NAND_GATE U1216 ( .I1(n832), .I2(donnee[3]), .O(n839) );
  NAND_GATE U1217 ( .I1(\registres[19][3] ), .I2(n833), .O(n838) );
  NAND_GATE U1218 ( .I1(n840), .I2(n841), .O(n5147) );
  NAND_GATE U1219 ( .I1(n832), .I2(donnee[4]), .O(n841) );
  NAND_GATE U1220 ( .I1(\registres[19][4] ), .I2(n833), .O(n840) );
  NAND_GATE U1221 ( .I1(n842), .I2(n843), .O(n5148) );
  NAND_GATE U1222 ( .I1(n832), .I2(donnee[5]), .O(n843) );
  NAND_GATE U1223 ( .I1(\registres[19][5] ), .I2(n833), .O(n842) );
  NAND_GATE U1224 ( .I1(n844), .I2(n845), .O(n5149) );
  NAND_GATE U1225 ( .I1(n832), .I2(donnee[6]), .O(n845) );
  NAND_GATE U1226 ( .I1(\registres[19][6] ), .I2(n833), .O(n844) );
  NAND_GATE U1227 ( .I1(n846), .I2(n847), .O(n5150) );
  NAND_GATE U1228 ( .I1(n832), .I2(donnee[7]), .O(n847) );
  NAND_GATE U1229 ( .I1(\registres[19][7] ), .I2(n833), .O(n846) );
  NAND_GATE U1230 ( .I1(n848), .I2(n849), .O(n5151) );
  NAND_GATE U1231 ( .I1(n832), .I2(donnee[8]), .O(n849) );
  NAND_GATE U1232 ( .I1(\registres[19][8] ), .I2(n833), .O(n848) );
  NAND_GATE U1233 ( .I1(n850), .I2(n851), .O(n5152) );
  NAND_GATE U1234 ( .I1(n832), .I2(donnee[9]), .O(n851) );
  NAND_GATE U1235 ( .I1(\registres[19][9] ), .I2(n833), .O(n850) );
  NAND_GATE U1236 ( .I1(n852), .I2(n853), .O(n5153) );
  NAND_GATE U1237 ( .I1(n832), .I2(donnee[10]), .O(n853) );
  NAND_GATE U1238 ( .I1(\registres[19][10] ), .I2(n833), .O(n852) );
  NAND_GATE U1239 ( .I1(n854), .I2(n855), .O(n5154) );
  NAND_GATE U1240 ( .I1(n832), .I2(donnee[11]), .O(n855) );
  NAND_GATE U1241 ( .I1(\registres[19][11] ), .I2(n833), .O(n854) );
  NAND_GATE U1242 ( .I1(n856), .I2(n857), .O(n5155) );
  NAND_GATE U1243 ( .I1(n832), .I2(donnee[12]), .O(n857) );
  NAND_GATE U1244 ( .I1(\registres[19][12] ), .I2(n833), .O(n856) );
  NAND_GATE U1245 ( .I1(n858), .I2(n859), .O(n5156) );
  NAND_GATE U1246 ( .I1(n832), .I2(donnee[13]), .O(n859) );
  NAND_GATE U1247 ( .I1(\registres[19][13] ), .I2(n833), .O(n858) );
  NAND_GATE U1248 ( .I1(n860), .I2(n861), .O(n5157) );
  NAND_GATE U1249 ( .I1(n832), .I2(donnee[14]), .O(n861) );
  NAND_GATE U1250 ( .I1(\registres[19][14] ), .I2(n833), .O(n860) );
  NAND_GATE U1251 ( .I1(n862), .I2(n863), .O(n5158) );
  NAND_GATE U1252 ( .I1(n832), .I2(donnee[15]), .O(n863) );
  NAND_GATE U1253 ( .I1(\registres[19][15] ), .I2(n833), .O(n862) );
  NAND_GATE U1254 ( .I1(n864), .I2(n865), .O(n5159) );
  NAND_GATE U1255 ( .I1(n832), .I2(donnee[16]), .O(n865) );
  NAND_GATE U1256 ( .I1(\registres[19][16] ), .I2(n833), .O(n864) );
  NAND_GATE U1257 ( .I1(n866), .I2(n867), .O(n5160) );
  NAND_GATE U1258 ( .I1(n832), .I2(donnee[17]), .O(n867) );
  NAND_GATE U1259 ( .I1(\registres[19][17] ), .I2(n833), .O(n866) );
  NAND_GATE U1260 ( .I1(n868), .I2(n869), .O(n5161) );
  NAND_GATE U1261 ( .I1(n832), .I2(donnee[18]), .O(n869) );
  NAND_GATE U1262 ( .I1(\registres[19][18] ), .I2(n833), .O(n868) );
  NAND_GATE U1263 ( .I1(n870), .I2(n871), .O(n5162) );
  NAND_GATE U1264 ( .I1(n832), .I2(donnee[19]), .O(n871) );
  NAND_GATE U1265 ( .I1(\registres[19][19] ), .I2(n833), .O(n870) );
  NAND_GATE U1266 ( .I1(n872), .I2(n873), .O(n5163) );
  NAND_GATE U1267 ( .I1(n832), .I2(donnee[20]), .O(n873) );
  NAND_GATE U1268 ( .I1(\registres[19][20] ), .I2(n833), .O(n872) );
  NAND_GATE U1269 ( .I1(n874), .I2(n875), .O(n5164) );
  NAND_GATE U1270 ( .I1(n832), .I2(donnee[21]), .O(n875) );
  NAND_GATE U1271 ( .I1(\registres[19][21] ), .I2(n833), .O(n874) );
  NAND_GATE U1272 ( .I1(n876), .I2(n877), .O(n5165) );
  NAND_GATE U1273 ( .I1(n832), .I2(donnee[22]), .O(n877) );
  NAND_GATE U1274 ( .I1(\registres[19][22] ), .I2(n833), .O(n876) );
  NAND_GATE U1275 ( .I1(n878), .I2(n879), .O(n5166) );
  NAND_GATE U1276 ( .I1(n832), .I2(donnee[23]), .O(n879) );
  NAND_GATE U1277 ( .I1(\registres[19][23] ), .I2(n833), .O(n878) );
  NAND_GATE U1278 ( .I1(n880), .I2(n881), .O(n5167) );
  NAND_GATE U1279 ( .I1(n832), .I2(donnee[24]), .O(n881) );
  NAND_GATE U1280 ( .I1(\registres[19][24] ), .I2(n833), .O(n880) );
  NAND_GATE U1281 ( .I1(n882), .I2(n883), .O(n5168) );
  NAND_GATE U1282 ( .I1(n832), .I2(donnee[25]), .O(n883) );
  NAND_GATE U1283 ( .I1(\registres[19][25] ), .I2(n833), .O(n882) );
  NAND_GATE U1284 ( .I1(n884), .I2(n885), .O(n5169) );
  NAND_GATE U1285 ( .I1(n832), .I2(donnee[26]), .O(n885) );
  NAND_GATE U1286 ( .I1(\registres[19][26] ), .I2(n833), .O(n884) );
  NAND_GATE U1287 ( .I1(n886), .I2(n887), .O(n5170) );
  NAND_GATE U1288 ( .I1(n832), .I2(donnee[27]), .O(n887) );
  NAND_GATE U1289 ( .I1(\registres[19][27] ), .I2(n833), .O(n886) );
  NAND_GATE U1290 ( .I1(n888), .I2(n889), .O(n5171) );
  NAND_GATE U1291 ( .I1(n832), .I2(donnee[28]), .O(n889) );
  NAND_GATE U1292 ( .I1(\registres[19][28] ), .I2(n833), .O(n888) );
  NAND_GATE U1293 ( .I1(n890), .I2(n891), .O(n5172) );
  NAND_GATE U1294 ( .I1(n832), .I2(donnee[29]), .O(n891) );
  NAND_GATE U1295 ( .I1(\registres[19][29] ), .I2(n833), .O(n890) );
  NAND_GATE U1296 ( .I1(n892), .I2(n893), .O(n5173) );
  NAND_GATE U1297 ( .I1(n832), .I2(donnee[30]), .O(n893) );
  NAND_GATE U1298 ( .I1(\registres[19][30] ), .I2(n833), .O(n892) );
  NAND_GATE U1299 ( .I1(n894), .I2(n895), .O(n5174) );
  NAND_GATE U1300 ( .I1(n832), .I2(donnee[31]), .O(n895) );
  AND_GATE U1301 ( .I1(n896), .I2(n1), .O(n832) );
  NAND_GATE U1302 ( .I1(\registres[19][31] ), .I2(n833), .O(n894) );
  NOR_GATE U1303 ( .I1(n896), .I2(reset), .O(n833) );
  AND3_GATE U1304 ( .I1(n356), .I2(cmd_ecr), .I3(n628), .O(n896) );
  NAND_GATE U1305 ( .I1(n897), .I2(n898), .O(n5175) );
  NAND_GATE U1306 ( .I1(n899), .I2(donnee[0]), .O(n898) );
  NAND_GATE U1307 ( .I1(\registres[18][0] ), .I2(n900), .O(n897) );
  NAND_GATE U1308 ( .I1(n901), .I2(n902), .O(n5176) );
  NAND_GATE U1309 ( .I1(n899), .I2(donnee[1]), .O(n902) );
  NAND_GATE U1310 ( .I1(\registres[18][1] ), .I2(n900), .O(n901) );
  NAND_GATE U1311 ( .I1(n903), .I2(n904), .O(n5177) );
  NAND_GATE U1312 ( .I1(n899), .I2(donnee[2]), .O(n904) );
  NAND_GATE U1313 ( .I1(\registres[18][2] ), .I2(n900), .O(n903) );
  NAND_GATE U1314 ( .I1(n905), .I2(n906), .O(n5178) );
  NAND_GATE U1315 ( .I1(n899), .I2(donnee[3]), .O(n906) );
  NAND_GATE U1316 ( .I1(\registres[18][3] ), .I2(n900), .O(n905) );
  NAND_GATE U1317 ( .I1(n907), .I2(n908), .O(n5179) );
  NAND_GATE U1318 ( .I1(n899), .I2(donnee[4]), .O(n908) );
  NAND_GATE U1319 ( .I1(\registres[18][4] ), .I2(n900), .O(n907) );
  NAND_GATE U1320 ( .I1(n909), .I2(n910), .O(n5180) );
  NAND_GATE U1321 ( .I1(n899), .I2(donnee[5]), .O(n910) );
  NAND_GATE U1322 ( .I1(\registres[18][5] ), .I2(n900), .O(n909) );
  NAND_GATE U1323 ( .I1(n911), .I2(n912), .O(n5181) );
  NAND_GATE U1324 ( .I1(n899), .I2(donnee[6]), .O(n912) );
  NAND_GATE U1325 ( .I1(\registres[18][6] ), .I2(n900), .O(n911) );
  NAND_GATE U1326 ( .I1(n913), .I2(n914), .O(n5182) );
  NAND_GATE U1327 ( .I1(n899), .I2(donnee[7]), .O(n914) );
  NAND_GATE U1328 ( .I1(\registres[18][7] ), .I2(n900), .O(n913) );
  NAND_GATE U1329 ( .I1(n915), .I2(n916), .O(n5183) );
  NAND_GATE U1330 ( .I1(n899), .I2(donnee[8]), .O(n916) );
  NAND_GATE U1331 ( .I1(\registres[18][8] ), .I2(n900), .O(n915) );
  NAND_GATE U1332 ( .I1(n917), .I2(n918), .O(n5184) );
  NAND_GATE U1333 ( .I1(n899), .I2(donnee[9]), .O(n918) );
  NAND_GATE U1334 ( .I1(\registres[18][9] ), .I2(n900), .O(n917) );
  NAND_GATE U1335 ( .I1(n919), .I2(n920), .O(n5185) );
  NAND_GATE U1336 ( .I1(n899), .I2(donnee[10]), .O(n920) );
  NAND_GATE U1337 ( .I1(\registres[18][10] ), .I2(n900), .O(n919) );
  NAND_GATE U1338 ( .I1(n921), .I2(n922), .O(n5186) );
  NAND_GATE U1339 ( .I1(n899), .I2(donnee[11]), .O(n922) );
  NAND_GATE U1340 ( .I1(\registres[18][11] ), .I2(n900), .O(n921) );
  NAND_GATE U1341 ( .I1(n923), .I2(n924), .O(n5187) );
  NAND_GATE U1342 ( .I1(n899), .I2(donnee[12]), .O(n924) );
  NAND_GATE U1343 ( .I1(\registres[18][12] ), .I2(n900), .O(n923) );
  NAND_GATE U1344 ( .I1(n925), .I2(n926), .O(n5188) );
  NAND_GATE U1345 ( .I1(n899), .I2(donnee[13]), .O(n926) );
  NAND_GATE U1346 ( .I1(\registres[18][13] ), .I2(n900), .O(n925) );
  NAND_GATE U1347 ( .I1(n927), .I2(n928), .O(n5189) );
  NAND_GATE U1348 ( .I1(n899), .I2(donnee[14]), .O(n928) );
  NAND_GATE U1349 ( .I1(\registres[18][14] ), .I2(n900), .O(n927) );
  NAND_GATE U1350 ( .I1(n929), .I2(n930), .O(n5190) );
  NAND_GATE U1351 ( .I1(n899), .I2(donnee[15]), .O(n930) );
  NAND_GATE U1352 ( .I1(\registres[18][15] ), .I2(n900), .O(n929) );
  NAND_GATE U1353 ( .I1(n931), .I2(n932), .O(n5191) );
  NAND_GATE U1354 ( .I1(n899), .I2(donnee[16]), .O(n932) );
  NAND_GATE U1355 ( .I1(\registres[18][16] ), .I2(n900), .O(n931) );
  NAND_GATE U1356 ( .I1(n933), .I2(n934), .O(n5192) );
  NAND_GATE U1357 ( .I1(n899), .I2(donnee[17]), .O(n934) );
  NAND_GATE U1358 ( .I1(\registres[18][17] ), .I2(n900), .O(n933) );
  NAND_GATE U1359 ( .I1(n935), .I2(n936), .O(n5193) );
  NAND_GATE U1360 ( .I1(n899), .I2(donnee[18]), .O(n936) );
  NAND_GATE U1361 ( .I1(\registres[18][18] ), .I2(n900), .O(n935) );
  NAND_GATE U1362 ( .I1(n937), .I2(n938), .O(n5194) );
  NAND_GATE U1363 ( .I1(n899), .I2(donnee[19]), .O(n938) );
  NAND_GATE U1364 ( .I1(\registres[18][19] ), .I2(n900), .O(n937) );
  NAND_GATE U1365 ( .I1(n939), .I2(n940), .O(n5195) );
  NAND_GATE U1366 ( .I1(n899), .I2(donnee[20]), .O(n940) );
  NAND_GATE U1367 ( .I1(\registres[18][20] ), .I2(n900), .O(n939) );
  NAND_GATE U1368 ( .I1(n941), .I2(n942), .O(n5196) );
  NAND_GATE U1369 ( .I1(n899), .I2(donnee[21]), .O(n942) );
  NAND_GATE U1370 ( .I1(\registres[18][21] ), .I2(n900), .O(n941) );
  NAND_GATE U1371 ( .I1(n943), .I2(n944), .O(n5197) );
  NAND_GATE U1372 ( .I1(n899), .I2(donnee[22]), .O(n944) );
  NAND_GATE U1373 ( .I1(\registres[18][22] ), .I2(n900), .O(n943) );
  NAND_GATE U1374 ( .I1(n945), .I2(n946), .O(n5198) );
  NAND_GATE U1375 ( .I1(n899), .I2(donnee[23]), .O(n946) );
  NAND_GATE U1376 ( .I1(\registres[18][23] ), .I2(n900), .O(n945) );
  NAND_GATE U1377 ( .I1(n947), .I2(n948), .O(n5199) );
  NAND_GATE U1378 ( .I1(n899), .I2(donnee[24]), .O(n948) );
  NAND_GATE U1379 ( .I1(\registres[18][24] ), .I2(n900), .O(n947) );
  NAND_GATE U1380 ( .I1(n949), .I2(n950), .O(n5200) );
  NAND_GATE U1381 ( .I1(n899), .I2(donnee[25]), .O(n950) );
  NAND_GATE U1382 ( .I1(\registres[18][25] ), .I2(n900), .O(n949) );
  NAND_GATE U1383 ( .I1(n951), .I2(n952), .O(n5201) );
  NAND_GATE U1384 ( .I1(n899), .I2(donnee[26]), .O(n952) );
  NAND_GATE U1385 ( .I1(\registres[18][26] ), .I2(n900), .O(n951) );
  NAND_GATE U1386 ( .I1(n953), .I2(n954), .O(n5202) );
  NAND_GATE U1387 ( .I1(n899), .I2(donnee[27]), .O(n954) );
  NAND_GATE U1388 ( .I1(\registres[18][27] ), .I2(n900), .O(n953) );
  NAND_GATE U1389 ( .I1(n955), .I2(n956), .O(n5203) );
  NAND_GATE U1390 ( .I1(n899), .I2(donnee[28]), .O(n956) );
  NAND_GATE U1391 ( .I1(\registres[18][28] ), .I2(n900), .O(n955) );
  NAND_GATE U1392 ( .I1(n957), .I2(n958), .O(n5204) );
  NAND_GATE U1393 ( .I1(n899), .I2(donnee[29]), .O(n958) );
  NAND_GATE U1394 ( .I1(\registres[18][29] ), .I2(n900), .O(n957) );
  NAND_GATE U1395 ( .I1(n959), .I2(n960), .O(n5205) );
  NAND_GATE U1396 ( .I1(n899), .I2(donnee[30]), .O(n960) );
  NAND_GATE U1397 ( .I1(\registres[18][30] ), .I2(n900), .O(n959) );
  NAND_GATE U1398 ( .I1(n961), .I2(n962), .O(n5206) );
  NAND_GATE U1399 ( .I1(n899), .I2(donnee[31]), .O(n962) );
  AND_GATE U1400 ( .I1(n963), .I2(n1), .O(n899) );
  NAND_GATE U1401 ( .I1(\registres[18][31] ), .I2(n900), .O(n961) );
  NOR_GATE U1402 ( .I1(n963), .I2(reset), .O(n900) );
  AND3_GATE U1403 ( .I1(n424), .I2(cmd_ecr), .I3(n628), .O(n963) );
  NAND_GATE U1404 ( .I1(n964), .I2(n965), .O(n5207) );
  NAND_GATE U1405 ( .I1(n966), .I2(donnee[0]), .O(n965) );
  NAND_GATE U1406 ( .I1(\registres[17][0] ), .I2(n967), .O(n964) );
  NAND_GATE U1407 ( .I1(n968), .I2(n969), .O(n5208) );
  NAND_GATE U1408 ( .I1(n966), .I2(donnee[1]), .O(n969) );
  NAND_GATE U1409 ( .I1(\registres[17][1] ), .I2(n967), .O(n968) );
  NAND_GATE U1410 ( .I1(n970), .I2(n971), .O(n5209) );
  NAND_GATE U1411 ( .I1(n966), .I2(donnee[2]), .O(n971) );
  NAND_GATE U1412 ( .I1(\registres[17][2] ), .I2(n967), .O(n970) );
  NAND_GATE U1413 ( .I1(n972), .I2(n973), .O(n5210) );
  NAND_GATE U1414 ( .I1(n966), .I2(donnee[3]), .O(n973) );
  NAND_GATE U1415 ( .I1(\registres[17][3] ), .I2(n967), .O(n972) );
  NAND_GATE U1416 ( .I1(n974), .I2(n975), .O(n5211) );
  NAND_GATE U1417 ( .I1(n966), .I2(donnee[4]), .O(n975) );
  NAND_GATE U1418 ( .I1(\registres[17][4] ), .I2(n967), .O(n974) );
  NAND_GATE U1419 ( .I1(n976), .I2(n977), .O(n5212) );
  NAND_GATE U1420 ( .I1(n966), .I2(donnee[5]), .O(n977) );
  NAND_GATE U1421 ( .I1(\registres[17][5] ), .I2(n967), .O(n976) );
  NAND_GATE U1422 ( .I1(n978), .I2(n979), .O(n5213) );
  NAND_GATE U1423 ( .I1(n966), .I2(donnee[6]), .O(n979) );
  NAND_GATE U1424 ( .I1(\registres[17][6] ), .I2(n967), .O(n978) );
  NAND_GATE U1425 ( .I1(n980), .I2(n981), .O(n5214) );
  NAND_GATE U1426 ( .I1(n966), .I2(donnee[7]), .O(n981) );
  NAND_GATE U1427 ( .I1(\registres[17][7] ), .I2(n967), .O(n980) );
  NAND_GATE U1428 ( .I1(n982), .I2(n983), .O(n5215) );
  NAND_GATE U1429 ( .I1(n966), .I2(donnee[8]), .O(n983) );
  NAND_GATE U1430 ( .I1(\registres[17][8] ), .I2(n967), .O(n982) );
  NAND_GATE U1431 ( .I1(n984), .I2(n985), .O(n5216) );
  NAND_GATE U1432 ( .I1(n966), .I2(donnee[9]), .O(n985) );
  NAND_GATE U1433 ( .I1(\registres[17][9] ), .I2(n967), .O(n984) );
  NAND_GATE U1434 ( .I1(n986), .I2(n987), .O(n5217) );
  NAND_GATE U1435 ( .I1(n966), .I2(donnee[10]), .O(n987) );
  NAND_GATE U1436 ( .I1(\registres[17][10] ), .I2(n967), .O(n986) );
  NAND_GATE U1437 ( .I1(n988), .I2(n989), .O(n5218) );
  NAND_GATE U1438 ( .I1(n966), .I2(donnee[11]), .O(n989) );
  NAND_GATE U1439 ( .I1(\registres[17][11] ), .I2(n967), .O(n988) );
  NAND_GATE U1440 ( .I1(n990), .I2(n991), .O(n5219) );
  NAND_GATE U1441 ( .I1(n966), .I2(donnee[12]), .O(n991) );
  NAND_GATE U1442 ( .I1(\registres[17][12] ), .I2(n967), .O(n990) );
  NAND_GATE U1443 ( .I1(n992), .I2(n993), .O(n5220) );
  NAND_GATE U1444 ( .I1(n966), .I2(donnee[13]), .O(n993) );
  NAND_GATE U1445 ( .I1(\registres[17][13] ), .I2(n967), .O(n992) );
  NAND_GATE U1446 ( .I1(n994), .I2(n995), .O(n5221) );
  NAND_GATE U1447 ( .I1(n966), .I2(donnee[14]), .O(n995) );
  NAND_GATE U1448 ( .I1(\registres[17][14] ), .I2(n967), .O(n994) );
  NAND_GATE U1449 ( .I1(n996), .I2(n997), .O(n5222) );
  NAND_GATE U1450 ( .I1(n966), .I2(donnee[15]), .O(n997) );
  NAND_GATE U1451 ( .I1(\registres[17][15] ), .I2(n967), .O(n996) );
  NAND_GATE U1452 ( .I1(n998), .I2(n999), .O(n5223) );
  NAND_GATE U1453 ( .I1(n966), .I2(donnee[16]), .O(n999) );
  NAND_GATE U1454 ( .I1(\registres[17][16] ), .I2(n967), .O(n998) );
  NAND_GATE U1455 ( .I1(n1000), .I2(n1001), .O(n5224) );
  NAND_GATE U1456 ( .I1(n966), .I2(donnee[17]), .O(n1001) );
  NAND_GATE U1457 ( .I1(\registres[17][17] ), .I2(n967), .O(n1000) );
  NAND_GATE U1458 ( .I1(n1002), .I2(n1003), .O(n5225) );
  NAND_GATE U1459 ( .I1(n966), .I2(donnee[18]), .O(n1003) );
  NAND_GATE U1460 ( .I1(\registres[17][18] ), .I2(n967), .O(n1002) );
  NAND_GATE U1461 ( .I1(n1004), .I2(n1005), .O(n5226) );
  NAND_GATE U1462 ( .I1(n966), .I2(donnee[19]), .O(n1005) );
  NAND_GATE U1463 ( .I1(\registres[17][19] ), .I2(n967), .O(n1004) );
  NAND_GATE U1464 ( .I1(n1006), .I2(n1007), .O(n5227) );
  NAND_GATE U1465 ( .I1(n966), .I2(donnee[20]), .O(n1007) );
  NAND_GATE U1466 ( .I1(\registres[17][20] ), .I2(n967), .O(n1006) );
  NAND_GATE U1467 ( .I1(n1008), .I2(n1009), .O(n5228) );
  NAND_GATE U1468 ( .I1(n966), .I2(donnee[21]), .O(n1009) );
  NAND_GATE U1469 ( .I1(\registres[17][21] ), .I2(n967), .O(n1008) );
  NAND_GATE U1470 ( .I1(n1010), .I2(n1011), .O(n5229) );
  NAND_GATE U1471 ( .I1(n966), .I2(donnee[22]), .O(n1011) );
  NAND_GATE U1472 ( .I1(\registres[17][22] ), .I2(n967), .O(n1010) );
  NAND_GATE U1473 ( .I1(n1012), .I2(n1013), .O(n5230) );
  NAND_GATE U1474 ( .I1(n966), .I2(donnee[23]), .O(n1013) );
  NAND_GATE U1475 ( .I1(\registres[17][23] ), .I2(n967), .O(n1012) );
  NAND_GATE U1476 ( .I1(n1014), .I2(n1015), .O(n5231) );
  NAND_GATE U1477 ( .I1(n966), .I2(donnee[24]), .O(n1015) );
  NAND_GATE U1478 ( .I1(\registres[17][24] ), .I2(n967), .O(n1014) );
  NAND_GATE U1479 ( .I1(n1016), .I2(n1017), .O(n5232) );
  NAND_GATE U1480 ( .I1(n966), .I2(donnee[25]), .O(n1017) );
  NAND_GATE U1481 ( .I1(\registres[17][25] ), .I2(n967), .O(n1016) );
  NAND_GATE U1482 ( .I1(n1018), .I2(n1019), .O(n5233) );
  NAND_GATE U1483 ( .I1(n966), .I2(donnee[26]), .O(n1019) );
  NAND_GATE U1484 ( .I1(\registres[17][26] ), .I2(n967), .O(n1018) );
  NAND_GATE U1485 ( .I1(n1020), .I2(n1021), .O(n5234) );
  NAND_GATE U1486 ( .I1(n966), .I2(donnee[27]), .O(n1021) );
  NAND_GATE U1487 ( .I1(\registres[17][27] ), .I2(n967), .O(n1020) );
  NAND_GATE U1488 ( .I1(n1022), .I2(n1023), .O(n5235) );
  NAND_GATE U1489 ( .I1(n966), .I2(donnee[28]), .O(n1023) );
  NAND_GATE U1490 ( .I1(\registres[17][28] ), .I2(n967), .O(n1022) );
  NAND_GATE U1491 ( .I1(n1024), .I2(n1025), .O(n5236) );
  NAND_GATE U1492 ( .I1(n966), .I2(donnee[29]), .O(n1025) );
  NAND_GATE U1493 ( .I1(\registres[17][29] ), .I2(n967), .O(n1024) );
  NAND_GATE U1494 ( .I1(n1026), .I2(n1027), .O(n5237) );
  NAND_GATE U1495 ( .I1(n966), .I2(donnee[30]), .O(n1027) );
  NAND_GATE U1496 ( .I1(\registres[17][30] ), .I2(n967), .O(n1026) );
  NAND_GATE U1497 ( .I1(n1028), .I2(n1029), .O(n5238) );
  NAND_GATE U1498 ( .I1(n966), .I2(donnee[31]), .O(n1029) );
  AND_GATE U1499 ( .I1(n1030), .I2(n1), .O(n966) );
  NAND_GATE U1500 ( .I1(\registres[17][31] ), .I2(n967), .O(n1028) );
  NOR_GATE U1501 ( .I1(n1030), .I2(reset), .O(n967) );
  AND3_GATE U1502 ( .I1(n492), .I2(cmd_ecr), .I3(n628), .O(n1030) );
  NAND_GATE U1503 ( .I1(n1031), .I2(n1032), .O(n5239) );
  NAND_GATE U1504 ( .I1(n1033), .I2(donnee[0]), .O(n1032) );
  NAND_GATE U1505 ( .I1(\registres[16][0] ), .I2(n1034), .O(n1031) );
  NAND_GATE U1506 ( .I1(n1035), .I2(n1036), .O(n5240) );
  NAND_GATE U1507 ( .I1(n1033), .I2(donnee[1]), .O(n1036) );
  NAND_GATE U1508 ( .I1(\registres[16][1] ), .I2(n1034), .O(n1035) );
  NAND_GATE U1509 ( .I1(n1037), .I2(n1038), .O(n5241) );
  NAND_GATE U1510 ( .I1(n1033), .I2(donnee[2]), .O(n1038) );
  NAND_GATE U1511 ( .I1(\registres[16][2] ), .I2(n1034), .O(n1037) );
  NAND_GATE U1512 ( .I1(n1039), .I2(n1040), .O(n5242) );
  NAND_GATE U1513 ( .I1(n1033), .I2(donnee[3]), .O(n1040) );
  NAND_GATE U1514 ( .I1(\registres[16][3] ), .I2(n1034), .O(n1039) );
  NAND_GATE U1515 ( .I1(n1041), .I2(n1042), .O(n5243) );
  NAND_GATE U1516 ( .I1(n1033), .I2(donnee[4]), .O(n1042) );
  NAND_GATE U1517 ( .I1(\registres[16][4] ), .I2(n1034), .O(n1041) );
  NAND_GATE U1518 ( .I1(n1043), .I2(n1044), .O(n5244) );
  NAND_GATE U1519 ( .I1(n1033), .I2(donnee[5]), .O(n1044) );
  NAND_GATE U1520 ( .I1(\registres[16][5] ), .I2(n1034), .O(n1043) );
  NAND_GATE U1521 ( .I1(n1045), .I2(n1046), .O(n5245) );
  NAND_GATE U1522 ( .I1(n1033), .I2(donnee[6]), .O(n1046) );
  NAND_GATE U1523 ( .I1(\registres[16][6] ), .I2(n1034), .O(n1045) );
  NAND_GATE U1524 ( .I1(n1047), .I2(n1048), .O(n5246) );
  NAND_GATE U1525 ( .I1(n1033), .I2(donnee[7]), .O(n1048) );
  NAND_GATE U1526 ( .I1(\registres[16][7] ), .I2(n1034), .O(n1047) );
  NAND_GATE U1527 ( .I1(n1049), .I2(n1050), .O(n5247) );
  NAND_GATE U1528 ( .I1(n1033), .I2(donnee[8]), .O(n1050) );
  NAND_GATE U1529 ( .I1(\registres[16][8] ), .I2(n1034), .O(n1049) );
  NAND_GATE U1530 ( .I1(n1051), .I2(n1052), .O(n5248) );
  NAND_GATE U1531 ( .I1(n1033), .I2(donnee[9]), .O(n1052) );
  NAND_GATE U1532 ( .I1(\registres[16][9] ), .I2(n1034), .O(n1051) );
  NAND_GATE U1533 ( .I1(n1053), .I2(n1054), .O(n5249) );
  NAND_GATE U1534 ( .I1(n1033), .I2(donnee[10]), .O(n1054) );
  NAND_GATE U1535 ( .I1(\registres[16][10] ), .I2(n1034), .O(n1053) );
  NAND_GATE U1536 ( .I1(n1055), .I2(n1056), .O(n5250) );
  NAND_GATE U1537 ( .I1(n1033), .I2(donnee[11]), .O(n1056) );
  NAND_GATE U1538 ( .I1(\registres[16][11] ), .I2(n1034), .O(n1055) );
  NAND_GATE U1539 ( .I1(n1057), .I2(n1058), .O(n5251) );
  NAND_GATE U1540 ( .I1(n1033), .I2(donnee[12]), .O(n1058) );
  NAND_GATE U1541 ( .I1(\registres[16][12] ), .I2(n1034), .O(n1057) );
  NAND_GATE U1542 ( .I1(n1059), .I2(n1060), .O(n5252) );
  NAND_GATE U1543 ( .I1(n1033), .I2(donnee[13]), .O(n1060) );
  NAND_GATE U1544 ( .I1(\registres[16][13] ), .I2(n1034), .O(n1059) );
  NAND_GATE U1545 ( .I1(n1061), .I2(n1062), .O(n5253) );
  NAND_GATE U1546 ( .I1(n1033), .I2(donnee[14]), .O(n1062) );
  NAND_GATE U1547 ( .I1(\registres[16][14] ), .I2(n1034), .O(n1061) );
  NAND_GATE U1548 ( .I1(n1063), .I2(n1064), .O(n5254) );
  NAND_GATE U1549 ( .I1(n1033), .I2(donnee[15]), .O(n1064) );
  NAND_GATE U1550 ( .I1(\registres[16][15] ), .I2(n1034), .O(n1063) );
  NAND_GATE U1551 ( .I1(n1065), .I2(n1066), .O(n5255) );
  NAND_GATE U1552 ( .I1(n1033), .I2(donnee[16]), .O(n1066) );
  NAND_GATE U1553 ( .I1(\registres[16][16] ), .I2(n1034), .O(n1065) );
  NAND_GATE U1554 ( .I1(n1067), .I2(n1068), .O(n5256) );
  NAND_GATE U1555 ( .I1(n1033), .I2(donnee[17]), .O(n1068) );
  NAND_GATE U1556 ( .I1(\registres[16][17] ), .I2(n1034), .O(n1067) );
  NAND_GATE U1557 ( .I1(n1069), .I2(n1070), .O(n5257) );
  NAND_GATE U1558 ( .I1(n1033), .I2(donnee[18]), .O(n1070) );
  NAND_GATE U1559 ( .I1(\registres[16][18] ), .I2(n1034), .O(n1069) );
  NAND_GATE U1560 ( .I1(n1071), .I2(n1072), .O(n5258) );
  NAND_GATE U1561 ( .I1(n1033), .I2(donnee[19]), .O(n1072) );
  NAND_GATE U1562 ( .I1(\registres[16][19] ), .I2(n1034), .O(n1071) );
  NAND_GATE U1563 ( .I1(n1073), .I2(n1074), .O(n5259) );
  NAND_GATE U1564 ( .I1(n1033), .I2(donnee[20]), .O(n1074) );
  NAND_GATE U1565 ( .I1(\registres[16][20] ), .I2(n1034), .O(n1073) );
  NAND_GATE U1566 ( .I1(n1075), .I2(n1076), .O(n5260) );
  NAND_GATE U1567 ( .I1(n1033), .I2(donnee[21]), .O(n1076) );
  NAND_GATE U1568 ( .I1(\registres[16][21] ), .I2(n1034), .O(n1075) );
  NAND_GATE U1569 ( .I1(n1077), .I2(n1078), .O(n5261) );
  NAND_GATE U1570 ( .I1(n1033), .I2(donnee[22]), .O(n1078) );
  NAND_GATE U1571 ( .I1(\registres[16][22] ), .I2(n1034), .O(n1077) );
  NAND_GATE U1572 ( .I1(n1079), .I2(n1080), .O(n5262) );
  NAND_GATE U1573 ( .I1(n1033), .I2(donnee[23]), .O(n1080) );
  NAND_GATE U1574 ( .I1(\registres[16][23] ), .I2(n1034), .O(n1079) );
  NAND_GATE U1575 ( .I1(n1081), .I2(n1082), .O(n5263) );
  NAND_GATE U1576 ( .I1(n1033), .I2(donnee[24]), .O(n1082) );
  NAND_GATE U1577 ( .I1(\registres[16][24] ), .I2(n1034), .O(n1081) );
  NAND_GATE U1578 ( .I1(n1083), .I2(n1084), .O(n5264) );
  NAND_GATE U1579 ( .I1(n1033), .I2(donnee[25]), .O(n1084) );
  NAND_GATE U1580 ( .I1(\registres[16][25] ), .I2(n1034), .O(n1083) );
  NAND_GATE U1581 ( .I1(n1085), .I2(n1086), .O(n5265) );
  NAND_GATE U1582 ( .I1(n1033), .I2(donnee[26]), .O(n1086) );
  NAND_GATE U1583 ( .I1(\registres[16][26] ), .I2(n1034), .O(n1085) );
  NAND_GATE U1584 ( .I1(n1087), .I2(n1088), .O(n5266) );
  NAND_GATE U1585 ( .I1(n1033), .I2(donnee[27]), .O(n1088) );
  NAND_GATE U1586 ( .I1(\registres[16][27] ), .I2(n1034), .O(n1087) );
  NAND_GATE U1587 ( .I1(n1089), .I2(n1090), .O(n5267) );
  NAND_GATE U1588 ( .I1(n1033), .I2(donnee[28]), .O(n1090) );
  NAND_GATE U1589 ( .I1(\registres[16][28] ), .I2(n1034), .O(n1089) );
  NAND_GATE U1590 ( .I1(n1091), .I2(n1092), .O(n5268) );
  NAND_GATE U1591 ( .I1(n1033), .I2(donnee[29]), .O(n1092) );
  NAND_GATE U1592 ( .I1(\registres[16][29] ), .I2(n1034), .O(n1091) );
  NAND_GATE U1593 ( .I1(n1093), .I2(n1094), .O(n5269) );
  NAND_GATE U1594 ( .I1(n1033), .I2(donnee[30]), .O(n1094) );
  NAND_GATE U1595 ( .I1(\registres[16][30] ), .I2(n1034), .O(n1093) );
  NAND_GATE U1596 ( .I1(n1095), .I2(n1096), .O(n5270) );
  NAND_GATE U1597 ( .I1(n1033), .I2(donnee[31]), .O(n1096) );
  AND_GATE U1598 ( .I1(n1097), .I2(n1), .O(n1033) );
  NAND_GATE U1599 ( .I1(\registres[16][31] ), .I2(n1034), .O(n1095) );
  NOR_GATE U1600 ( .I1(n1097), .I2(reset), .O(n1034) );
  AND3_GATE U1601 ( .I1(n560), .I2(cmd_ecr), .I3(n628), .O(n1097) );
  NOR_GATE U1602 ( .I1(n2), .I2(reg_dest[3]), .O(n628) );
  NAND_GATE U1603 ( .I1(n1098), .I2(n1099), .O(n5271) );
  NAND_GATE U1604 ( .I1(n1100), .I2(donnee[0]), .O(n1099) );
  NAND_GATE U1605 ( .I1(\registres[15][0] ), .I2(n1101), .O(n1098) );
  NAND_GATE U1606 ( .I1(n1102), .I2(n1103), .O(n5272) );
  NAND_GATE U1607 ( .I1(n1100), .I2(donnee[1]), .O(n1103) );
  NAND_GATE U1608 ( .I1(\registres[15][1] ), .I2(n1101), .O(n1102) );
  NAND_GATE U1609 ( .I1(n1104), .I2(n1105), .O(n5273) );
  NAND_GATE U1610 ( .I1(n1100), .I2(donnee[2]), .O(n1105) );
  NAND_GATE U1611 ( .I1(\registres[15][2] ), .I2(n1101), .O(n1104) );
  NAND_GATE U1612 ( .I1(n1106), .I2(n1107), .O(n5274) );
  NAND_GATE U1613 ( .I1(n1100), .I2(donnee[3]), .O(n1107) );
  NAND_GATE U1614 ( .I1(\registres[15][3] ), .I2(n1101), .O(n1106) );
  NAND_GATE U1615 ( .I1(n1108), .I2(n1109), .O(n5275) );
  NAND_GATE U1616 ( .I1(n1100), .I2(donnee[4]), .O(n1109) );
  NAND_GATE U1617 ( .I1(\registres[15][4] ), .I2(n1101), .O(n1108) );
  NAND_GATE U1618 ( .I1(n1110), .I2(n1111), .O(n5276) );
  NAND_GATE U1619 ( .I1(n1100), .I2(donnee[5]), .O(n1111) );
  NAND_GATE U1620 ( .I1(\registres[15][5] ), .I2(n1101), .O(n1110) );
  NAND_GATE U1621 ( .I1(n1112), .I2(n1113), .O(n5277) );
  NAND_GATE U1622 ( .I1(n1100), .I2(donnee[6]), .O(n1113) );
  NAND_GATE U1623 ( .I1(\registres[15][6] ), .I2(n1101), .O(n1112) );
  NAND_GATE U1624 ( .I1(n1114), .I2(n1115), .O(n5278) );
  NAND_GATE U1625 ( .I1(n1100), .I2(donnee[7]), .O(n1115) );
  NAND_GATE U1626 ( .I1(\registres[15][7] ), .I2(n1101), .O(n1114) );
  NAND_GATE U1627 ( .I1(n1116), .I2(n1117), .O(n5279) );
  NAND_GATE U1628 ( .I1(n1100), .I2(donnee[8]), .O(n1117) );
  NAND_GATE U1629 ( .I1(\registres[15][8] ), .I2(n1101), .O(n1116) );
  NAND_GATE U1630 ( .I1(n1118), .I2(n1119), .O(n5280) );
  NAND_GATE U1631 ( .I1(n1100), .I2(donnee[9]), .O(n1119) );
  NAND_GATE U1632 ( .I1(\registres[15][9] ), .I2(n1101), .O(n1118) );
  NAND_GATE U1633 ( .I1(n1120), .I2(n1121), .O(n5281) );
  NAND_GATE U1634 ( .I1(n1100), .I2(donnee[10]), .O(n1121) );
  NAND_GATE U1635 ( .I1(\registres[15][10] ), .I2(n1101), .O(n1120) );
  NAND_GATE U1636 ( .I1(n1122), .I2(n1123), .O(n5282) );
  NAND_GATE U1637 ( .I1(n1100), .I2(donnee[11]), .O(n1123) );
  NAND_GATE U1638 ( .I1(\registres[15][11] ), .I2(n1101), .O(n1122) );
  NAND_GATE U1639 ( .I1(n1124), .I2(n1125), .O(n5283) );
  NAND_GATE U1640 ( .I1(n1100), .I2(donnee[12]), .O(n1125) );
  NAND_GATE U1641 ( .I1(\registres[15][12] ), .I2(n1101), .O(n1124) );
  NAND_GATE U1642 ( .I1(n1126), .I2(n1127), .O(n5284) );
  NAND_GATE U1643 ( .I1(n1100), .I2(donnee[13]), .O(n1127) );
  NAND_GATE U1644 ( .I1(\registres[15][13] ), .I2(n1101), .O(n1126) );
  NAND_GATE U1645 ( .I1(n1128), .I2(n1129), .O(n5285) );
  NAND_GATE U1646 ( .I1(n1100), .I2(donnee[14]), .O(n1129) );
  NAND_GATE U1647 ( .I1(\registres[15][14] ), .I2(n1101), .O(n1128) );
  NAND_GATE U1648 ( .I1(n1130), .I2(n1131), .O(n5286) );
  NAND_GATE U1649 ( .I1(n1100), .I2(donnee[15]), .O(n1131) );
  NAND_GATE U1650 ( .I1(\registres[15][15] ), .I2(n1101), .O(n1130) );
  NAND_GATE U1651 ( .I1(n1132), .I2(n1133), .O(n5287) );
  NAND_GATE U1652 ( .I1(n1100), .I2(donnee[16]), .O(n1133) );
  NAND_GATE U1653 ( .I1(\registres[15][16] ), .I2(n1101), .O(n1132) );
  NAND_GATE U1654 ( .I1(n1134), .I2(n1135), .O(n5288) );
  NAND_GATE U1655 ( .I1(n1100), .I2(donnee[17]), .O(n1135) );
  NAND_GATE U1656 ( .I1(\registres[15][17] ), .I2(n1101), .O(n1134) );
  NAND_GATE U1657 ( .I1(n1136), .I2(n1137), .O(n5289) );
  NAND_GATE U1658 ( .I1(n1100), .I2(donnee[18]), .O(n1137) );
  NAND_GATE U1659 ( .I1(\registres[15][18] ), .I2(n1101), .O(n1136) );
  NAND_GATE U1660 ( .I1(n1138), .I2(n1139), .O(n5290) );
  NAND_GATE U1661 ( .I1(n1100), .I2(donnee[19]), .O(n1139) );
  NAND_GATE U1662 ( .I1(\registres[15][19] ), .I2(n1101), .O(n1138) );
  NAND_GATE U1663 ( .I1(n1140), .I2(n1141), .O(n5291) );
  NAND_GATE U1664 ( .I1(n1100), .I2(donnee[20]), .O(n1141) );
  NAND_GATE U1665 ( .I1(\registres[15][20] ), .I2(n1101), .O(n1140) );
  NAND_GATE U1666 ( .I1(n1142), .I2(n1143), .O(n5292) );
  NAND_GATE U1667 ( .I1(n1100), .I2(donnee[21]), .O(n1143) );
  NAND_GATE U1668 ( .I1(\registres[15][21] ), .I2(n1101), .O(n1142) );
  NAND_GATE U1669 ( .I1(n1144), .I2(n1145), .O(n5293) );
  NAND_GATE U1670 ( .I1(n1100), .I2(donnee[22]), .O(n1145) );
  NAND_GATE U1671 ( .I1(\registres[15][22] ), .I2(n1101), .O(n1144) );
  NAND_GATE U1672 ( .I1(n1146), .I2(n1147), .O(n5294) );
  NAND_GATE U1673 ( .I1(n1100), .I2(donnee[23]), .O(n1147) );
  NAND_GATE U1674 ( .I1(\registres[15][23] ), .I2(n1101), .O(n1146) );
  NAND_GATE U1675 ( .I1(n1148), .I2(n1149), .O(n5295) );
  NAND_GATE U1676 ( .I1(n1100), .I2(donnee[24]), .O(n1149) );
  NAND_GATE U1677 ( .I1(\registres[15][24] ), .I2(n1101), .O(n1148) );
  NAND_GATE U1678 ( .I1(n1150), .I2(n1151), .O(n5296) );
  NAND_GATE U1679 ( .I1(n1100), .I2(donnee[25]), .O(n1151) );
  NAND_GATE U1680 ( .I1(\registres[15][25] ), .I2(n1101), .O(n1150) );
  NAND_GATE U1681 ( .I1(n1152), .I2(n1153), .O(n5297) );
  NAND_GATE U1682 ( .I1(n1100), .I2(donnee[26]), .O(n1153) );
  NAND_GATE U1683 ( .I1(\registres[15][26] ), .I2(n1101), .O(n1152) );
  NAND_GATE U1684 ( .I1(n1154), .I2(n1155), .O(n5298) );
  NAND_GATE U1685 ( .I1(n1100), .I2(donnee[27]), .O(n1155) );
  NAND_GATE U1686 ( .I1(\registres[15][27] ), .I2(n1101), .O(n1154) );
  NAND_GATE U1687 ( .I1(n1156), .I2(n1157), .O(n5299) );
  NAND_GATE U1688 ( .I1(n1100), .I2(donnee[28]), .O(n1157) );
  NAND_GATE U1689 ( .I1(\registres[15][28] ), .I2(n1101), .O(n1156) );
  NAND_GATE U1690 ( .I1(n1158), .I2(n1159), .O(n5300) );
  NAND_GATE U1691 ( .I1(n1100), .I2(donnee[29]), .O(n1159) );
  NAND_GATE U1692 ( .I1(\registres[15][29] ), .I2(n1101), .O(n1158) );
  NAND_GATE U1693 ( .I1(n1160), .I2(n1161), .O(n5301) );
  NAND_GATE U1694 ( .I1(n1100), .I2(donnee[30]), .O(n1161) );
  NAND_GATE U1695 ( .I1(\registres[15][30] ), .I2(n1101), .O(n1160) );
  NAND_GATE U1696 ( .I1(n1162), .I2(n1163), .O(n5302) );
  NAND_GATE U1697 ( .I1(n1100), .I2(donnee[31]), .O(n1163) );
  AND_GATE U1698 ( .I1(n1164), .I2(n1), .O(n1100) );
  NAND_GATE U1699 ( .I1(\registres[15][31] ), .I2(n1101), .O(n1162) );
  NOR_GATE U1700 ( .I1(n1164), .I2(reset), .O(n1101) );
  AND3_GATE U1701 ( .I1(n84), .I2(cmd_ecr), .I3(n1165), .O(n1164) );
  NAND_GATE U1702 ( .I1(n1166), .I2(n1167), .O(n5303) );
  NAND_GATE U1703 ( .I1(n1168), .I2(donnee[0]), .O(n1167) );
  NAND_GATE U1704 ( .I1(\registres[14][0] ), .I2(n1169), .O(n1166) );
  NAND_GATE U1705 ( .I1(n1170), .I2(n1171), .O(n5304) );
  NAND_GATE U1706 ( .I1(n1168), .I2(donnee[1]), .O(n1171) );
  NAND_GATE U1707 ( .I1(\registres[14][1] ), .I2(n1169), .O(n1170) );
  NAND_GATE U1708 ( .I1(n1172), .I2(n1173), .O(n5305) );
  NAND_GATE U1709 ( .I1(n1168), .I2(donnee[2]), .O(n1173) );
  NAND_GATE U1710 ( .I1(\registres[14][2] ), .I2(n1169), .O(n1172) );
  NAND_GATE U1711 ( .I1(n1174), .I2(n1175), .O(n5306) );
  NAND_GATE U1712 ( .I1(n1168), .I2(donnee[3]), .O(n1175) );
  NAND_GATE U1713 ( .I1(\registres[14][3] ), .I2(n1169), .O(n1174) );
  NAND_GATE U1714 ( .I1(n1176), .I2(n1177), .O(n5307) );
  NAND_GATE U1715 ( .I1(n1168), .I2(donnee[4]), .O(n1177) );
  NAND_GATE U1716 ( .I1(\registres[14][4] ), .I2(n1169), .O(n1176) );
  NAND_GATE U1717 ( .I1(n1178), .I2(n1179), .O(n5308) );
  NAND_GATE U1718 ( .I1(n1168), .I2(donnee[5]), .O(n1179) );
  NAND_GATE U1719 ( .I1(\registres[14][5] ), .I2(n1169), .O(n1178) );
  NAND_GATE U1720 ( .I1(n1180), .I2(n1181), .O(n5309) );
  NAND_GATE U1721 ( .I1(n1168), .I2(donnee[6]), .O(n1181) );
  NAND_GATE U1722 ( .I1(\registres[14][6] ), .I2(n1169), .O(n1180) );
  NAND_GATE U1723 ( .I1(n1182), .I2(n1183), .O(n5310) );
  NAND_GATE U1724 ( .I1(n1168), .I2(donnee[7]), .O(n1183) );
  NAND_GATE U1725 ( .I1(\registres[14][7] ), .I2(n1169), .O(n1182) );
  NAND_GATE U1726 ( .I1(n1184), .I2(n1185), .O(n5311) );
  NAND_GATE U1727 ( .I1(n1168), .I2(donnee[8]), .O(n1185) );
  NAND_GATE U1728 ( .I1(\registres[14][8] ), .I2(n1169), .O(n1184) );
  NAND_GATE U1729 ( .I1(n1186), .I2(n1187), .O(n5312) );
  NAND_GATE U1730 ( .I1(n1168), .I2(donnee[9]), .O(n1187) );
  NAND_GATE U1731 ( .I1(\registres[14][9] ), .I2(n1169), .O(n1186) );
  NAND_GATE U1732 ( .I1(n1188), .I2(n1189), .O(n5313) );
  NAND_GATE U1733 ( .I1(n1168), .I2(donnee[10]), .O(n1189) );
  NAND_GATE U1734 ( .I1(\registres[14][10] ), .I2(n1169), .O(n1188) );
  NAND_GATE U1735 ( .I1(n1190), .I2(n1191), .O(n5314) );
  NAND_GATE U1736 ( .I1(n1168), .I2(donnee[11]), .O(n1191) );
  NAND_GATE U1737 ( .I1(\registres[14][11] ), .I2(n1169), .O(n1190) );
  NAND_GATE U1738 ( .I1(n1192), .I2(n1193), .O(n5315) );
  NAND_GATE U1739 ( .I1(n1168), .I2(donnee[12]), .O(n1193) );
  NAND_GATE U1740 ( .I1(\registres[14][12] ), .I2(n1169), .O(n1192) );
  NAND_GATE U1741 ( .I1(n1194), .I2(n1195), .O(n5316) );
  NAND_GATE U1742 ( .I1(n1168), .I2(donnee[13]), .O(n1195) );
  NAND_GATE U1743 ( .I1(\registres[14][13] ), .I2(n1169), .O(n1194) );
  NAND_GATE U1744 ( .I1(n1196), .I2(n1197), .O(n5317) );
  NAND_GATE U1745 ( .I1(n1168), .I2(donnee[14]), .O(n1197) );
  NAND_GATE U1746 ( .I1(\registres[14][14] ), .I2(n1169), .O(n1196) );
  NAND_GATE U1747 ( .I1(n1198), .I2(n1199), .O(n5318) );
  NAND_GATE U1748 ( .I1(n1168), .I2(donnee[15]), .O(n1199) );
  NAND_GATE U1749 ( .I1(\registres[14][15] ), .I2(n1169), .O(n1198) );
  NAND_GATE U1750 ( .I1(n1200), .I2(n1201), .O(n5319) );
  NAND_GATE U1751 ( .I1(n1168), .I2(donnee[16]), .O(n1201) );
  NAND_GATE U1752 ( .I1(\registres[14][16] ), .I2(n1169), .O(n1200) );
  NAND_GATE U1753 ( .I1(n1202), .I2(n1203), .O(n5320) );
  NAND_GATE U1754 ( .I1(n1168), .I2(donnee[17]), .O(n1203) );
  NAND_GATE U1755 ( .I1(\registres[14][17] ), .I2(n1169), .O(n1202) );
  NAND_GATE U1756 ( .I1(n1204), .I2(n1205), .O(n5321) );
  NAND_GATE U1757 ( .I1(n1168), .I2(donnee[18]), .O(n1205) );
  NAND_GATE U1758 ( .I1(\registres[14][18] ), .I2(n1169), .O(n1204) );
  NAND_GATE U1759 ( .I1(n1206), .I2(n1207), .O(n5322) );
  NAND_GATE U1760 ( .I1(n1168), .I2(donnee[19]), .O(n1207) );
  NAND_GATE U1761 ( .I1(\registres[14][19] ), .I2(n1169), .O(n1206) );
  NAND_GATE U1762 ( .I1(n1208), .I2(n1209), .O(n5323) );
  NAND_GATE U1763 ( .I1(n1168), .I2(donnee[20]), .O(n1209) );
  NAND_GATE U1764 ( .I1(\registres[14][20] ), .I2(n1169), .O(n1208) );
  NAND_GATE U1765 ( .I1(n1210), .I2(n1211), .O(n5324) );
  NAND_GATE U1766 ( .I1(n1168), .I2(donnee[21]), .O(n1211) );
  NAND_GATE U1767 ( .I1(\registres[14][21] ), .I2(n1169), .O(n1210) );
  NAND_GATE U1768 ( .I1(n1212), .I2(n1213), .O(n5325) );
  NAND_GATE U1769 ( .I1(n1168), .I2(donnee[22]), .O(n1213) );
  NAND_GATE U1770 ( .I1(\registres[14][22] ), .I2(n1169), .O(n1212) );
  NAND_GATE U1771 ( .I1(n1214), .I2(n1215), .O(n5326) );
  NAND_GATE U1772 ( .I1(n1168), .I2(donnee[23]), .O(n1215) );
  NAND_GATE U1773 ( .I1(\registres[14][23] ), .I2(n1169), .O(n1214) );
  NAND_GATE U1774 ( .I1(n1216), .I2(n1217), .O(n5327) );
  NAND_GATE U1775 ( .I1(n1168), .I2(donnee[24]), .O(n1217) );
  NAND_GATE U1776 ( .I1(\registres[14][24] ), .I2(n1169), .O(n1216) );
  NAND_GATE U1777 ( .I1(n1218), .I2(n1219), .O(n5328) );
  NAND_GATE U1778 ( .I1(n1168), .I2(donnee[25]), .O(n1219) );
  NAND_GATE U1779 ( .I1(\registres[14][25] ), .I2(n1169), .O(n1218) );
  NAND_GATE U1780 ( .I1(n1220), .I2(n1221), .O(n5329) );
  NAND_GATE U1781 ( .I1(n1168), .I2(donnee[26]), .O(n1221) );
  NAND_GATE U1782 ( .I1(\registres[14][26] ), .I2(n1169), .O(n1220) );
  NAND_GATE U1783 ( .I1(n1222), .I2(n1223), .O(n5330) );
  NAND_GATE U1784 ( .I1(n1168), .I2(donnee[27]), .O(n1223) );
  NAND_GATE U1785 ( .I1(\registres[14][27] ), .I2(n1169), .O(n1222) );
  NAND_GATE U1786 ( .I1(n1224), .I2(n1225), .O(n5331) );
  NAND_GATE U1787 ( .I1(n1168), .I2(donnee[28]), .O(n1225) );
  NAND_GATE U1788 ( .I1(\registres[14][28] ), .I2(n1169), .O(n1224) );
  NAND_GATE U1789 ( .I1(n1226), .I2(n1227), .O(n5332) );
  NAND_GATE U1790 ( .I1(n1168), .I2(donnee[29]), .O(n1227) );
  NAND_GATE U1791 ( .I1(\registres[14][29] ), .I2(n1169), .O(n1226) );
  NAND_GATE U1792 ( .I1(n1228), .I2(n1229), .O(n5333) );
  NAND_GATE U1793 ( .I1(n1168), .I2(donnee[30]), .O(n1229) );
  NAND_GATE U1794 ( .I1(\registres[14][30] ), .I2(n1169), .O(n1228) );
  NAND_GATE U1795 ( .I1(n1230), .I2(n1231), .O(n5334) );
  NAND_GATE U1796 ( .I1(n1168), .I2(donnee[31]), .O(n1231) );
  AND_GATE U1797 ( .I1(n1232), .I2(n1), .O(n1168) );
  NAND_GATE U1798 ( .I1(\registres[14][31] ), .I2(n1169), .O(n1230) );
  NOR_GATE U1799 ( .I1(n1232), .I2(reset), .O(n1169) );
  AND3_GATE U1800 ( .I1(n152), .I2(cmd_ecr), .I3(n1165), .O(n1232) );
  NAND_GATE U1801 ( .I1(n1233), .I2(n1234), .O(n5335) );
  NAND_GATE U1802 ( .I1(n1235), .I2(donnee[0]), .O(n1234) );
  NAND_GATE U1803 ( .I1(\registres[13][0] ), .I2(n1236), .O(n1233) );
  NAND_GATE U1804 ( .I1(n1237), .I2(n1238), .O(n5336) );
  NAND_GATE U1805 ( .I1(n1235), .I2(donnee[1]), .O(n1238) );
  NAND_GATE U1806 ( .I1(\registres[13][1] ), .I2(n1236), .O(n1237) );
  NAND_GATE U1807 ( .I1(n1239), .I2(n1240), .O(n5337) );
  NAND_GATE U1808 ( .I1(n1235), .I2(donnee[2]), .O(n1240) );
  NAND_GATE U1809 ( .I1(\registres[13][2] ), .I2(n1236), .O(n1239) );
  NAND_GATE U1810 ( .I1(n1241), .I2(n1242), .O(n5338) );
  NAND_GATE U1811 ( .I1(n1235), .I2(donnee[3]), .O(n1242) );
  NAND_GATE U1812 ( .I1(\registres[13][3] ), .I2(n1236), .O(n1241) );
  NAND_GATE U1813 ( .I1(n1243), .I2(n1244), .O(n5339) );
  NAND_GATE U1814 ( .I1(n1235), .I2(donnee[4]), .O(n1244) );
  NAND_GATE U1815 ( .I1(\registres[13][4] ), .I2(n1236), .O(n1243) );
  NAND_GATE U1816 ( .I1(n1245), .I2(n1246), .O(n5340) );
  NAND_GATE U1817 ( .I1(n1235), .I2(donnee[5]), .O(n1246) );
  NAND_GATE U1818 ( .I1(\registres[13][5] ), .I2(n1236), .O(n1245) );
  NAND_GATE U1819 ( .I1(n1247), .I2(n1248), .O(n5341) );
  NAND_GATE U1820 ( .I1(n1235), .I2(donnee[6]), .O(n1248) );
  NAND_GATE U1821 ( .I1(\registres[13][6] ), .I2(n1236), .O(n1247) );
  NAND_GATE U1822 ( .I1(n1249), .I2(n1250), .O(n5342) );
  NAND_GATE U1823 ( .I1(n1235), .I2(donnee[7]), .O(n1250) );
  NAND_GATE U1824 ( .I1(\registres[13][7] ), .I2(n1236), .O(n1249) );
  NAND_GATE U1825 ( .I1(n1251), .I2(n1252), .O(n5343) );
  NAND_GATE U1826 ( .I1(n1235), .I2(donnee[8]), .O(n1252) );
  NAND_GATE U1827 ( .I1(\registres[13][8] ), .I2(n1236), .O(n1251) );
  NAND_GATE U1828 ( .I1(n1253), .I2(n1254), .O(n5344) );
  NAND_GATE U1829 ( .I1(n1235), .I2(donnee[9]), .O(n1254) );
  NAND_GATE U1830 ( .I1(\registres[13][9] ), .I2(n1236), .O(n1253) );
  NAND_GATE U1831 ( .I1(n1255), .I2(n1256), .O(n5345) );
  NAND_GATE U1832 ( .I1(n1235), .I2(donnee[10]), .O(n1256) );
  NAND_GATE U1833 ( .I1(\registres[13][10] ), .I2(n1236), .O(n1255) );
  NAND_GATE U1834 ( .I1(n1257), .I2(n1258), .O(n5346) );
  NAND_GATE U1835 ( .I1(n1235), .I2(donnee[11]), .O(n1258) );
  NAND_GATE U1836 ( .I1(\registres[13][11] ), .I2(n1236), .O(n1257) );
  NAND_GATE U1837 ( .I1(n1259), .I2(n1260), .O(n5347) );
  NAND_GATE U1838 ( .I1(n1235), .I2(donnee[12]), .O(n1260) );
  NAND_GATE U1839 ( .I1(\registres[13][12] ), .I2(n1236), .O(n1259) );
  NAND_GATE U1840 ( .I1(n1261), .I2(n1262), .O(n5348) );
  NAND_GATE U1841 ( .I1(n1235), .I2(donnee[13]), .O(n1262) );
  NAND_GATE U1842 ( .I1(\registres[13][13] ), .I2(n1236), .O(n1261) );
  NAND_GATE U1843 ( .I1(n1263), .I2(n1264), .O(n5349) );
  NAND_GATE U1844 ( .I1(n1235), .I2(donnee[14]), .O(n1264) );
  NAND_GATE U1845 ( .I1(\registres[13][14] ), .I2(n1236), .O(n1263) );
  NAND_GATE U1846 ( .I1(n1265), .I2(n1266), .O(n5350) );
  NAND_GATE U1847 ( .I1(n1235), .I2(donnee[15]), .O(n1266) );
  NAND_GATE U1848 ( .I1(\registres[13][15] ), .I2(n1236), .O(n1265) );
  NAND_GATE U1849 ( .I1(n1267), .I2(n1268), .O(n5351) );
  NAND_GATE U1850 ( .I1(n1235), .I2(donnee[16]), .O(n1268) );
  NAND_GATE U1851 ( .I1(\registres[13][16] ), .I2(n1236), .O(n1267) );
  NAND_GATE U1852 ( .I1(n1269), .I2(n1270), .O(n5352) );
  NAND_GATE U1853 ( .I1(n1235), .I2(donnee[17]), .O(n1270) );
  NAND_GATE U1854 ( .I1(\registres[13][17] ), .I2(n1236), .O(n1269) );
  NAND_GATE U1855 ( .I1(n1271), .I2(n1272), .O(n5353) );
  NAND_GATE U1856 ( .I1(n1235), .I2(donnee[18]), .O(n1272) );
  NAND_GATE U1857 ( .I1(\registres[13][18] ), .I2(n1236), .O(n1271) );
  NAND_GATE U1858 ( .I1(n1273), .I2(n1274), .O(n5354) );
  NAND_GATE U1859 ( .I1(n1235), .I2(donnee[19]), .O(n1274) );
  NAND_GATE U1860 ( .I1(\registres[13][19] ), .I2(n1236), .O(n1273) );
  NAND_GATE U1861 ( .I1(n1275), .I2(n1276), .O(n5355) );
  NAND_GATE U1862 ( .I1(n1235), .I2(donnee[20]), .O(n1276) );
  NAND_GATE U1863 ( .I1(\registres[13][20] ), .I2(n1236), .O(n1275) );
  NAND_GATE U1864 ( .I1(n1277), .I2(n1278), .O(n5356) );
  NAND_GATE U1865 ( .I1(n1235), .I2(donnee[21]), .O(n1278) );
  NAND_GATE U1866 ( .I1(\registres[13][21] ), .I2(n1236), .O(n1277) );
  NAND_GATE U1867 ( .I1(n1279), .I2(n1280), .O(n5357) );
  NAND_GATE U1868 ( .I1(n1235), .I2(donnee[22]), .O(n1280) );
  NAND_GATE U1869 ( .I1(\registres[13][22] ), .I2(n1236), .O(n1279) );
  NAND_GATE U1870 ( .I1(n1281), .I2(n1282), .O(n5358) );
  NAND_GATE U1871 ( .I1(n1235), .I2(donnee[23]), .O(n1282) );
  NAND_GATE U1872 ( .I1(\registres[13][23] ), .I2(n1236), .O(n1281) );
  NAND_GATE U1873 ( .I1(n1283), .I2(n1284), .O(n5359) );
  NAND_GATE U1874 ( .I1(n1235), .I2(donnee[24]), .O(n1284) );
  NAND_GATE U1875 ( .I1(\registres[13][24] ), .I2(n1236), .O(n1283) );
  NAND_GATE U1876 ( .I1(n1285), .I2(n1286), .O(n5360) );
  NAND_GATE U1877 ( .I1(n1235), .I2(donnee[25]), .O(n1286) );
  NAND_GATE U1878 ( .I1(\registres[13][25] ), .I2(n1236), .O(n1285) );
  NAND_GATE U1879 ( .I1(n1287), .I2(n1288), .O(n5361) );
  NAND_GATE U1880 ( .I1(n1235), .I2(donnee[26]), .O(n1288) );
  NAND_GATE U1881 ( .I1(\registres[13][26] ), .I2(n1236), .O(n1287) );
  NAND_GATE U1882 ( .I1(n1289), .I2(n1290), .O(n5362) );
  NAND_GATE U1883 ( .I1(n1235), .I2(donnee[27]), .O(n1290) );
  NAND_GATE U1884 ( .I1(\registres[13][27] ), .I2(n1236), .O(n1289) );
  NAND_GATE U1885 ( .I1(n1291), .I2(n1292), .O(n5363) );
  NAND_GATE U1886 ( .I1(n1235), .I2(donnee[28]), .O(n1292) );
  NAND_GATE U1887 ( .I1(\registres[13][28] ), .I2(n1236), .O(n1291) );
  NAND_GATE U1888 ( .I1(n1293), .I2(n1294), .O(n5364) );
  NAND_GATE U1889 ( .I1(n1235), .I2(donnee[29]), .O(n1294) );
  NAND_GATE U1890 ( .I1(\registres[13][29] ), .I2(n1236), .O(n1293) );
  NAND_GATE U1891 ( .I1(n1295), .I2(n1296), .O(n5365) );
  NAND_GATE U1892 ( .I1(n1235), .I2(donnee[30]), .O(n1296) );
  NAND_GATE U1893 ( .I1(\registres[13][30] ), .I2(n1236), .O(n1295) );
  NAND_GATE U1894 ( .I1(n1297), .I2(n1298), .O(n5366) );
  NAND_GATE U1895 ( .I1(n1235), .I2(donnee[31]), .O(n1298) );
  AND_GATE U1896 ( .I1(n1299), .I2(n1), .O(n1235) );
  NAND_GATE U1897 ( .I1(\registres[13][31] ), .I2(n1236), .O(n1297) );
  NOR_GATE U1898 ( .I1(n1299), .I2(reset), .O(n1236) );
  AND3_GATE U1899 ( .I1(n220), .I2(cmd_ecr), .I3(n1165), .O(n1299) );
  NAND_GATE U1900 ( .I1(n1300), .I2(n1301), .O(n5367) );
  NAND_GATE U1901 ( .I1(n1302), .I2(donnee[0]), .O(n1301) );
  NAND_GATE U1902 ( .I1(\registres[12][0] ), .I2(n1303), .O(n1300) );
  NAND_GATE U1903 ( .I1(n1304), .I2(n1305), .O(n5368) );
  NAND_GATE U1904 ( .I1(n1302), .I2(donnee[1]), .O(n1305) );
  NAND_GATE U1905 ( .I1(\registres[12][1] ), .I2(n1303), .O(n1304) );
  NAND_GATE U1906 ( .I1(n1306), .I2(n1307), .O(n5369) );
  NAND_GATE U1907 ( .I1(n1302), .I2(donnee[2]), .O(n1307) );
  NAND_GATE U1908 ( .I1(\registres[12][2] ), .I2(n1303), .O(n1306) );
  NAND_GATE U1909 ( .I1(n1308), .I2(n1309), .O(n5370) );
  NAND_GATE U1910 ( .I1(n1302), .I2(donnee[3]), .O(n1309) );
  NAND_GATE U1911 ( .I1(\registres[12][3] ), .I2(n1303), .O(n1308) );
  NAND_GATE U1912 ( .I1(n1310), .I2(n1311), .O(n5371) );
  NAND_GATE U1913 ( .I1(n1302), .I2(donnee[4]), .O(n1311) );
  NAND_GATE U1914 ( .I1(\registres[12][4] ), .I2(n1303), .O(n1310) );
  NAND_GATE U1915 ( .I1(n1312), .I2(n1313), .O(n5372) );
  NAND_GATE U1916 ( .I1(n1302), .I2(donnee[5]), .O(n1313) );
  NAND_GATE U1917 ( .I1(\registres[12][5] ), .I2(n1303), .O(n1312) );
  NAND_GATE U1918 ( .I1(n1314), .I2(n1315), .O(n5373) );
  NAND_GATE U1919 ( .I1(n1302), .I2(donnee[6]), .O(n1315) );
  NAND_GATE U1920 ( .I1(\registres[12][6] ), .I2(n1303), .O(n1314) );
  NAND_GATE U1921 ( .I1(n1316), .I2(n1317), .O(n5374) );
  NAND_GATE U1922 ( .I1(n1302), .I2(donnee[7]), .O(n1317) );
  NAND_GATE U1923 ( .I1(\registres[12][7] ), .I2(n1303), .O(n1316) );
  NAND_GATE U1924 ( .I1(n1318), .I2(n1319), .O(n5375) );
  NAND_GATE U1925 ( .I1(n1302), .I2(donnee[8]), .O(n1319) );
  NAND_GATE U1926 ( .I1(\registres[12][8] ), .I2(n1303), .O(n1318) );
  NAND_GATE U1927 ( .I1(n1320), .I2(n1321), .O(n5376) );
  NAND_GATE U1928 ( .I1(n1302), .I2(donnee[9]), .O(n1321) );
  NAND_GATE U1929 ( .I1(\registres[12][9] ), .I2(n1303), .O(n1320) );
  NAND_GATE U1930 ( .I1(n1322), .I2(n1323), .O(n5377) );
  NAND_GATE U1931 ( .I1(n1302), .I2(donnee[10]), .O(n1323) );
  NAND_GATE U1932 ( .I1(\registres[12][10] ), .I2(n1303), .O(n1322) );
  NAND_GATE U1933 ( .I1(n1324), .I2(n1325), .O(n5378) );
  NAND_GATE U1934 ( .I1(n1302), .I2(donnee[11]), .O(n1325) );
  NAND_GATE U1935 ( .I1(\registres[12][11] ), .I2(n1303), .O(n1324) );
  NAND_GATE U1936 ( .I1(n1326), .I2(n1327), .O(n5379) );
  NAND_GATE U1937 ( .I1(n1302), .I2(donnee[12]), .O(n1327) );
  NAND_GATE U1938 ( .I1(\registres[12][12] ), .I2(n1303), .O(n1326) );
  NAND_GATE U1939 ( .I1(n1328), .I2(n1329), .O(n5380) );
  NAND_GATE U1940 ( .I1(n1302), .I2(donnee[13]), .O(n1329) );
  NAND_GATE U1941 ( .I1(\registres[12][13] ), .I2(n1303), .O(n1328) );
  NAND_GATE U1942 ( .I1(n1330), .I2(n1331), .O(n5381) );
  NAND_GATE U1943 ( .I1(n1302), .I2(donnee[14]), .O(n1331) );
  NAND_GATE U1944 ( .I1(\registres[12][14] ), .I2(n1303), .O(n1330) );
  NAND_GATE U1945 ( .I1(n1332), .I2(n1333), .O(n5382) );
  NAND_GATE U1946 ( .I1(n1302), .I2(donnee[15]), .O(n1333) );
  NAND_GATE U1947 ( .I1(\registres[12][15] ), .I2(n1303), .O(n1332) );
  NAND_GATE U1948 ( .I1(n1334), .I2(n1335), .O(n5383) );
  NAND_GATE U1949 ( .I1(n1302), .I2(donnee[16]), .O(n1335) );
  NAND_GATE U1950 ( .I1(\registres[12][16] ), .I2(n1303), .O(n1334) );
  NAND_GATE U1951 ( .I1(n1336), .I2(n1337), .O(n5384) );
  NAND_GATE U1952 ( .I1(n1302), .I2(donnee[17]), .O(n1337) );
  NAND_GATE U1953 ( .I1(\registres[12][17] ), .I2(n1303), .O(n1336) );
  NAND_GATE U1954 ( .I1(n1338), .I2(n1339), .O(n5385) );
  NAND_GATE U1955 ( .I1(n1302), .I2(donnee[18]), .O(n1339) );
  NAND_GATE U1956 ( .I1(\registres[12][18] ), .I2(n1303), .O(n1338) );
  NAND_GATE U1957 ( .I1(n1340), .I2(n1341), .O(n5386) );
  NAND_GATE U1958 ( .I1(n1302), .I2(donnee[19]), .O(n1341) );
  NAND_GATE U1959 ( .I1(\registres[12][19] ), .I2(n1303), .O(n1340) );
  NAND_GATE U1960 ( .I1(n1342), .I2(n1343), .O(n5387) );
  NAND_GATE U1961 ( .I1(n1302), .I2(donnee[20]), .O(n1343) );
  NAND_GATE U1962 ( .I1(\registres[12][20] ), .I2(n1303), .O(n1342) );
  NAND_GATE U1963 ( .I1(n1344), .I2(n1345), .O(n5388) );
  NAND_GATE U1964 ( .I1(n1302), .I2(donnee[21]), .O(n1345) );
  NAND_GATE U1965 ( .I1(\registres[12][21] ), .I2(n1303), .O(n1344) );
  NAND_GATE U1966 ( .I1(n1346), .I2(n1347), .O(n5389) );
  NAND_GATE U1967 ( .I1(n1302), .I2(donnee[22]), .O(n1347) );
  NAND_GATE U1968 ( .I1(\registres[12][22] ), .I2(n1303), .O(n1346) );
  NAND_GATE U1969 ( .I1(n1348), .I2(n1349), .O(n5390) );
  NAND_GATE U1970 ( .I1(n1302), .I2(donnee[23]), .O(n1349) );
  NAND_GATE U1971 ( .I1(\registres[12][23] ), .I2(n1303), .O(n1348) );
  NAND_GATE U1972 ( .I1(n1350), .I2(n1351), .O(n5391) );
  NAND_GATE U1973 ( .I1(n1302), .I2(donnee[24]), .O(n1351) );
  NAND_GATE U1974 ( .I1(\registres[12][24] ), .I2(n1303), .O(n1350) );
  NAND_GATE U1975 ( .I1(n1352), .I2(n1353), .O(n5392) );
  NAND_GATE U1976 ( .I1(n1302), .I2(donnee[25]), .O(n1353) );
  NAND_GATE U1977 ( .I1(\registres[12][25] ), .I2(n1303), .O(n1352) );
  NAND_GATE U1978 ( .I1(n1354), .I2(n1355), .O(n5393) );
  NAND_GATE U1979 ( .I1(n1302), .I2(donnee[26]), .O(n1355) );
  NAND_GATE U1980 ( .I1(\registres[12][26] ), .I2(n1303), .O(n1354) );
  NAND_GATE U1981 ( .I1(n1356), .I2(n1357), .O(n5394) );
  NAND_GATE U1982 ( .I1(n1302), .I2(donnee[27]), .O(n1357) );
  NAND_GATE U1983 ( .I1(\registres[12][27] ), .I2(n1303), .O(n1356) );
  NAND_GATE U1984 ( .I1(n1358), .I2(n1359), .O(n5395) );
  NAND_GATE U1985 ( .I1(n1302), .I2(donnee[28]), .O(n1359) );
  NAND_GATE U1986 ( .I1(\registres[12][28] ), .I2(n1303), .O(n1358) );
  NAND_GATE U1987 ( .I1(n1360), .I2(n1361), .O(n5396) );
  NAND_GATE U1988 ( .I1(n1302), .I2(donnee[29]), .O(n1361) );
  NAND_GATE U1989 ( .I1(\registres[12][29] ), .I2(n1303), .O(n1360) );
  NAND_GATE U1990 ( .I1(n1362), .I2(n1363), .O(n5397) );
  NAND_GATE U1991 ( .I1(n1302), .I2(donnee[30]), .O(n1363) );
  NAND_GATE U1992 ( .I1(\registres[12][30] ), .I2(n1303), .O(n1362) );
  NAND_GATE U1993 ( .I1(n1364), .I2(n1365), .O(n5398) );
  NAND_GATE U1994 ( .I1(n1302), .I2(donnee[31]), .O(n1365) );
  AND_GATE U1995 ( .I1(n1366), .I2(n1), .O(n1302) );
  NAND_GATE U1996 ( .I1(\registres[12][31] ), .I2(n1303), .O(n1364) );
  NOR_GATE U1997 ( .I1(n1366), .I2(reset), .O(n1303) );
  AND3_GATE U1998 ( .I1(n288), .I2(cmd_ecr), .I3(n1165), .O(n1366) );
  NAND_GATE U1999 ( .I1(n1367), .I2(n1368), .O(n5399) );
  NAND_GATE U2000 ( .I1(n1369), .I2(donnee[0]), .O(n1368) );
  NAND_GATE U2001 ( .I1(\registres[11][0] ), .I2(n1370), .O(n1367) );
  NAND_GATE U2002 ( .I1(n1371), .I2(n1372), .O(n5400) );
  NAND_GATE U2003 ( .I1(n1369), .I2(donnee[1]), .O(n1372) );
  NAND_GATE U2004 ( .I1(\registres[11][1] ), .I2(n1370), .O(n1371) );
  NAND_GATE U2005 ( .I1(n1373), .I2(n1374), .O(n5401) );
  NAND_GATE U2006 ( .I1(n1369), .I2(donnee[2]), .O(n1374) );
  NAND_GATE U2007 ( .I1(\registres[11][2] ), .I2(n1370), .O(n1373) );
  NAND_GATE U2008 ( .I1(n1375), .I2(n1376), .O(n5402) );
  NAND_GATE U2009 ( .I1(n1369), .I2(donnee[3]), .O(n1376) );
  NAND_GATE U2010 ( .I1(\registres[11][3] ), .I2(n1370), .O(n1375) );
  NAND_GATE U2011 ( .I1(n1377), .I2(n1378), .O(n5403) );
  NAND_GATE U2012 ( .I1(n1369), .I2(donnee[4]), .O(n1378) );
  NAND_GATE U2013 ( .I1(\registres[11][4] ), .I2(n1370), .O(n1377) );
  NAND_GATE U2014 ( .I1(n1379), .I2(n1380), .O(n5404) );
  NAND_GATE U2015 ( .I1(n1369), .I2(donnee[5]), .O(n1380) );
  NAND_GATE U2016 ( .I1(\registres[11][5] ), .I2(n1370), .O(n1379) );
  NAND_GATE U2017 ( .I1(n1381), .I2(n1382), .O(n5405) );
  NAND_GATE U2018 ( .I1(n1369), .I2(donnee[6]), .O(n1382) );
  NAND_GATE U2019 ( .I1(\registres[11][6] ), .I2(n1370), .O(n1381) );
  NAND_GATE U2020 ( .I1(n1383), .I2(n1384), .O(n5406) );
  NAND_GATE U2021 ( .I1(n1369), .I2(donnee[7]), .O(n1384) );
  NAND_GATE U2022 ( .I1(\registres[11][7] ), .I2(n1370), .O(n1383) );
  NAND_GATE U2023 ( .I1(n1385), .I2(n1386), .O(n5407) );
  NAND_GATE U2024 ( .I1(n1369), .I2(donnee[8]), .O(n1386) );
  NAND_GATE U2025 ( .I1(\registres[11][8] ), .I2(n1370), .O(n1385) );
  NAND_GATE U2026 ( .I1(n1387), .I2(n1388), .O(n5408) );
  NAND_GATE U2027 ( .I1(n1369), .I2(donnee[9]), .O(n1388) );
  NAND_GATE U2028 ( .I1(\registres[11][9] ), .I2(n1370), .O(n1387) );
  NAND_GATE U2029 ( .I1(n1389), .I2(n1390), .O(n5409) );
  NAND_GATE U2030 ( .I1(n1369), .I2(donnee[10]), .O(n1390) );
  NAND_GATE U2031 ( .I1(\registres[11][10] ), .I2(n1370), .O(n1389) );
  NAND_GATE U2032 ( .I1(n1391), .I2(n1392), .O(n5410) );
  NAND_GATE U2033 ( .I1(n1369), .I2(donnee[11]), .O(n1392) );
  NAND_GATE U2034 ( .I1(\registres[11][11] ), .I2(n1370), .O(n1391) );
  NAND_GATE U2035 ( .I1(n1393), .I2(n1394), .O(n5411) );
  NAND_GATE U2036 ( .I1(n1369), .I2(donnee[12]), .O(n1394) );
  NAND_GATE U2037 ( .I1(\registres[11][12] ), .I2(n1370), .O(n1393) );
  NAND_GATE U2038 ( .I1(n1395), .I2(n1396), .O(n5412) );
  NAND_GATE U2039 ( .I1(n1369), .I2(donnee[13]), .O(n1396) );
  NAND_GATE U2040 ( .I1(\registres[11][13] ), .I2(n1370), .O(n1395) );
  NAND_GATE U2041 ( .I1(n1397), .I2(n1398), .O(n5413) );
  NAND_GATE U2042 ( .I1(n1369), .I2(donnee[14]), .O(n1398) );
  NAND_GATE U2043 ( .I1(\registres[11][14] ), .I2(n1370), .O(n1397) );
  NAND_GATE U2044 ( .I1(n1399), .I2(n1400), .O(n5414) );
  NAND_GATE U2045 ( .I1(n1369), .I2(donnee[15]), .O(n1400) );
  NAND_GATE U2046 ( .I1(\registres[11][15] ), .I2(n1370), .O(n1399) );
  NAND_GATE U2047 ( .I1(n1401), .I2(n1402), .O(n5415) );
  NAND_GATE U2048 ( .I1(n1369), .I2(donnee[16]), .O(n1402) );
  NAND_GATE U2049 ( .I1(\registres[11][16] ), .I2(n1370), .O(n1401) );
  NAND_GATE U2050 ( .I1(n1403), .I2(n1404), .O(n5416) );
  NAND_GATE U2051 ( .I1(n1369), .I2(donnee[17]), .O(n1404) );
  NAND_GATE U2052 ( .I1(\registres[11][17] ), .I2(n1370), .O(n1403) );
  NAND_GATE U2053 ( .I1(n1405), .I2(n1406), .O(n5417) );
  NAND_GATE U2054 ( .I1(n1369), .I2(donnee[18]), .O(n1406) );
  NAND_GATE U2055 ( .I1(\registres[11][18] ), .I2(n1370), .O(n1405) );
  NAND_GATE U2056 ( .I1(n1407), .I2(n1408), .O(n5418) );
  NAND_GATE U2057 ( .I1(n1369), .I2(donnee[19]), .O(n1408) );
  NAND_GATE U2058 ( .I1(\registres[11][19] ), .I2(n1370), .O(n1407) );
  NAND_GATE U2059 ( .I1(n1409), .I2(n1410), .O(n5419) );
  NAND_GATE U2060 ( .I1(n1369), .I2(donnee[20]), .O(n1410) );
  NAND_GATE U2061 ( .I1(\registres[11][20] ), .I2(n1370), .O(n1409) );
  NAND_GATE U2062 ( .I1(n1411), .I2(n1412), .O(n5420) );
  NAND_GATE U2063 ( .I1(n1369), .I2(donnee[21]), .O(n1412) );
  NAND_GATE U2064 ( .I1(\registres[11][21] ), .I2(n1370), .O(n1411) );
  NAND_GATE U2065 ( .I1(n1413), .I2(n1414), .O(n5421) );
  NAND_GATE U2066 ( .I1(n1369), .I2(donnee[22]), .O(n1414) );
  NAND_GATE U2067 ( .I1(\registres[11][22] ), .I2(n1370), .O(n1413) );
  NAND_GATE U2068 ( .I1(n1415), .I2(n1416), .O(n5422) );
  NAND_GATE U2069 ( .I1(n1369), .I2(donnee[23]), .O(n1416) );
  NAND_GATE U2070 ( .I1(\registres[11][23] ), .I2(n1370), .O(n1415) );
  NAND_GATE U2071 ( .I1(n1417), .I2(n1418), .O(n5423) );
  NAND_GATE U2072 ( .I1(n1369), .I2(donnee[24]), .O(n1418) );
  NAND_GATE U2073 ( .I1(\registres[11][24] ), .I2(n1370), .O(n1417) );
  NAND_GATE U2074 ( .I1(n1419), .I2(n1420), .O(n5424) );
  NAND_GATE U2075 ( .I1(n1369), .I2(donnee[25]), .O(n1420) );
  NAND_GATE U2076 ( .I1(\registres[11][25] ), .I2(n1370), .O(n1419) );
  NAND_GATE U2077 ( .I1(n1421), .I2(n1422), .O(n5425) );
  NAND_GATE U2078 ( .I1(n1369), .I2(donnee[26]), .O(n1422) );
  NAND_GATE U2079 ( .I1(\registres[11][26] ), .I2(n1370), .O(n1421) );
  NAND_GATE U2080 ( .I1(n1423), .I2(n1424), .O(n5426) );
  NAND_GATE U2081 ( .I1(n1369), .I2(donnee[27]), .O(n1424) );
  NAND_GATE U2082 ( .I1(\registres[11][27] ), .I2(n1370), .O(n1423) );
  NAND_GATE U2083 ( .I1(n1425), .I2(n1426), .O(n5427) );
  NAND_GATE U2084 ( .I1(n1369), .I2(donnee[28]), .O(n1426) );
  NAND_GATE U2085 ( .I1(\registres[11][28] ), .I2(n1370), .O(n1425) );
  NAND_GATE U2086 ( .I1(n1427), .I2(n1428), .O(n5428) );
  NAND_GATE U2087 ( .I1(n1369), .I2(donnee[29]), .O(n1428) );
  NAND_GATE U2088 ( .I1(\registres[11][29] ), .I2(n1370), .O(n1427) );
  NAND_GATE U2089 ( .I1(n1429), .I2(n1430), .O(n5429) );
  NAND_GATE U2090 ( .I1(n1369), .I2(donnee[30]), .O(n1430) );
  NAND_GATE U2091 ( .I1(\registres[11][30] ), .I2(n1370), .O(n1429) );
  NAND_GATE U2092 ( .I1(n1431), .I2(n1432), .O(n5430) );
  NAND_GATE U2093 ( .I1(n1369), .I2(donnee[31]), .O(n1432) );
  AND_GATE U2094 ( .I1(n1433), .I2(n1), .O(n1369) );
  NAND_GATE U2095 ( .I1(\registres[11][31] ), .I2(n1370), .O(n1431) );
  NOR_GATE U2096 ( .I1(n1433), .I2(reset), .O(n1370) );
  AND3_GATE U2097 ( .I1(n356), .I2(cmd_ecr), .I3(n1165), .O(n1433) );
  NAND_GATE U2098 ( .I1(n1434), .I2(n1435), .O(n5431) );
  NAND_GATE U2099 ( .I1(n1436), .I2(donnee[0]), .O(n1435) );
  NAND_GATE U2100 ( .I1(\registres[10][0] ), .I2(n1437), .O(n1434) );
  NAND_GATE U2101 ( .I1(n1438), .I2(n1439), .O(n5432) );
  NAND_GATE U2102 ( .I1(n1436), .I2(donnee[1]), .O(n1439) );
  NAND_GATE U2103 ( .I1(\registres[10][1] ), .I2(n1437), .O(n1438) );
  NAND_GATE U2104 ( .I1(n1440), .I2(n1441), .O(n5433) );
  NAND_GATE U2105 ( .I1(n1436), .I2(donnee[2]), .O(n1441) );
  NAND_GATE U2106 ( .I1(\registres[10][2] ), .I2(n1437), .O(n1440) );
  NAND_GATE U2107 ( .I1(n1442), .I2(n1443), .O(n5434) );
  NAND_GATE U2108 ( .I1(n1436), .I2(donnee[3]), .O(n1443) );
  NAND_GATE U2109 ( .I1(\registres[10][3] ), .I2(n1437), .O(n1442) );
  NAND_GATE U2110 ( .I1(n1444), .I2(n1445), .O(n5435) );
  NAND_GATE U2111 ( .I1(n1436), .I2(donnee[4]), .O(n1445) );
  NAND_GATE U2112 ( .I1(\registres[10][4] ), .I2(n1437), .O(n1444) );
  NAND_GATE U2113 ( .I1(n1446), .I2(n1447), .O(n5436) );
  NAND_GATE U2114 ( .I1(n1436), .I2(donnee[5]), .O(n1447) );
  NAND_GATE U2115 ( .I1(\registres[10][5] ), .I2(n1437), .O(n1446) );
  NAND_GATE U2116 ( .I1(n1448), .I2(n1449), .O(n5437) );
  NAND_GATE U2117 ( .I1(n1436), .I2(donnee[6]), .O(n1449) );
  NAND_GATE U2118 ( .I1(\registres[10][6] ), .I2(n1437), .O(n1448) );
  NAND_GATE U2119 ( .I1(n1450), .I2(n1451), .O(n5438) );
  NAND_GATE U2120 ( .I1(n1436), .I2(donnee[7]), .O(n1451) );
  NAND_GATE U2121 ( .I1(\registres[10][7] ), .I2(n1437), .O(n1450) );
  NAND_GATE U2122 ( .I1(n1452), .I2(n1453), .O(n5439) );
  NAND_GATE U2123 ( .I1(n1436), .I2(donnee[8]), .O(n1453) );
  NAND_GATE U2124 ( .I1(\registres[10][8] ), .I2(n1437), .O(n1452) );
  NAND_GATE U2125 ( .I1(n1454), .I2(n1455), .O(n5440) );
  NAND_GATE U2126 ( .I1(n1436), .I2(donnee[9]), .O(n1455) );
  NAND_GATE U2127 ( .I1(\registres[10][9] ), .I2(n1437), .O(n1454) );
  NAND_GATE U2128 ( .I1(n1456), .I2(n1457), .O(n5441) );
  NAND_GATE U2129 ( .I1(n1436), .I2(donnee[10]), .O(n1457) );
  NAND_GATE U2130 ( .I1(\registres[10][10] ), .I2(n1437), .O(n1456) );
  NAND_GATE U2131 ( .I1(n1458), .I2(n1459), .O(n5442) );
  NAND_GATE U2132 ( .I1(n1436), .I2(donnee[11]), .O(n1459) );
  NAND_GATE U2133 ( .I1(\registres[10][11] ), .I2(n1437), .O(n1458) );
  NAND_GATE U2134 ( .I1(n1460), .I2(n1461), .O(n5443) );
  NAND_GATE U2135 ( .I1(n1436), .I2(donnee[12]), .O(n1461) );
  NAND_GATE U2136 ( .I1(\registres[10][12] ), .I2(n1437), .O(n1460) );
  NAND_GATE U2137 ( .I1(n1462), .I2(n1463), .O(n5444) );
  NAND_GATE U2138 ( .I1(n1436), .I2(donnee[13]), .O(n1463) );
  NAND_GATE U2139 ( .I1(\registres[10][13] ), .I2(n1437), .O(n1462) );
  NAND_GATE U2140 ( .I1(n1464), .I2(n1465), .O(n5445) );
  NAND_GATE U2141 ( .I1(n1436), .I2(donnee[14]), .O(n1465) );
  NAND_GATE U2142 ( .I1(\registres[10][14] ), .I2(n1437), .O(n1464) );
  NAND_GATE U2143 ( .I1(n1466), .I2(n1467), .O(n5446) );
  NAND_GATE U2144 ( .I1(n1436), .I2(donnee[15]), .O(n1467) );
  NAND_GATE U2145 ( .I1(\registres[10][15] ), .I2(n1437), .O(n1466) );
  NAND_GATE U2146 ( .I1(n1468), .I2(n1469), .O(n5447) );
  NAND_GATE U2147 ( .I1(n1436), .I2(donnee[16]), .O(n1469) );
  NAND_GATE U2148 ( .I1(\registres[10][16] ), .I2(n1437), .O(n1468) );
  NAND_GATE U2149 ( .I1(n1470), .I2(n1471), .O(n5448) );
  NAND_GATE U2150 ( .I1(n1436), .I2(donnee[17]), .O(n1471) );
  NAND_GATE U2151 ( .I1(\registres[10][17] ), .I2(n1437), .O(n1470) );
  NAND_GATE U2152 ( .I1(n1472), .I2(n1473), .O(n5449) );
  NAND_GATE U2153 ( .I1(n1436), .I2(donnee[18]), .O(n1473) );
  NAND_GATE U2154 ( .I1(\registres[10][18] ), .I2(n1437), .O(n1472) );
  NAND_GATE U2155 ( .I1(n1474), .I2(n1475), .O(n5450) );
  NAND_GATE U2156 ( .I1(n1436), .I2(donnee[19]), .O(n1475) );
  NAND_GATE U2157 ( .I1(\registres[10][19] ), .I2(n1437), .O(n1474) );
  NAND_GATE U2158 ( .I1(n1476), .I2(n1477), .O(n5451) );
  NAND_GATE U2159 ( .I1(n1436), .I2(donnee[20]), .O(n1477) );
  NAND_GATE U2160 ( .I1(\registres[10][20] ), .I2(n1437), .O(n1476) );
  NAND_GATE U2161 ( .I1(n1478), .I2(n1479), .O(n5452) );
  NAND_GATE U2162 ( .I1(n1436), .I2(donnee[21]), .O(n1479) );
  NAND_GATE U2163 ( .I1(\registres[10][21] ), .I2(n1437), .O(n1478) );
  NAND_GATE U2164 ( .I1(n1480), .I2(n1481), .O(n5453) );
  NAND_GATE U2165 ( .I1(n1436), .I2(donnee[22]), .O(n1481) );
  NAND_GATE U2166 ( .I1(\registres[10][22] ), .I2(n1437), .O(n1480) );
  NAND_GATE U2167 ( .I1(n1482), .I2(n1483), .O(n5454) );
  NAND_GATE U2168 ( .I1(n1436), .I2(donnee[23]), .O(n1483) );
  NAND_GATE U2169 ( .I1(\registres[10][23] ), .I2(n1437), .O(n1482) );
  NAND_GATE U2170 ( .I1(n1484), .I2(n1485), .O(n5455) );
  NAND_GATE U2171 ( .I1(n1436), .I2(donnee[24]), .O(n1485) );
  NAND_GATE U2172 ( .I1(\registres[10][24] ), .I2(n1437), .O(n1484) );
  NAND_GATE U2173 ( .I1(n1486), .I2(n1487), .O(n5456) );
  NAND_GATE U2174 ( .I1(n1436), .I2(donnee[25]), .O(n1487) );
  NAND_GATE U2175 ( .I1(\registres[10][25] ), .I2(n1437), .O(n1486) );
  NAND_GATE U2176 ( .I1(n1488), .I2(n1489), .O(n5457) );
  NAND_GATE U2177 ( .I1(n1436), .I2(donnee[26]), .O(n1489) );
  NAND_GATE U2178 ( .I1(\registres[10][26] ), .I2(n1437), .O(n1488) );
  NAND_GATE U2179 ( .I1(n1490), .I2(n1491), .O(n5458) );
  NAND_GATE U2180 ( .I1(n1436), .I2(donnee[27]), .O(n1491) );
  NAND_GATE U2181 ( .I1(\registres[10][27] ), .I2(n1437), .O(n1490) );
  NAND_GATE U2182 ( .I1(n1492), .I2(n1493), .O(n5459) );
  NAND_GATE U2183 ( .I1(n1436), .I2(donnee[28]), .O(n1493) );
  NAND_GATE U2184 ( .I1(\registres[10][28] ), .I2(n1437), .O(n1492) );
  NAND_GATE U2185 ( .I1(n1494), .I2(n1495), .O(n5460) );
  NAND_GATE U2186 ( .I1(n1436), .I2(donnee[29]), .O(n1495) );
  NAND_GATE U2187 ( .I1(\registres[10][29] ), .I2(n1437), .O(n1494) );
  NAND_GATE U2188 ( .I1(n1496), .I2(n1497), .O(n5461) );
  NAND_GATE U2189 ( .I1(n1436), .I2(donnee[30]), .O(n1497) );
  NAND_GATE U2190 ( .I1(\registres[10][30] ), .I2(n1437), .O(n1496) );
  NAND_GATE U2191 ( .I1(n1498), .I2(n1499), .O(n5462) );
  NAND_GATE U2192 ( .I1(n1436), .I2(donnee[31]), .O(n1499) );
  AND_GATE U2193 ( .I1(n1500), .I2(n1), .O(n1436) );
  NAND_GATE U2194 ( .I1(\registres[10][31] ), .I2(n1437), .O(n1498) );
  NOR_GATE U2195 ( .I1(n1500), .I2(reset), .O(n1437) );
  AND3_GATE U2196 ( .I1(n424), .I2(cmd_ecr), .I3(n1165), .O(n1500) );
  NAND_GATE U2197 ( .I1(n1501), .I2(n1502), .O(n5463) );
  NAND_GATE U2198 ( .I1(n1503), .I2(donnee[0]), .O(n1502) );
  NAND_GATE U2199 ( .I1(\registres[9][0] ), .I2(n1504), .O(n1501) );
  NAND_GATE U2200 ( .I1(n1505), .I2(n1506), .O(n5464) );
  NAND_GATE U2201 ( .I1(n1503), .I2(donnee[1]), .O(n1506) );
  NAND_GATE U2202 ( .I1(\registres[9][1] ), .I2(n1504), .O(n1505) );
  NAND_GATE U2203 ( .I1(n1507), .I2(n1508), .O(n5465) );
  NAND_GATE U2204 ( .I1(n1503), .I2(donnee[2]), .O(n1508) );
  NAND_GATE U2205 ( .I1(\registres[9][2] ), .I2(n1504), .O(n1507) );
  NAND_GATE U2206 ( .I1(n1509), .I2(n1510), .O(n5466) );
  NAND_GATE U2207 ( .I1(n1503), .I2(donnee[3]), .O(n1510) );
  NAND_GATE U2208 ( .I1(\registres[9][3] ), .I2(n1504), .O(n1509) );
  NAND_GATE U2209 ( .I1(n1511), .I2(n1512), .O(n5467) );
  NAND_GATE U2210 ( .I1(n1503), .I2(donnee[4]), .O(n1512) );
  NAND_GATE U2211 ( .I1(\registres[9][4] ), .I2(n1504), .O(n1511) );
  NAND_GATE U2212 ( .I1(n1513), .I2(n1514), .O(n5468) );
  NAND_GATE U2213 ( .I1(n1503), .I2(donnee[5]), .O(n1514) );
  NAND_GATE U2214 ( .I1(\registres[9][5] ), .I2(n1504), .O(n1513) );
  NAND_GATE U2215 ( .I1(n1515), .I2(n1516), .O(n5469) );
  NAND_GATE U2216 ( .I1(n1503), .I2(donnee[6]), .O(n1516) );
  NAND_GATE U2217 ( .I1(\registres[9][6] ), .I2(n1504), .O(n1515) );
  NAND_GATE U2218 ( .I1(n1517), .I2(n1518), .O(n5470) );
  NAND_GATE U2219 ( .I1(n1503), .I2(donnee[7]), .O(n1518) );
  NAND_GATE U2220 ( .I1(\registres[9][7] ), .I2(n1504), .O(n1517) );
  NAND_GATE U2221 ( .I1(n1519), .I2(n1520), .O(n5471) );
  NAND_GATE U2222 ( .I1(n1503), .I2(donnee[8]), .O(n1520) );
  NAND_GATE U2223 ( .I1(\registres[9][8] ), .I2(n1504), .O(n1519) );
  NAND_GATE U2224 ( .I1(n1521), .I2(n1522), .O(n5472) );
  NAND_GATE U2225 ( .I1(n1503), .I2(donnee[9]), .O(n1522) );
  NAND_GATE U2226 ( .I1(\registres[9][9] ), .I2(n1504), .O(n1521) );
  NAND_GATE U2227 ( .I1(n1523), .I2(n1524), .O(n5473) );
  NAND_GATE U2228 ( .I1(n1503), .I2(donnee[10]), .O(n1524) );
  NAND_GATE U2229 ( .I1(\registres[9][10] ), .I2(n1504), .O(n1523) );
  NAND_GATE U2230 ( .I1(n1525), .I2(n1526), .O(n5474) );
  NAND_GATE U2231 ( .I1(n1503), .I2(donnee[11]), .O(n1526) );
  NAND_GATE U2232 ( .I1(\registres[9][11] ), .I2(n1504), .O(n1525) );
  NAND_GATE U2233 ( .I1(n1527), .I2(n1528), .O(n5475) );
  NAND_GATE U2234 ( .I1(n1503), .I2(donnee[12]), .O(n1528) );
  NAND_GATE U2235 ( .I1(\registres[9][12] ), .I2(n1504), .O(n1527) );
  NAND_GATE U2236 ( .I1(n1529), .I2(n1530), .O(n5476) );
  NAND_GATE U2237 ( .I1(n1503), .I2(donnee[13]), .O(n1530) );
  NAND_GATE U2238 ( .I1(\registres[9][13] ), .I2(n1504), .O(n1529) );
  NAND_GATE U2239 ( .I1(n1531), .I2(n1532), .O(n5477) );
  NAND_GATE U2240 ( .I1(n1503), .I2(donnee[14]), .O(n1532) );
  NAND_GATE U2241 ( .I1(\registres[9][14] ), .I2(n1504), .O(n1531) );
  NAND_GATE U2242 ( .I1(n1533), .I2(n1534), .O(n5478) );
  NAND_GATE U2243 ( .I1(n1503), .I2(donnee[15]), .O(n1534) );
  NAND_GATE U2244 ( .I1(\registres[9][15] ), .I2(n1504), .O(n1533) );
  NAND_GATE U2245 ( .I1(n1535), .I2(n1536), .O(n5479) );
  NAND_GATE U2246 ( .I1(n1503), .I2(donnee[16]), .O(n1536) );
  NAND_GATE U2247 ( .I1(\registres[9][16] ), .I2(n1504), .O(n1535) );
  NAND_GATE U2248 ( .I1(n1537), .I2(n1538), .O(n5480) );
  NAND_GATE U2249 ( .I1(n1503), .I2(donnee[17]), .O(n1538) );
  NAND_GATE U2250 ( .I1(\registres[9][17] ), .I2(n1504), .O(n1537) );
  NAND_GATE U2251 ( .I1(n1539), .I2(n1540), .O(n5481) );
  NAND_GATE U2252 ( .I1(n1503), .I2(donnee[18]), .O(n1540) );
  NAND_GATE U2253 ( .I1(\registres[9][18] ), .I2(n1504), .O(n1539) );
  NAND_GATE U2254 ( .I1(n1541), .I2(n1542), .O(n5482) );
  NAND_GATE U2255 ( .I1(n1503), .I2(donnee[19]), .O(n1542) );
  NAND_GATE U2256 ( .I1(\registres[9][19] ), .I2(n1504), .O(n1541) );
  NAND_GATE U2257 ( .I1(n1543), .I2(n1544), .O(n5483) );
  NAND_GATE U2258 ( .I1(n1503), .I2(donnee[20]), .O(n1544) );
  NAND_GATE U2259 ( .I1(\registres[9][20] ), .I2(n1504), .O(n1543) );
  NAND_GATE U2260 ( .I1(n1545), .I2(n1546), .O(n5484) );
  NAND_GATE U2261 ( .I1(n1503), .I2(donnee[21]), .O(n1546) );
  NAND_GATE U2262 ( .I1(\registres[9][21] ), .I2(n1504), .O(n1545) );
  NAND_GATE U2263 ( .I1(n1547), .I2(n1548), .O(n5485) );
  NAND_GATE U2264 ( .I1(n1503), .I2(donnee[22]), .O(n1548) );
  NAND_GATE U2265 ( .I1(\registres[9][22] ), .I2(n1504), .O(n1547) );
  NAND_GATE U2266 ( .I1(n1549), .I2(n1550), .O(n5486) );
  NAND_GATE U2267 ( .I1(n1503), .I2(donnee[23]), .O(n1550) );
  NAND_GATE U2268 ( .I1(\registres[9][23] ), .I2(n1504), .O(n1549) );
  NAND_GATE U2269 ( .I1(n1551), .I2(n1552), .O(n5487) );
  NAND_GATE U2270 ( .I1(n1503), .I2(donnee[24]), .O(n1552) );
  NAND_GATE U2271 ( .I1(\registres[9][24] ), .I2(n1504), .O(n1551) );
  NAND_GATE U2272 ( .I1(n1553), .I2(n1554), .O(n5488) );
  NAND_GATE U2273 ( .I1(n1503), .I2(donnee[25]), .O(n1554) );
  NAND_GATE U2274 ( .I1(\registres[9][25] ), .I2(n1504), .O(n1553) );
  NAND_GATE U2275 ( .I1(n1555), .I2(n1556), .O(n5489) );
  NAND_GATE U2276 ( .I1(n1503), .I2(donnee[26]), .O(n1556) );
  NAND_GATE U2277 ( .I1(\registres[9][26] ), .I2(n1504), .O(n1555) );
  NAND_GATE U2278 ( .I1(n1557), .I2(n1558), .O(n5490) );
  NAND_GATE U2279 ( .I1(n1503), .I2(donnee[27]), .O(n1558) );
  NAND_GATE U2280 ( .I1(\registres[9][27] ), .I2(n1504), .O(n1557) );
  NAND_GATE U2281 ( .I1(n1559), .I2(n1560), .O(n5491) );
  NAND_GATE U2282 ( .I1(n1503), .I2(donnee[28]), .O(n1560) );
  NAND_GATE U2283 ( .I1(\registres[9][28] ), .I2(n1504), .O(n1559) );
  NAND_GATE U2284 ( .I1(n1561), .I2(n1562), .O(n5492) );
  NAND_GATE U2285 ( .I1(n1503), .I2(donnee[29]), .O(n1562) );
  NAND_GATE U2286 ( .I1(\registres[9][29] ), .I2(n1504), .O(n1561) );
  NAND_GATE U2287 ( .I1(n1563), .I2(n1564), .O(n5493) );
  NAND_GATE U2288 ( .I1(n1503), .I2(donnee[30]), .O(n1564) );
  NAND_GATE U2289 ( .I1(\registres[9][30] ), .I2(n1504), .O(n1563) );
  NAND_GATE U2290 ( .I1(n1565), .I2(n1566), .O(n5494) );
  NAND_GATE U2291 ( .I1(n1503), .I2(donnee[31]), .O(n1566) );
  AND_GATE U2292 ( .I1(n1567), .I2(n1), .O(n1503) );
  NAND_GATE U2293 ( .I1(\registres[9][31] ), .I2(n1504), .O(n1565) );
  NOR_GATE U2294 ( .I1(n1567), .I2(reset), .O(n1504) );
  AND3_GATE U2295 ( .I1(n492), .I2(cmd_ecr), .I3(n1165), .O(n1567) );
  NAND_GATE U2296 ( .I1(n1568), .I2(n1569), .O(n5495) );
  NAND_GATE U2297 ( .I1(n1570), .I2(donnee[0]), .O(n1569) );
  NAND_GATE U2298 ( .I1(\registres[8][0] ), .I2(n1571), .O(n1568) );
  NAND_GATE U2299 ( .I1(n1572), .I2(n1573), .O(n5496) );
  NAND_GATE U2300 ( .I1(n1570), .I2(donnee[1]), .O(n1573) );
  NAND_GATE U2301 ( .I1(\registres[8][1] ), .I2(n1571), .O(n1572) );
  NAND_GATE U2302 ( .I1(n1574), .I2(n1575), .O(n5497) );
  NAND_GATE U2303 ( .I1(n1570), .I2(donnee[2]), .O(n1575) );
  NAND_GATE U2304 ( .I1(\registres[8][2] ), .I2(n1571), .O(n1574) );
  NAND_GATE U2305 ( .I1(n1576), .I2(n1577), .O(n5498) );
  NAND_GATE U2306 ( .I1(n1570), .I2(donnee[3]), .O(n1577) );
  NAND_GATE U2307 ( .I1(\registres[8][3] ), .I2(n1571), .O(n1576) );
  NAND_GATE U2308 ( .I1(n1578), .I2(n1579), .O(n5499) );
  NAND_GATE U2309 ( .I1(n1570), .I2(donnee[4]), .O(n1579) );
  NAND_GATE U2310 ( .I1(\registres[8][4] ), .I2(n1571), .O(n1578) );
  NAND_GATE U2311 ( .I1(n1580), .I2(n1581), .O(n5500) );
  NAND_GATE U2312 ( .I1(n1570), .I2(donnee[5]), .O(n1581) );
  NAND_GATE U2313 ( .I1(\registres[8][5] ), .I2(n1571), .O(n1580) );
  NAND_GATE U2314 ( .I1(n1582), .I2(n1583), .O(n5501) );
  NAND_GATE U2315 ( .I1(n1570), .I2(donnee[6]), .O(n1583) );
  NAND_GATE U2316 ( .I1(\registres[8][6] ), .I2(n1571), .O(n1582) );
  NAND_GATE U2317 ( .I1(n1584), .I2(n1585), .O(n5502) );
  NAND_GATE U2318 ( .I1(n1570), .I2(donnee[7]), .O(n1585) );
  NAND_GATE U2319 ( .I1(\registres[8][7] ), .I2(n1571), .O(n1584) );
  NAND_GATE U2320 ( .I1(n1586), .I2(n1587), .O(n5503) );
  NAND_GATE U2321 ( .I1(n1570), .I2(donnee[8]), .O(n1587) );
  NAND_GATE U2322 ( .I1(\registres[8][8] ), .I2(n1571), .O(n1586) );
  NAND_GATE U2323 ( .I1(n1588), .I2(n1589), .O(n5504) );
  NAND_GATE U2324 ( .I1(n1570), .I2(donnee[9]), .O(n1589) );
  NAND_GATE U2325 ( .I1(\registres[8][9] ), .I2(n1571), .O(n1588) );
  NAND_GATE U2326 ( .I1(n1590), .I2(n1591), .O(n5505) );
  NAND_GATE U2327 ( .I1(n1570), .I2(donnee[10]), .O(n1591) );
  NAND_GATE U2328 ( .I1(\registres[8][10] ), .I2(n1571), .O(n1590) );
  NAND_GATE U2329 ( .I1(n1592), .I2(n1593), .O(n5506) );
  NAND_GATE U2330 ( .I1(n1570), .I2(donnee[11]), .O(n1593) );
  NAND_GATE U2331 ( .I1(\registres[8][11] ), .I2(n1571), .O(n1592) );
  NAND_GATE U2332 ( .I1(n1594), .I2(n1595), .O(n5507) );
  NAND_GATE U2333 ( .I1(n1570), .I2(donnee[12]), .O(n1595) );
  NAND_GATE U2334 ( .I1(\registres[8][12] ), .I2(n1571), .O(n1594) );
  NAND_GATE U2335 ( .I1(n1596), .I2(n1597), .O(n5508) );
  NAND_GATE U2336 ( .I1(n1570), .I2(donnee[13]), .O(n1597) );
  NAND_GATE U2337 ( .I1(\registres[8][13] ), .I2(n1571), .O(n1596) );
  NAND_GATE U2338 ( .I1(n1598), .I2(n1599), .O(n5509) );
  NAND_GATE U2339 ( .I1(n1570), .I2(donnee[14]), .O(n1599) );
  NAND_GATE U2340 ( .I1(\registres[8][14] ), .I2(n1571), .O(n1598) );
  NAND_GATE U2341 ( .I1(n1600), .I2(n1601), .O(n5510) );
  NAND_GATE U2342 ( .I1(n1570), .I2(donnee[15]), .O(n1601) );
  NAND_GATE U2343 ( .I1(\registres[8][15] ), .I2(n1571), .O(n1600) );
  NAND_GATE U2344 ( .I1(n1602), .I2(n1603), .O(n5511) );
  NAND_GATE U2345 ( .I1(n1570), .I2(donnee[16]), .O(n1603) );
  NAND_GATE U2346 ( .I1(\registres[8][16] ), .I2(n1571), .O(n1602) );
  NAND_GATE U2347 ( .I1(n1604), .I2(n1605), .O(n5512) );
  NAND_GATE U2348 ( .I1(n1570), .I2(donnee[17]), .O(n1605) );
  NAND_GATE U2349 ( .I1(\registres[8][17] ), .I2(n1571), .O(n1604) );
  NAND_GATE U2350 ( .I1(n1606), .I2(n1607), .O(n5513) );
  NAND_GATE U2351 ( .I1(n1570), .I2(donnee[18]), .O(n1607) );
  NAND_GATE U2352 ( .I1(\registres[8][18] ), .I2(n1571), .O(n1606) );
  NAND_GATE U2353 ( .I1(n1608), .I2(n1609), .O(n5514) );
  NAND_GATE U2354 ( .I1(n1570), .I2(donnee[19]), .O(n1609) );
  NAND_GATE U2355 ( .I1(\registres[8][19] ), .I2(n1571), .O(n1608) );
  NAND_GATE U2356 ( .I1(n1610), .I2(n1611), .O(n5515) );
  NAND_GATE U2357 ( .I1(n1570), .I2(donnee[20]), .O(n1611) );
  NAND_GATE U2358 ( .I1(\registres[8][20] ), .I2(n1571), .O(n1610) );
  NAND_GATE U2359 ( .I1(n1612), .I2(n1613), .O(n5516) );
  NAND_GATE U2360 ( .I1(n1570), .I2(donnee[21]), .O(n1613) );
  NAND_GATE U2361 ( .I1(\registres[8][21] ), .I2(n1571), .O(n1612) );
  NAND_GATE U2362 ( .I1(n1614), .I2(n1615), .O(n5517) );
  NAND_GATE U2363 ( .I1(n1570), .I2(donnee[22]), .O(n1615) );
  NAND_GATE U2364 ( .I1(\registres[8][22] ), .I2(n1571), .O(n1614) );
  NAND_GATE U2365 ( .I1(n1616), .I2(n1617), .O(n5518) );
  NAND_GATE U2366 ( .I1(n1570), .I2(donnee[23]), .O(n1617) );
  NAND_GATE U2367 ( .I1(\registres[8][23] ), .I2(n1571), .O(n1616) );
  NAND_GATE U2368 ( .I1(n1618), .I2(n1619), .O(n5519) );
  NAND_GATE U2369 ( .I1(n1570), .I2(donnee[24]), .O(n1619) );
  NAND_GATE U2370 ( .I1(\registres[8][24] ), .I2(n1571), .O(n1618) );
  NAND_GATE U2371 ( .I1(n1620), .I2(n1621), .O(n5520) );
  NAND_GATE U2372 ( .I1(n1570), .I2(donnee[25]), .O(n1621) );
  NAND_GATE U2373 ( .I1(\registres[8][25] ), .I2(n1571), .O(n1620) );
  NAND_GATE U2374 ( .I1(n1622), .I2(n1623), .O(n5521) );
  NAND_GATE U2375 ( .I1(n1570), .I2(donnee[26]), .O(n1623) );
  NAND_GATE U2376 ( .I1(\registres[8][26] ), .I2(n1571), .O(n1622) );
  NAND_GATE U2377 ( .I1(n1624), .I2(n1625), .O(n5522) );
  NAND_GATE U2378 ( .I1(n1570), .I2(donnee[27]), .O(n1625) );
  NAND_GATE U2379 ( .I1(\registres[8][27] ), .I2(n1571), .O(n1624) );
  NAND_GATE U2380 ( .I1(n1626), .I2(n1627), .O(n5523) );
  NAND_GATE U2381 ( .I1(n1570), .I2(donnee[28]), .O(n1627) );
  NAND_GATE U2382 ( .I1(\registres[8][28] ), .I2(n1571), .O(n1626) );
  NAND_GATE U2383 ( .I1(n1628), .I2(n1629), .O(n5524) );
  NAND_GATE U2384 ( .I1(n1570), .I2(donnee[29]), .O(n1629) );
  NAND_GATE U2385 ( .I1(\registres[8][29] ), .I2(n1571), .O(n1628) );
  NAND_GATE U2386 ( .I1(n1630), .I2(n1631), .O(n5525) );
  NAND_GATE U2387 ( .I1(n1570), .I2(donnee[30]), .O(n1631) );
  NAND_GATE U2388 ( .I1(\registres[8][30] ), .I2(n1571), .O(n1630) );
  NAND_GATE U2389 ( .I1(n1632), .I2(n1633), .O(n5526) );
  NAND_GATE U2390 ( .I1(n1570), .I2(donnee[31]), .O(n1633) );
  AND_GATE U2391 ( .I1(n1634), .I2(n1), .O(n1570) );
  NAND_GATE U2392 ( .I1(\registres[8][31] ), .I2(n1571), .O(n1632) );
  NOR_GATE U2393 ( .I1(n1634), .I2(reset), .O(n1571) );
  AND3_GATE U2394 ( .I1(n560), .I2(cmd_ecr), .I3(n1165), .O(n1634) );
  AND_GATE U2395 ( .I1(reg_dest[3]), .I2(n2), .O(n1165) );
  NOR3_GATE U2396 ( .I1(reg_dest[2]), .I2(reg_dest[1]), .I3(reg_dest[0]), .O(
        n560) );
  NAND_GATE U2397 ( .I1(n1635), .I2(n1636), .O(n5527) );
  NAND_GATE U2398 ( .I1(n1637), .I2(donnee[0]), .O(n1636) );
  NAND_GATE U2399 ( .I1(\registres[7][0] ), .I2(n1638), .O(n1635) );
  NAND_GATE U2400 ( .I1(n1639), .I2(n1640), .O(n5528) );
  NAND_GATE U2401 ( .I1(n1637), .I2(donnee[1]), .O(n1640) );
  NAND_GATE U2402 ( .I1(\registres[7][1] ), .I2(n1638), .O(n1639) );
  NAND_GATE U2403 ( .I1(n1641), .I2(n1642), .O(n5529) );
  NAND_GATE U2404 ( .I1(n1637), .I2(donnee[2]), .O(n1642) );
  NAND_GATE U2405 ( .I1(\registres[7][2] ), .I2(n1638), .O(n1641) );
  NAND_GATE U2406 ( .I1(n1643), .I2(n1644), .O(n5530) );
  NAND_GATE U2407 ( .I1(n1637), .I2(donnee[3]), .O(n1644) );
  NAND_GATE U2408 ( .I1(\registres[7][3] ), .I2(n1638), .O(n1643) );
  NAND_GATE U2409 ( .I1(n1645), .I2(n1646), .O(n5531) );
  NAND_GATE U2410 ( .I1(n1637), .I2(donnee[4]), .O(n1646) );
  NAND_GATE U2411 ( .I1(\registres[7][4] ), .I2(n1638), .O(n1645) );
  NAND_GATE U2412 ( .I1(n1647), .I2(n1648), .O(n5532) );
  NAND_GATE U2413 ( .I1(n1637), .I2(donnee[5]), .O(n1648) );
  NAND_GATE U2414 ( .I1(\registres[7][5] ), .I2(n1638), .O(n1647) );
  NAND_GATE U2415 ( .I1(n1649), .I2(n1650), .O(n5533) );
  NAND_GATE U2416 ( .I1(n1637), .I2(donnee[6]), .O(n1650) );
  NAND_GATE U2417 ( .I1(\registres[7][6] ), .I2(n1638), .O(n1649) );
  NAND_GATE U2418 ( .I1(n1651), .I2(n1652), .O(n5534) );
  NAND_GATE U2419 ( .I1(n1637), .I2(donnee[7]), .O(n1652) );
  NAND_GATE U2420 ( .I1(\registres[7][7] ), .I2(n1638), .O(n1651) );
  NAND_GATE U2421 ( .I1(n1653), .I2(n1654), .O(n5535) );
  NAND_GATE U2422 ( .I1(n1637), .I2(donnee[8]), .O(n1654) );
  NAND_GATE U2423 ( .I1(\registres[7][8] ), .I2(n1638), .O(n1653) );
  NAND_GATE U2424 ( .I1(n1655), .I2(n1656), .O(n5536) );
  NAND_GATE U2425 ( .I1(n1637), .I2(donnee[9]), .O(n1656) );
  NAND_GATE U2426 ( .I1(\registres[7][9] ), .I2(n1638), .O(n1655) );
  NAND_GATE U2427 ( .I1(n1657), .I2(n1658), .O(n5537) );
  NAND_GATE U2428 ( .I1(n1637), .I2(donnee[10]), .O(n1658) );
  NAND_GATE U2429 ( .I1(\registres[7][10] ), .I2(n1638), .O(n1657) );
  NAND_GATE U2430 ( .I1(n1659), .I2(n1660), .O(n5538) );
  NAND_GATE U2431 ( .I1(n1637), .I2(donnee[11]), .O(n1660) );
  NAND_GATE U2432 ( .I1(\registres[7][11] ), .I2(n1638), .O(n1659) );
  NAND_GATE U2433 ( .I1(n1661), .I2(n1662), .O(n5539) );
  NAND_GATE U2434 ( .I1(n1637), .I2(donnee[12]), .O(n1662) );
  NAND_GATE U2435 ( .I1(\registres[7][12] ), .I2(n1638), .O(n1661) );
  NAND_GATE U2436 ( .I1(n1663), .I2(n1664), .O(n5540) );
  NAND_GATE U2437 ( .I1(n1637), .I2(donnee[13]), .O(n1664) );
  NAND_GATE U2438 ( .I1(\registres[7][13] ), .I2(n1638), .O(n1663) );
  NAND_GATE U2439 ( .I1(n1665), .I2(n1666), .O(n5541) );
  NAND_GATE U2440 ( .I1(n1637), .I2(donnee[14]), .O(n1666) );
  NAND_GATE U2441 ( .I1(\registres[7][14] ), .I2(n1638), .O(n1665) );
  NAND_GATE U2442 ( .I1(n1667), .I2(n1668), .O(n5542) );
  NAND_GATE U2443 ( .I1(n1637), .I2(donnee[15]), .O(n1668) );
  NAND_GATE U2444 ( .I1(\registres[7][15] ), .I2(n1638), .O(n1667) );
  NAND_GATE U2445 ( .I1(n1669), .I2(n1670), .O(n5543) );
  NAND_GATE U2446 ( .I1(n1637), .I2(donnee[16]), .O(n1670) );
  NAND_GATE U2447 ( .I1(\registres[7][16] ), .I2(n1638), .O(n1669) );
  NAND_GATE U2448 ( .I1(n1671), .I2(n1672), .O(n5544) );
  NAND_GATE U2449 ( .I1(n1637), .I2(donnee[17]), .O(n1672) );
  NAND_GATE U2450 ( .I1(\registres[7][17] ), .I2(n1638), .O(n1671) );
  NAND_GATE U2451 ( .I1(n1673), .I2(n1674), .O(n5545) );
  NAND_GATE U2452 ( .I1(n1637), .I2(donnee[18]), .O(n1674) );
  NAND_GATE U2453 ( .I1(\registres[7][18] ), .I2(n1638), .O(n1673) );
  NAND_GATE U2454 ( .I1(n1675), .I2(n1676), .O(n5546) );
  NAND_GATE U2455 ( .I1(n1637), .I2(donnee[19]), .O(n1676) );
  NAND_GATE U2456 ( .I1(\registres[7][19] ), .I2(n1638), .O(n1675) );
  NAND_GATE U2457 ( .I1(n1677), .I2(n1678), .O(n5547) );
  NAND_GATE U2458 ( .I1(n1637), .I2(donnee[20]), .O(n1678) );
  NAND_GATE U2459 ( .I1(\registres[7][20] ), .I2(n1638), .O(n1677) );
  NAND_GATE U2460 ( .I1(n1679), .I2(n1680), .O(n5548) );
  NAND_GATE U2461 ( .I1(n1637), .I2(donnee[21]), .O(n1680) );
  NAND_GATE U2462 ( .I1(\registres[7][21] ), .I2(n1638), .O(n1679) );
  NAND_GATE U2463 ( .I1(n1681), .I2(n1682), .O(n5549) );
  NAND_GATE U2464 ( .I1(n1637), .I2(donnee[22]), .O(n1682) );
  NAND_GATE U2465 ( .I1(\registres[7][22] ), .I2(n1638), .O(n1681) );
  NAND_GATE U2466 ( .I1(n1683), .I2(n1684), .O(n5550) );
  NAND_GATE U2467 ( .I1(n1637), .I2(donnee[23]), .O(n1684) );
  NAND_GATE U2468 ( .I1(\registres[7][23] ), .I2(n1638), .O(n1683) );
  NAND_GATE U2469 ( .I1(n1685), .I2(n1686), .O(n5551) );
  NAND_GATE U2470 ( .I1(n1637), .I2(donnee[24]), .O(n1686) );
  NAND_GATE U2471 ( .I1(\registres[7][24] ), .I2(n1638), .O(n1685) );
  NAND_GATE U2472 ( .I1(n1687), .I2(n1688), .O(n5552) );
  NAND_GATE U2473 ( .I1(n1637), .I2(donnee[25]), .O(n1688) );
  NAND_GATE U2474 ( .I1(\registres[7][25] ), .I2(n1638), .O(n1687) );
  NAND_GATE U2475 ( .I1(n1689), .I2(n1690), .O(n5553) );
  NAND_GATE U2476 ( .I1(n1637), .I2(donnee[26]), .O(n1690) );
  NAND_GATE U2477 ( .I1(\registres[7][26] ), .I2(n1638), .O(n1689) );
  NAND_GATE U2478 ( .I1(n1691), .I2(n1692), .O(n5554) );
  NAND_GATE U2479 ( .I1(n1637), .I2(donnee[27]), .O(n1692) );
  NAND_GATE U2480 ( .I1(\registres[7][27] ), .I2(n1638), .O(n1691) );
  NAND_GATE U2481 ( .I1(n1693), .I2(n1694), .O(n5555) );
  NAND_GATE U2482 ( .I1(n1637), .I2(donnee[28]), .O(n1694) );
  NAND_GATE U2483 ( .I1(\registres[7][28] ), .I2(n1638), .O(n1693) );
  NAND_GATE U2484 ( .I1(n1695), .I2(n1696), .O(n5556) );
  NAND_GATE U2485 ( .I1(n1637), .I2(donnee[29]), .O(n1696) );
  NAND_GATE U2486 ( .I1(\registres[7][29] ), .I2(n1638), .O(n1695) );
  NAND_GATE U2487 ( .I1(n1697), .I2(n1698), .O(n5557) );
  NAND_GATE U2488 ( .I1(n1637), .I2(donnee[30]), .O(n1698) );
  NAND_GATE U2489 ( .I1(\registres[7][30] ), .I2(n1638), .O(n1697) );
  NAND_GATE U2490 ( .I1(n1699), .I2(n1700), .O(n5558) );
  NAND_GATE U2491 ( .I1(n1637), .I2(donnee[31]), .O(n1700) );
  AND_GATE U2492 ( .I1(n1701), .I2(n1), .O(n1637) );
  NAND_GATE U2493 ( .I1(\registres[7][31] ), .I2(n1638), .O(n1699) );
  NOR_GATE U2494 ( .I1(n1701), .I2(reset), .O(n1638) );
  AND3_GATE U2495 ( .I1(n84), .I2(cmd_ecr), .I3(n1702), .O(n1701) );
  AND3_GATE U2496 ( .I1(reg_dest[1]), .I2(reg_dest[0]), .I3(reg_dest[2]), .O(
        n84) );
  NAND_GATE U2497 ( .I1(n1703), .I2(n1704), .O(n5559) );
  NAND_GATE U2498 ( .I1(n1705), .I2(donnee[0]), .O(n1704) );
  NAND_GATE U2499 ( .I1(\registres[6][0] ), .I2(n1706), .O(n1703) );
  NAND_GATE U2500 ( .I1(n1707), .I2(n1708), .O(n5560) );
  NAND_GATE U2501 ( .I1(n1705), .I2(donnee[1]), .O(n1708) );
  NAND_GATE U2502 ( .I1(\registres[6][1] ), .I2(n1706), .O(n1707) );
  NAND_GATE U2503 ( .I1(n1709), .I2(n1710), .O(n5561) );
  NAND_GATE U2504 ( .I1(n1705), .I2(donnee[2]), .O(n1710) );
  NAND_GATE U2505 ( .I1(\registres[6][2] ), .I2(n1706), .O(n1709) );
  NAND_GATE U2506 ( .I1(n1711), .I2(n1712), .O(n5562) );
  NAND_GATE U2507 ( .I1(n1705), .I2(donnee[3]), .O(n1712) );
  NAND_GATE U2508 ( .I1(\registres[6][3] ), .I2(n1706), .O(n1711) );
  NAND_GATE U2509 ( .I1(n1713), .I2(n1714), .O(n5563) );
  NAND_GATE U2510 ( .I1(n1705), .I2(donnee[4]), .O(n1714) );
  NAND_GATE U2511 ( .I1(\registres[6][4] ), .I2(n1706), .O(n1713) );
  NAND_GATE U2512 ( .I1(n1715), .I2(n1716), .O(n5564) );
  NAND_GATE U2513 ( .I1(n1705), .I2(donnee[5]), .O(n1716) );
  NAND_GATE U2514 ( .I1(\registres[6][5] ), .I2(n1706), .O(n1715) );
  NAND_GATE U2515 ( .I1(n1717), .I2(n1718), .O(n5565) );
  NAND_GATE U2516 ( .I1(n1705), .I2(donnee[6]), .O(n1718) );
  NAND_GATE U2517 ( .I1(\registres[6][6] ), .I2(n1706), .O(n1717) );
  NAND_GATE U2518 ( .I1(n1719), .I2(n1720), .O(n5566) );
  NAND_GATE U2519 ( .I1(n1705), .I2(donnee[7]), .O(n1720) );
  NAND_GATE U2520 ( .I1(\registres[6][7] ), .I2(n1706), .O(n1719) );
  NAND_GATE U2521 ( .I1(n1721), .I2(n1722), .O(n5567) );
  NAND_GATE U2522 ( .I1(n1705), .I2(donnee[8]), .O(n1722) );
  NAND_GATE U2523 ( .I1(\registres[6][8] ), .I2(n1706), .O(n1721) );
  NAND_GATE U2524 ( .I1(n1723), .I2(n1724), .O(n5568) );
  NAND_GATE U2525 ( .I1(n1705), .I2(donnee[9]), .O(n1724) );
  NAND_GATE U2526 ( .I1(\registres[6][9] ), .I2(n1706), .O(n1723) );
  NAND_GATE U2527 ( .I1(n1725), .I2(n1726), .O(n5569) );
  NAND_GATE U2528 ( .I1(n1705), .I2(donnee[10]), .O(n1726) );
  NAND_GATE U2529 ( .I1(\registres[6][10] ), .I2(n1706), .O(n1725) );
  NAND_GATE U2530 ( .I1(n1727), .I2(n1728), .O(n5570) );
  NAND_GATE U2531 ( .I1(n1705), .I2(donnee[11]), .O(n1728) );
  NAND_GATE U2532 ( .I1(\registres[6][11] ), .I2(n1706), .O(n1727) );
  NAND_GATE U2533 ( .I1(n1729), .I2(n1730), .O(n5571) );
  NAND_GATE U2534 ( .I1(n1705), .I2(donnee[12]), .O(n1730) );
  NAND_GATE U2535 ( .I1(\registres[6][12] ), .I2(n1706), .O(n1729) );
  NAND_GATE U2536 ( .I1(n1731), .I2(n1732), .O(n5572) );
  NAND_GATE U2537 ( .I1(n1705), .I2(donnee[13]), .O(n1732) );
  NAND_GATE U2538 ( .I1(\registres[6][13] ), .I2(n1706), .O(n1731) );
  NAND_GATE U2539 ( .I1(n1733), .I2(n1734), .O(n5573) );
  NAND_GATE U2540 ( .I1(n1705), .I2(donnee[14]), .O(n1734) );
  NAND_GATE U2541 ( .I1(\registres[6][14] ), .I2(n1706), .O(n1733) );
  NAND_GATE U2542 ( .I1(n1735), .I2(n1736), .O(n5574) );
  NAND_GATE U2543 ( .I1(n1705), .I2(donnee[15]), .O(n1736) );
  NAND_GATE U2544 ( .I1(\registres[6][15] ), .I2(n1706), .O(n1735) );
  NAND_GATE U2545 ( .I1(n1737), .I2(n1738), .O(n5575) );
  NAND_GATE U2546 ( .I1(n1705), .I2(donnee[16]), .O(n1738) );
  NAND_GATE U2547 ( .I1(\registres[6][16] ), .I2(n1706), .O(n1737) );
  NAND_GATE U2548 ( .I1(n1739), .I2(n1740), .O(n5576) );
  NAND_GATE U2549 ( .I1(n1705), .I2(donnee[17]), .O(n1740) );
  NAND_GATE U2550 ( .I1(\registres[6][17] ), .I2(n1706), .O(n1739) );
  NAND_GATE U2551 ( .I1(n1741), .I2(n1742), .O(n5577) );
  NAND_GATE U2552 ( .I1(n1705), .I2(donnee[18]), .O(n1742) );
  NAND_GATE U2553 ( .I1(\registres[6][18] ), .I2(n1706), .O(n1741) );
  NAND_GATE U2554 ( .I1(n1743), .I2(n1744), .O(n5578) );
  NAND_GATE U2555 ( .I1(n1705), .I2(donnee[19]), .O(n1744) );
  NAND_GATE U2556 ( .I1(\registres[6][19] ), .I2(n1706), .O(n1743) );
  NAND_GATE U2557 ( .I1(n1745), .I2(n1746), .O(n5579) );
  NAND_GATE U2558 ( .I1(n1705), .I2(donnee[20]), .O(n1746) );
  NAND_GATE U2559 ( .I1(\registres[6][20] ), .I2(n1706), .O(n1745) );
  NAND_GATE U2560 ( .I1(n1747), .I2(n1748), .O(n5580) );
  NAND_GATE U2561 ( .I1(n1705), .I2(donnee[21]), .O(n1748) );
  NAND_GATE U2562 ( .I1(\registres[6][21] ), .I2(n1706), .O(n1747) );
  NAND_GATE U2563 ( .I1(n1749), .I2(n1750), .O(n5581) );
  NAND_GATE U2564 ( .I1(n1705), .I2(donnee[22]), .O(n1750) );
  NAND_GATE U2565 ( .I1(\registres[6][22] ), .I2(n1706), .O(n1749) );
  NAND_GATE U2566 ( .I1(n1751), .I2(n1752), .O(n5582) );
  NAND_GATE U2567 ( .I1(n1705), .I2(donnee[23]), .O(n1752) );
  NAND_GATE U2568 ( .I1(\registres[6][23] ), .I2(n1706), .O(n1751) );
  NAND_GATE U2569 ( .I1(n1753), .I2(n1754), .O(n5583) );
  NAND_GATE U2570 ( .I1(n1705), .I2(donnee[24]), .O(n1754) );
  NAND_GATE U2571 ( .I1(\registres[6][24] ), .I2(n1706), .O(n1753) );
  NAND_GATE U2572 ( .I1(n1755), .I2(n1756), .O(n5584) );
  NAND_GATE U2573 ( .I1(n1705), .I2(donnee[25]), .O(n1756) );
  NAND_GATE U2574 ( .I1(\registres[6][25] ), .I2(n1706), .O(n1755) );
  NAND_GATE U2575 ( .I1(n1757), .I2(n1758), .O(n5585) );
  NAND_GATE U2576 ( .I1(n1705), .I2(donnee[26]), .O(n1758) );
  NAND_GATE U2577 ( .I1(\registres[6][26] ), .I2(n1706), .O(n1757) );
  NAND_GATE U2578 ( .I1(n1759), .I2(n1760), .O(n5586) );
  NAND_GATE U2579 ( .I1(n1705), .I2(donnee[27]), .O(n1760) );
  NAND_GATE U2580 ( .I1(\registres[6][27] ), .I2(n1706), .O(n1759) );
  NAND_GATE U2581 ( .I1(n1761), .I2(n1762), .O(n5587) );
  NAND_GATE U2582 ( .I1(n1705), .I2(donnee[28]), .O(n1762) );
  NAND_GATE U2583 ( .I1(\registres[6][28] ), .I2(n1706), .O(n1761) );
  NAND_GATE U2584 ( .I1(n1763), .I2(n1764), .O(n5588) );
  NAND_GATE U2585 ( .I1(n1705), .I2(donnee[29]), .O(n1764) );
  NAND_GATE U2586 ( .I1(\registres[6][29] ), .I2(n1706), .O(n1763) );
  NAND_GATE U2587 ( .I1(n1765), .I2(n1766), .O(n5589) );
  NAND_GATE U2588 ( .I1(n1705), .I2(donnee[30]), .O(n1766) );
  NAND_GATE U2589 ( .I1(\registres[6][30] ), .I2(n1706), .O(n1765) );
  NAND_GATE U2590 ( .I1(n1767), .I2(n1768), .O(n5590) );
  NAND_GATE U2591 ( .I1(n1705), .I2(donnee[31]), .O(n1768) );
  AND_GATE U2592 ( .I1(n1769), .I2(n1), .O(n1705) );
  NAND_GATE U2593 ( .I1(\registres[6][31] ), .I2(n1706), .O(n1767) );
  NOR_GATE U2594 ( .I1(n1769), .I2(reset), .O(n1706) );
  AND3_GATE U2595 ( .I1(n152), .I2(cmd_ecr), .I3(n1702), .O(n1769) );
  AND3_GATE U2596 ( .I1(reg_dest[1]), .I2(n4), .I3(reg_dest[2]), .O(n152) );
  NAND_GATE U2597 ( .I1(n1770), .I2(n1771), .O(n5591) );
  NAND_GATE U2598 ( .I1(n1772), .I2(donnee[0]), .O(n1771) );
  NAND_GATE U2599 ( .I1(\registres[5][0] ), .I2(n1773), .O(n1770) );
  NAND_GATE U2600 ( .I1(n1774), .I2(n1775), .O(n5592) );
  NAND_GATE U2601 ( .I1(n1772), .I2(donnee[1]), .O(n1775) );
  NAND_GATE U2602 ( .I1(\registres[5][1] ), .I2(n1773), .O(n1774) );
  NAND_GATE U2603 ( .I1(n1776), .I2(n1777), .O(n5593) );
  NAND_GATE U2604 ( .I1(n1772), .I2(donnee[2]), .O(n1777) );
  NAND_GATE U2605 ( .I1(\registres[5][2] ), .I2(n1773), .O(n1776) );
  NAND_GATE U2606 ( .I1(n1778), .I2(n1779), .O(n5594) );
  NAND_GATE U2607 ( .I1(n1772), .I2(donnee[3]), .O(n1779) );
  NAND_GATE U2608 ( .I1(\registres[5][3] ), .I2(n1773), .O(n1778) );
  NAND_GATE U2609 ( .I1(n1780), .I2(n1781), .O(n5595) );
  NAND_GATE U2610 ( .I1(n1772), .I2(donnee[4]), .O(n1781) );
  NAND_GATE U2611 ( .I1(\registres[5][4] ), .I2(n1773), .O(n1780) );
  NAND_GATE U2612 ( .I1(n1782), .I2(n1783), .O(n5596) );
  NAND_GATE U2613 ( .I1(n1772), .I2(donnee[5]), .O(n1783) );
  NAND_GATE U2614 ( .I1(\registres[5][5] ), .I2(n1773), .O(n1782) );
  NAND_GATE U2615 ( .I1(n1784), .I2(n1785), .O(n5597) );
  NAND_GATE U2616 ( .I1(n1772), .I2(donnee[6]), .O(n1785) );
  NAND_GATE U2617 ( .I1(\registres[5][6] ), .I2(n1773), .O(n1784) );
  NAND_GATE U2618 ( .I1(n1786), .I2(n1787), .O(n5598) );
  NAND_GATE U2619 ( .I1(n1772), .I2(donnee[7]), .O(n1787) );
  NAND_GATE U2620 ( .I1(\registres[5][7] ), .I2(n1773), .O(n1786) );
  NAND_GATE U2621 ( .I1(n1788), .I2(n1789), .O(n5599) );
  NAND_GATE U2622 ( .I1(n1772), .I2(donnee[8]), .O(n1789) );
  NAND_GATE U2623 ( .I1(\registres[5][8] ), .I2(n1773), .O(n1788) );
  NAND_GATE U2624 ( .I1(n1790), .I2(n1791), .O(n5600) );
  NAND_GATE U2625 ( .I1(n1772), .I2(donnee[9]), .O(n1791) );
  NAND_GATE U2626 ( .I1(\registres[5][9] ), .I2(n1773), .O(n1790) );
  NAND_GATE U2627 ( .I1(n1792), .I2(n1793), .O(n5601) );
  NAND_GATE U2628 ( .I1(n1772), .I2(donnee[10]), .O(n1793) );
  NAND_GATE U2629 ( .I1(\registres[5][10] ), .I2(n1773), .O(n1792) );
  NAND_GATE U2630 ( .I1(n1794), .I2(n1795), .O(n5602) );
  NAND_GATE U2631 ( .I1(n1772), .I2(donnee[11]), .O(n1795) );
  NAND_GATE U2632 ( .I1(\registres[5][11] ), .I2(n1773), .O(n1794) );
  NAND_GATE U2633 ( .I1(n1796), .I2(n1797), .O(n5603) );
  NAND_GATE U2634 ( .I1(n1772), .I2(donnee[12]), .O(n1797) );
  NAND_GATE U2635 ( .I1(\registres[5][12] ), .I2(n1773), .O(n1796) );
  NAND_GATE U2636 ( .I1(n1798), .I2(n1799), .O(n5604) );
  NAND_GATE U2637 ( .I1(n1772), .I2(donnee[13]), .O(n1799) );
  NAND_GATE U2638 ( .I1(\registres[5][13] ), .I2(n1773), .O(n1798) );
  NAND_GATE U2639 ( .I1(n1800), .I2(n1801), .O(n5605) );
  NAND_GATE U2640 ( .I1(n1772), .I2(donnee[14]), .O(n1801) );
  NAND_GATE U2641 ( .I1(\registres[5][14] ), .I2(n1773), .O(n1800) );
  NAND_GATE U2642 ( .I1(n1802), .I2(n1803), .O(n5606) );
  NAND_GATE U2643 ( .I1(n1772), .I2(donnee[15]), .O(n1803) );
  NAND_GATE U2644 ( .I1(\registres[5][15] ), .I2(n1773), .O(n1802) );
  NAND_GATE U2645 ( .I1(n1804), .I2(n1805), .O(n5607) );
  NAND_GATE U2646 ( .I1(n1772), .I2(donnee[16]), .O(n1805) );
  NAND_GATE U2647 ( .I1(\registres[5][16] ), .I2(n1773), .O(n1804) );
  NAND_GATE U2648 ( .I1(n1806), .I2(n1807), .O(n5608) );
  NAND_GATE U2649 ( .I1(n1772), .I2(donnee[17]), .O(n1807) );
  NAND_GATE U2650 ( .I1(\registres[5][17] ), .I2(n1773), .O(n1806) );
  NAND_GATE U2651 ( .I1(n1808), .I2(n1809), .O(n5609) );
  NAND_GATE U2652 ( .I1(n1772), .I2(donnee[18]), .O(n1809) );
  NAND_GATE U2653 ( .I1(\registres[5][18] ), .I2(n1773), .O(n1808) );
  NAND_GATE U2654 ( .I1(n1810), .I2(n1811), .O(n5610) );
  NAND_GATE U2655 ( .I1(n1772), .I2(donnee[19]), .O(n1811) );
  NAND_GATE U2656 ( .I1(\registres[5][19] ), .I2(n1773), .O(n1810) );
  NAND_GATE U2657 ( .I1(n1812), .I2(n1813), .O(n5611) );
  NAND_GATE U2658 ( .I1(n1772), .I2(donnee[20]), .O(n1813) );
  NAND_GATE U2659 ( .I1(\registres[5][20] ), .I2(n1773), .O(n1812) );
  NAND_GATE U2660 ( .I1(n1814), .I2(n1815), .O(n5612) );
  NAND_GATE U2661 ( .I1(n1772), .I2(donnee[21]), .O(n1815) );
  NAND_GATE U2662 ( .I1(\registres[5][21] ), .I2(n1773), .O(n1814) );
  NAND_GATE U2663 ( .I1(n1816), .I2(n1817), .O(n5613) );
  NAND_GATE U2664 ( .I1(n1772), .I2(donnee[22]), .O(n1817) );
  NAND_GATE U2665 ( .I1(\registres[5][22] ), .I2(n1773), .O(n1816) );
  NAND_GATE U2666 ( .I1(n1818), .I2(n1819), .O(n5614) );
  NAND_GATE U2667 ( .I1(n1772), .I2(donnee[23]), .O(n1819) );
  NAND_GATE U2668 ( .I1(\registres[5][23] ), .I2(n1773), .O(n1818) );
  NAND_GATE U2669 ( .I1(n1820), .I2(n1821), .O(n5615) );
  NAND_GATE U2670 ( .I1(n1772), .I2(donnee[24]), .O(n1821) );
  NAND_GATE U2671 ( .I1(\registres[5][24] ), .I2(n1773), .O(n1820) );
  NAND_GATE U2672 ( .I1(n1822), .I2(n1823), .O(n5616) );
  NAND_GATE U2673 ( .I1(n1772), .I2(donnee[25]), .O(n1823) );
  NAND_GATE U2674 ( .I1(\registres[5][25] ), .I2(n1773), .O(n1822) );
  NAND_GATE U2675 ( .I1(n1824), .I2(n1825), .O(n5617) );
  NAND_GATE U2676 ( .I1(n1772), .I2(donnee[26]), .O(n1825) );
  NAND_GATE U2677 ( .I1(\registres[5][26] ), .I2(n1773), .O(n1824) );
  NAND_GATE U2678 ( .I1(n1826), .I2(n1827), .O(n5618) );
  NAND_GATE U2679 ( .I1(n1772), .I2(donnee[27]), .O(n1827) );
  NAND_GATE U2680 ( .I1(\registres[5][27] ), .I2(n1773), .O(n1826) );
  NAND_GATE U2681 ( .I1(n1828), .I2(n1829), .O(n5619) );
  NAND_GATE U2682 ( .I1(n1772), .I2(donnee[28]), .O(n1829) );
  NAND_GATE U2683 ( .I1(\registres[5][28] ), .I2(n1773), .O(n1828) );
  NAND_GATE U2684 ( .I1(n1830), .I2(n1831), .O(n5620) );
  NAND_GATE U2685 ( .I1(n1772), .I2(donnee[29]), .O(n1831) );
  NAND_GATE U2686 ( .I1(\registres[5][29] ), .I2(n1773), .O(n1830) );
  NAND_GATE U2687 ( .I1(n1832), .I2(n1833), .O(n5621) );
  NAND_GATE U2688 ( .I1(n1772), .I2(donnee[30]), .O(n1833) );
  NAND_GATE U2689 ( .I1(\registres[5][30] ), .I2(n1773), .O(n1832) );
  NAND_GATE U2690 ( .I1(n1834), .I2(n1835), .O(n5622) );
  NAND_GATE U2691 ( .I1(n1772), .I2(donnee[31]), .O(n1835) );
  AND_GATE U2692 ( .I1(n1836), .I2(n1), .O(n1772) );
  NAND_GATE U2693 ( .I1(\registres[5][31] ), .I2(n1773), .O(n1834) );
  NOR_GATE U2694 ( .I1(n1836), .I2(reset), .O(n1773) );
  AND3_GATE U2695 ( .I1(n220), .I2(cmd_ecr), .I3(n1702), .O(n1836) );
  AND3_GATE U2696 ( .I1(reg_dest[0]), .I2(n3), .I3(reg_dest[2]), .O(n220) );
  NAND_GATE U2697 ( .I1(n1837), .I2(n1838), .O(n5623) );
  NAND_GATE U2698 ( .I1(n1839), .I2(donnee[0]), .O(n1838) );
  NAND_GATE U2699 ( .I1(\registres[4][0] ), .I2(n1840), .O(n1837) );
  NAND_GATE U2700 ( .I1(n1841), .I2(n1842), .O(n5624) );
  NAND_GATE U2701 ( .I1(n1839), .I2(donnee[1]), .O(n1842) );
  NAND_GATE U2702 ( .I1(\registres[4][1] ), .I2(n1840), .O(n1841) );
  NAND_GATE U2703 ( .I1(n1843), .I2(n1844), .O(n5625) );
  NAND_GATE U2704 ( .I1(n1839), .I2(donnee[2]), .O(n1844) );
  NAND_GATE U2705 ( .I1(\registres[4][2] ), .I2(n1840), .O(n1843) );
  NAND_GATE U2706 ( .I1(n1845), .I2(n1846), .O(n5626) );
  NAND_GATE U2707 ( .I1(n1839), .I2(donnee[3]), .O(n1846) );
  NAND_GATE U2708 ( .I1(\registres[4][3] ), .I2(n1840), .O(n1845) );
  NAND_GATE U2709 ( .I1(n1847), .I2(n1848), .O(n5627) );
  NAND_GATE U2710 ( .I1(n1839), .I2(donnee[4]), .O(n1848) );
  NAND_GATE U2711 ( .I1(\registres[4][4] ), .I2(n1840), .O(n1847) );
  NAND_GATE U2712 ( .I1(n1849), .I2(n1850), .O(n5628) );
  NAND_GATE U2713 ( .I1(n1839), .I2(donnee[5]), .O(n1850) );
  NAND_GATE U2714 ( .I1(\registres[4][5] ), .I2(n1840), .O(n1849) );
  NAND_GATE U2715 ( .I1(n1851), .I2(n1852), .O(n5629) );
  NAND_GATE U2716 ( .I1(n1839), .I2(donnee[6]), .O(n1852) );
  NAND_GATE U2717 ( .I1(\registres[4][6] ), .I2(n1840), .O(n1851) );
  NAND_GATE U2718 ( .I1(n1853), .I2(n1854), .O(n5630) );
  NAND_GATE U2719 ( .I1(n1839), .I2(donnee[7]), .O(n1854) );
  NAND_GATE U2720 ( .I1(\registres[4][7] ), .I2(n1840), .O(n1853) );
  NAND_GATE U2721 ( .I1(n1855), .I2(n1856), .O(n5631) );
  NAND_GATE U2722 ( .I1(n1839), .I2(donnee[8]), .O(n1856) );
  NAND_GATE U2723 ( .I1(\registres[4][8] ), .I2(n1840), .O(n1855) );
  NAND_GATE U2724 ( .I1(n1857), .I2(n1858), .O(n5632) );
  NAND_GATE U2725 ( .I1(n1839), .I2(donnee[9]), .O(n1858) );
  NAND_GATE U2726 ( .I1(\registres[4][9] ), .I2(n1840), .O(n1857) );
  NAND_GATE U2727 ( .I1(n1859), .I2(n1860), .O(n5633) );
  NAND_GATE U2728 ( .I1(n1839), .I2(donnee[10]), .O(n1860) );
  NAND_GATE U2729 ( .I1(\registres[4][10] ), .I2(n1840), .O(n1859) );
  NAND_GATE U2730 ( .I1(n1861), .I2(n1862), .O(n5634) );
  NAND_GATE U2731 ( .I1(n1839), .I2(donnee[11]), .O(n1862) );
  NAND_GATE U2732 ( .I1(\registres[4][11] ), .I2(n1840), .O(n1861) );
  NAND_GATE U2733 ( .I1(n1863), .I2(n1864), .O(n5635) );
  NAND_GATE U2734 ( .I1(n1839), .I2(donnee[12]), .O(n1864) );
  NAND_GATE U2735 ( .I1(\registres[4][12] ), .I2(n1840), .O(n1863) );
  NAND_GATE U2736 ( .I1(n1865), .I2(n1866), .O(n5636) );
  NAND_GATE U2737 ( .I1(n1839), .I2(donnee[13]), .O(n1866) );
  NAND_GATE U2738 ( .I1(\registres[4][13] ), .I2(n1840), .O(n1865) );
  NAND_GATE U2739 ( .I1(n1867), .I2(n1868), .O(n5637) );
  NAND_GATE U2740 ( .I1(n1839), .I2(donnee[14]), .O(n1868) );
  NAND_GATE U2741 ( .I1(\registres[4][14] ), .I2(n1840), .O(n1867) );
  NAND_GATE U2742 ( .I1(n1869), .I2(n1870), .O(n5638) );
  NAND_GATE U2743 ( .I1(n1839), .I2(donnee[15]), .O(n1870) );
  NAND_GATE U2744 ( .I1(\registres[4][15] ), .I2(n1840), .O(n1869) );
  NAND_GATE U2745 ( .I1(n1871), .I2(n1872), .O(n5639) );
  NAND_GATE U2746 ( .I1(n1839), .I2(donnee[16]), .O(n1872) );
  NAND_GATE U2747 ( .I1(\registres[4][16] ), .I2(n1840), .O(n1871) );
  NAND_GATE U2748 ( .I1(n1873), .I2(n1874), .O(n5640) );
  NAND_GATE U2749 ( .I1(n1839), .I2(donnee[17]), .O(n1874) );
  NAND_GATE U2750 ( .I1(\registres[4][17] ), .I2(n1840), .O(n1873) );
  NAND_GATE U2751 ( .I1(n1875), .I2(n1876), .O(n5641) );
  NAND_GATE U2752 ( .I1(n1839), .I2(donnee[18]), .O(n1876) );
  NAND_GATE U2753 ( .I1(\registres[4][18] ), .I2(n1840), .O(n1875) );
  NAND_GATE U2754 ( .I1(n1877), .I2(n1878), .O(n5642) );
  NAND_GATE U2755 ( .I1(n1839), .I2(donnee[19]), .O(n1878) );
  NAND_GATE U2756 ( .I1(\registres[4][19] ), .I2(n1840), .O(n1877) );
  NAND_GATE U2757 ( .I1(n1879), .I2(n1880), .O(n5643) );
  NAND_GATE U2758 ( .I1(n1839), .I2(donnee[20]), .O(n1880) );
  NAND_GATE U2759 ( .I1(\registres[4][20] ), .I2(n1840), .O(n1879) );
  NAND_GATE U2760 ( .I1(n1881), .I2(n1882), .O(n5644) );
  NAND_GATE U2761 ( .I1(n1839), .I2(donnee[21]), .O(n1882) );
  NAND_GATE U2762 ( .I1(\registres[4][21] ), .I2(n1840), .O(n1881) );
  NAND_GATE U2763 ( .I1(n1883), .I2(n1884), .O(n5645) );
  NAND_GATE U2764 ( .I1(n1839), .I2(donnee[22]), .O(n1884) );
  NAND_GATE U2765 ( .I1(\registres[4][22] ), .I2(n1840), .O(n1883) );
  NAND_GATE U2766 ( .I1(n1885), .I2(n1886), .O(n5646) );
  NAND_GATE U2767 ( .I1(n1839), .I2(donnee[23]), .O(n1886) );
  NAND_GATE U2768 ( .I1(\registres[4][23] ), .I2(n1840), .O(n1885) );
  NAND_GATE U2769 ( .I1(n1887), .I2(n1888), .O(n5647) );
  NAND_GATE U2770 ( .I1(n1839), .I2(donnee[24]), .O(n1888) );
  NAND_GATE U2771 ( .I1(\registres[4][24] ), .I2(n1840), .O(n1887) );
  NAND_GATE U2772 ( .I1(n1889), .I2(n1890), .O(n5648) );
  NAND_GATE U2773 ( .I1(n1839), .I2(donnee[25]), .O(n1890) );
  NAND_GATE U2774 ( .I1(\registres[4][25] ), .I2(n1840), .O(n1889) );
  NAND_GATE U2775 ( .I1(n1891), .I2(n1892), .O(n5649) );
  NAND_GATE U2776 ( .I1(n1839), .I2(donnee[26]), .O(n1892) );
  NAND_GATE U2777 ( .I1(\registres[4][26] ), .I2(n1840), .O(n1891) );
  NAND_GATE U2778 ( .I1(n1893), .I2(n1894), .O(n5650) );
  NAND_GATE U2779 ( .I1(n1839), .I2(donnee[27]), .O(n1894) );
  NAND_GATE U2780 ( .I1(\registres[4][27] ), .I2(n1840), .O(n1893) );
  NAND_GATE U2781 ( .I1(n1895), .I2(n1896), .O(n5651) );
  NAND_GATE U2782 ( .I1(n1839), .I2(donnee[28]), .O(n1896) );
  NAND_GATE U2783 ( .I1(\registres[4][28] ), .I2(n1840), .O(n1895) );
  NAND_GATE U2784 ( .I1(n1897), .I2(n1898), .O(n5652) );
  NAND_GATE U2785 ( .I1(n1839), .I2(donnee[29]), .O(n1898) );
  NAND_GATE U2786 ( .I1(\registres[4][29] ), .I2(n1840), .O(n1897) );
  NAND_GATE U2787 ( .I1(n1899), .I2(n1900), .O(n5653) );
  NAND_GATE U2788 ( .I1(n1839), .I2(donnee[30]), .O(n1900) );
  NAND_GATE U2789 ( .I1(\registres[4][30] ), .I2(n1840), .O(n1899) );
  NAND_GATE U2790 ( .I1(n1901), .I2(n1902), .O(n5654) );
  NAND_GATE U2791 ( .I1(n1839), .I2(donnee[31]), .O(n1902) );
  AND_GATE U2792 ( .I1(n1903), .I2(n1), .O(n1839) );
  NAND_GATE U2793 ( .I1(\registres[4][31] ), .I2(n1840), .O(n1901) );
  NOR_GATE U2794 ( .I1(n1903), .I2(reset), .O(n1840) );
  AND3_GATE U2795 ( .I1(n288), .I2(cmd_ecr), .I3(n1702), .O(n1903) );
  AND3_GATE U2796 ( .I1(n4), .I2(n3), .I3(reg_dest[2]), .O(n288) );
  NAND_GATE U2797 ( .I1(n1904), .I2(n1905), .O(n5655) );
  NAND_GATE U2798 ( .I1(n1906), .I2(donnee[0]), .O(n1905) );
  NAND_GATE U2799 ( .I1(\registres[3][0] ), .I2(n1907), .O(n1904) );
  NAND_GATE U2800 ( .I1(n1908), .I2(n1909), .O(n5656) );
  NAND_GATE U2801 ( .I1(n1906), .I2(donnee[1]), .O(n1909) );
  NAND_GATE U2802 ( .I1(\registres[3][1] ), .I2(n1907), .O(n1908) );
  NAND_GATE U2803 ( .I1(n1910), .I2(n1911), .O(n5657) );
  NAND_GATE U2804 ( .I1(n1906), .I2(donnee[2]), .O(n1911) );
  NAND_GATE U2805 ( .I1(\registres[3][2] ), .I2(n1907), .O(n1910) );
  NAND_GATE U2806 ( .I1(n1912), .I2(n1913), .O(n5658) );
  NAND_GATE U2807 ( .I1(n1906), .I2(donnee[3]), .O(n1913) );
  NAND_GATE U2808 ( .I1(\registres[3][3] ), .I2(n1907), .O(n1912) );
  NAND_GATE U2809 ( .I1(n1914), .I2(n1915), .O(n5659) );
  NAND_GATE U2810 ( .I1(n1906), .I2(donnee[4]), .O(n1915) );
  NAND_GATE U2811 ( .I1(\registres[3][4] ), .I2(n1907), .O(n1914) );
  NAND_GATE U2812 ( .I1(n1916), .I2(n1917), .O(n5660) );
  NAND_GATE U2813 ( .I1(n1906), .I2(donnee[5]), .O(n1917) );
  NAND_GATE U2814 ( .I1(\registres[3][5] ), .I2(n1907), .O(n1916) );
  NAND_GATE U2815 ( .I1(n1918), .I2(n1919), .O(n5661) );
  NAND_GATE U2816 ( .I1(n1906), .I2(donnee[6]), .O(n1919) );
  NAND_GATE U2817 ( .I1(\registres[3][6] ), .I2(n1907), .O(n1918) );
  NAND_GATE U2818 ( .I1(n1920), .I2(n1921), .O(n5662) );
  NAND_GATE U2819 ( .I1(n1906), .I2(donnee[7]), .O(n1921) );
  NAND_GATE U2820 ( .I1(\registres[3][7] ), .I2(n1907), .O(n1920) );
  NAND_GATE U2821 ( .I1(n1922), .I2(n1923), .O(n5663) );
  NAND_GATE U2822 ( .I1(n1906), .I2(donnee[8]), .O(n1923) );
  NAND_GATE U2823 ( .I1(\registres[3][8] ), .I2(n1907), .O(n1922) );
  NAND_GATE U2824 ( .I1(n1924), .I2(n1925), .O(n5664) );
  NAND_GATE U2825 ( .I1(n1906), .I2(donnee[9]), .O(n1925) );
  NAND_GATE U2826 ( .I1(\registres[3][9] ), .I2(n1907), .O(n1924) );
  NAND_GATE U2827 ( .I1(n1926), .I2(n1927), .O(n5665) );
  NAND_GATE U2828 ( .I1(n1906), .I2(donnee[10]), .O(n1927) );
  NAND_GATE U2829 ( .I1(\registres[3][10] ), .I2(n1907), .O(n1926) );
  NAND_GATE U2830 ( .I1(n1928), .I2(n1929), .O(n5666) );
  NAND_GATE U2831 ( .I1(n1906), .I2(donnee[11]), .O(n1929) );
  NAND_GATE U2832 ( .I1(\registres[3][11] ), .I2(n1907), .O(n1928) );
  NAND_GATE U2833 ( .I1(n1930), .I2(n1931), .O(n5667) );
  NAND_GATE U2834 ( .I1(n1906), .I2(donnee[12]), .O(n1931) );
  NAND_GATE U2835 ( .I1(\registres[3][12] ), .I2(n1907), .O(n1930) );
  NAND_GATE U2836 ( .I1(n1932), .I2(n1933), .O(n5668) );
  NAND_GATE U2837 ( .I1(n1906), .I2(donnee[13]), .O(n1933) );
  NAND_GATE U2838 ( .I1(\registres[3][13] ), .I2(n1907), .O(n1932) );
  NAND_GATE U2839 ( .I1(n1934), .I2(n1935), .O(n5669) );
  NAND_GATE U2840 ( .I1(n1906), .I2(donnee[14]), .O(n1935) );
  NAND_GATE U2841 ( .I1(\registres[3][14] ), .I2(n1907), .O(n1934) );
  NAND_GATE U2842 ( .I1(n1936), .I2(n1937), .O(n5670) );
  NAND_GATE U2843 ( .I1(n1906), .I2(donnee[15]), .O(n1937) );
  NAND_GATE U2844 ( .I1(\registres[3][15] ), .I2(n1907), .O(n1936) );
  NAND_GATE U2845 ( .I1(n1938), .I2(n1939), .O(n5671) );
  NAND_GATE U2846 ( .I1(n1906), .I2(donnee[16]), .O(n1939) );
  NAND_GATE U2847 ( .I1(\registres[3][16] ), .I2(n1907), .O(n1938) );
  NAND_GATE U2848 ( .I1(n1940), .I2(n1941), .O(n5672) );
  NAND_GATE U2849 ( .I1(n1906), .I2(donnee[17]), .O(n1941) );
  NAND_GATE U2850 ( .I1(\registres[3][17] ), .I2(n1907), .O(n1940) );
  NAND_GATE U2851 ( .I1(n1942), .I2(n1943), .O(n5673) );
  NAND_GATE U2852 ( .I1(n1906), .I2(donnee[18]), .O(n1943) );
  NAND_GATE U2853 ( .I1(\registres[3][18] ), .I2(n1907), .O(n1942) );
  NAND_GATE U2854 ( .I1(n1944), .I2(n1945), .O(n5674) );
  NAND_GATE U2855 ( .I1(n1906), .I2(donnee[19]), .O(n1945) );
  NAND_GATE U2856 ( .I1(\registres[3][19] ), .I2(n1907), .O(n1944) );
  NAND_GATE U2857 ( .I1(n1946), .I2(n1947), .O(n5675) );
  NAND_GATE U2858 ( .I1(n1906), .I2(donnee[20]), .O(n1947) );
  NAND_GATE U2859 ( .I1(\registres[3][20] ), .I2(n1907), .O(n1946) );
  NAND_GATE U2860 ( .I1(n1948), .I2(n1949), .O(n5676) );
  NAND_GATE U2861 ( .I1(n1906), .I2(donnee[21]), .O(n1949) );
  NAND_GATE U2862 ( .I1(\registres[3][21] ), .I2(n1907), .O(n1948) );
  NAND_GATE U2863 ( .I1(n1950), .I2(n1951), .O(n5677) );
  NAND_GATE U2864 ( .I1(n1906), .I2(donnee[22]), .O(n1951) );
  NAND_GATE U2865 ( .I1(\registres[3][22] ), .I2(n1907), .O(n1950) );
  NAND_GATE U2866 ( .I1(n1952), .I2(n1953), .O(n5678) );
  NAND_GATE U2867 ( .I1(n1906), .I2(donnee[23]), .O(n1953) );
  NAND_GATE U2868 ( .I1(\registres[3][23] ), .I2(n1907), .O(n1952) );
  NAND_GATE U2869 ( .I1(n1954), .I2(n1955), .O(n5679) );
  NAND_GATE U2870 ( .I1(n1906), .I2(donnee[24]), .O(n1955) );
  NAND_GATE U2871 ( .I1(\registres[3][24] ), .I2(n1907), .O(n1954) );
  NAND_GATE U2872 ( .I1(n1956), .I2(n1957), .O(n5680) );
  NAND_GATE U2873 ( .I1(n1906), .I2(donnee[25]), .O(n1957) );
  NAND_GATE U2874 ( .I1(\registres[3][25] ), .I2(n1907), .O(n1956) );
  NAND_GATE U2875 ( .I1(n1958), .I2(n1959), .O(n5681) );
  NAND_GATE U2876 ( .I1(n1906), .I2(donnee[26]), .O(n1959) );
  NAND_GATE U2877 ( .I1(\registres[3][26] ), .I2(n1907), .O(n1958) );
  NAND_GATE U2878 ( .I1(n1960), .I2(n1961), .O(n5682) );
  NAND_GATE U2879 ( .I1(n1906), .I2(donnee[27]), .O(n1961) );
  NAND_GATE U2880 ( .I1(\registres[3][27] ), .I2(n1907), .O(n1960) );
  NAND_GATE U2881 ( .I1(n1962), .I2(n1963), .O(n5683) );
  NAND_GATE U2882 ( .I1(n1906), .I2(donnee[28]), .O(n1963) );
  NAND_GATE U2883 ( .I1(\registres[3][28] ), .I2(n1907), .O(n1962) );
  NAND_GATE U2884 ( .I1(n1964), .I2(n1965), .O(n5684) );
  NAND_GATE U2885 ( .I1(n1906), .I2(donnee[29]), .O(n1965) );
  NAND_GATE U2886 ( .I1(\registres[3][29] ), .I2(n1907), .O(n1964) );
  NAND_GATE U2887 ( .I1(n1966), .I2(n1967), .O(n5685) );
  NAND_GATE U2888 ( .I1(n1906), .I2(donnee[30]), .O(n1967) );
  NAND_GATE U2889 ( .I1(\registres[3][30] ), .I2(n1907), .O(n1966) );
  NAND_GATE U2890 ( .I1(n1968), .I2(n1969), .O(n5686) );
  NAND_GATE U2891 ( .I1(n1906), .I2(donnee[31]), .O(n1969) );
  AND_GATE U2892 ( .I1(n1970), .I2(n1), .O(n1906) );
  NAND_GATE U2893 ( .I1(\registres[3][31] ), .I2(n1907), .O(n1968) );
  NOR_GATE U2894 ( .I1(n1970), .I2(reset), .O(n1907) );
  AND3_GATE U2895 ( .I1(n356), .I2(cmd_ecr), .I3(n1702), .O(n1970) );
  NOR3_GATE U2896 ( .I1(n4), .I2(reg_dest[2]), .I3(n3), .O(n356) );
  NAND_GATE U2897 ( .I1(n1971), .I2(n1972), .O(n5687) );
  NAND_GATE U2898 ( .I1(n1973), .I2(donnee[0]), .O(n1972) );
  NAND_GATE U2899 ( .I1(\registres[2][0] ), .I2(n1974), .O(n1971) );
  NAND_GATE U2900 ( .I1(n1975), .I2(n1976), .O(n5688) );
  NAND_GATE U2901 ( .I1(n1973), .I2(donnee[1]), .O(n1976) );
  NAND_GATE U2902 ( .I1(\registres[2][1] ), .I2(n1974), .O(n1975) );
  NAND_GATE U2903 ( .I1(n1977), .I2(n1978), .O(n5689) );
  NAND_GATE U2904 ( .I1(n1973), .I2(donnee[2]), .O(n1978) );
  NAND_GATE U2905 ( .I1(\registres[2][2] ), .I2(n1974), .O(n1977) );
  NAND_GATE U2906 ( .I1(n1979), .I2(n1980), .O(n5690) );
  NAND_GATE U2907 ( .I1(n1973), .I2(donnee[3]), .O(n1980) );
  NAND_GATE U2908 ( .I1(\registres[2][3] ), .I2(n1974), .O(n1979) );
  NAND_GATE U2909 ( .I1(n1981), .I2(n1982), .O(n5691) );
  NAND_GATE U2910 ( .I1(n1973), .I2(donnee[4]), .O(n1982) );
  NAND_GATE U2911 ( .I1(\registres[2][4] ), .I2(n1974), .O(n1981) );
  NAND_GATE U2912 ( .I1(n1983), .I2(n1984), .O(n5692) );
  NAND_GATE U2913 ( .I1(n1973), .I2(donnee[5]), .O(n1984) );
  NAND_GATE U2914 ( .I1(\registres[2][5] ), .I2(n1974), .O(n1983) );
  NAND_GATE U2915 ( .I1(n1985), .I2(n1986), .O(n5693) );
  NAND_GATE U2916 ( .I1(n1973), .I2(donnee[6]), .O(n1986) );
  NAND_GATE U2917 ( .I1(\registres[2][6] ), .I2(n1974), .O(n1985) );
  NAND_GATE U2918 ( .I1(n1987), .I2(n1988), .O(n5694) );
  NAND_GATE U2919 ( .I1(n1973), .I2(donnee[7]), .O(n1988) );
  NAND_GATE U2920 ( .I1(\registres[2][7] ), .I2(n1974), .O(n1987) );
  NAND_GATE U2921 ( .I1(n1989), .I2(n1990), .O(n5695) );
  NAND_GATE U2922 ( .I1(n1973), .I2(donnee[8]), .O(n1990) );
  NAND_GATE U2923 ( .I1(\registres[2][8] ), .I2(n1974), .O(n1989) );
  NAND_GATE U2924 ( .I1(n1991), .I2(n1992), .O(n5696) );
  NAND_GATE U2925 ( .I1(n1973), .I2(donnee[9]), .O(n1992) );
  NAND_GATE U2926 ( .I1(\registres[2][9] ), .I2(n1974), .O(n1991) );
  NAND_GATE U2927 ( .I1(n1993), .I2(n1994), .O(n5697) );
  NAND_GATE U2928 ( .I1(n1973), .I2(donnee[10]), .O(n1994) );
  NAND_GATE U2929 ( .I1(\registres[2][10] ), .I2(n1974), .O(n1993) );
  NAND_GATE U2930 ( .I1(n1995), .I2(n1996), .O(n5698) );
  NAND_GATE U2931 ( .I1(n1973), .I2(donnee[11]), .O(n1996) );
  NAND_GATE U2932 ( .I1(\registres[2][11] ), .I2(n1974), .O(n1995) );
  NAND_GATE U2933 ( .I1(n1997), .I2(n1998), .O(n5699) );
  NAND_GATE U2934 ( .I1(n1973), .I2(donnee[12]), .O(n1998) );
  NAND_GATE U2935 ( .I1(\registres[2][12] ), .I2(n1974), .O(n1997) );
  NAND_GATE U2936 ( .I1(n1999), .I2(n2000), .O(n5700) );
  NAND_GATE U2937 ( .I1(n1973), .I2(donnee[13]), .O(n2000) );
  NAND_GATE U2938 ( .I1(\registres[2][13] ), .I2(n1974), .O(n1999) );
  NAND_GATE U2939 ( .I1(n2001), .I2(n2002), .O(n5701) );
  NAND_GATE U2940 ( .I1(n1973), .I2(donnee[14]), .O(n2002) );
  NAND_GATE U2941 ( .I1(\registres[2][14] ), .I2(n1974), .O(n2001) );
  NAND_GATE U2942 ( .I1(n2003), .I2(n2004), .O(n5702) );
  NAND_GATE U2943 ( .I1(n1973), .I2(donnee[15]), .O(n2004) );
  NAND_GATE U2944 ( .I1(\registres[2][15] ), .I2(n1974), .O(n2003) );
  NAND_GATE U2945 ( .I1(n2005), .I2(n2006), .O(n5703) );
  NAND_GATE U2946 ( .I1(n1973), .I2(donnee[16]), .O(n2006) );
  NAND_GATE U2947 ( .I1(\registres[2][16] ), .I2(n1974), .O(n2005) );
  NAND_GATE U2948 ( .I1(n2007), .I2(n2008), .O(n5704) );
  NAND_GATE U2949 ( .I1(n1973), .I2(donnee[17]), .O(n2008) );
  NAND_GATE U2950 ( .I1(\registres[2][17] ), .I2(n1974), .O(n2007) );
  NAND_GATE U2951 ( .I1(n2009), .I2(n2010), .O(n5705) );
  NAND_GATE U2952 ( .I1(n1973), .I2(donnee[18]), .O(n2010) );
  NAND_GATE U2953 ( .I1(\registres[2][18] ), .I2(n1974), .O(n2009) );
  NAND_GATE U2954 ( .I1(n2011), .I2(n2012), .O(n5706) );
  NAND_GATE U2955 ( .I1(n1973), .I2(donnee[19]), .O(n2012) );
  NAND_GATE U2956 ( .I1(\registres[2][19] ), .I2(n1974), .O(n2011) );
  NAND_GATE U2957 ( .I1(n2013), .I2(n2014), .O(n5707) );
  NAND_GATE U2958 ( .I1(n1973), .I2(donnee[20]), .O(n2014) );
  NAND_GATE U2959 ( .I1(\registres[2][20] ), .I2(n1974), .O(n2013) );
  NAND_GATE U2960 ( .I1(n2015), .I2(n2016), .O(n5708) );
  NAND_GATE U2961 ( .I1(n1973), .I2(donnee[21]), .O(n2016) );
  NAND_GATE U2962 ( .I1(\registres[2][21] ), .I2(n1974), .O(n2015) );
  NAND_GATE U2963 ( .I1(n2017), .I2(n2018), .O(n5709) );
  NAND_GATE U2964 ( .I1(n1973), .I2(donnee[22]), .O(n2018) );
  NAND_GATE U2965 ( .I1(\registres[2][22] ), .I2(n1974), .O(n2017) );
  NAND_GATE U2966 ( .I1(n2019), .I2(n2020), .O(n5710) );
  NAND_GATE U2967 ( .I1(n1973), .I2(donnee[23]), .O(n2020) );
  NAND_GATE U2968 ( .I1(\registres[2][23] ), .I2(n1974), .O(n2019) );
  NAND_GATE U2969 ( .I1(n2021), .I2(n2022), .O(n5711) );
  NAND_GATE U2970 ( .I1(n1973), .I2(donnee[24]), .O(n2022) );
  NAND_GATE U2971 ( .I1(\registres[2][24] ), .I2(n1974), .O(n2021) );
  NAND_GATE U2972 ( .I1(n2023), .I2(n2024), .O(n5712) );
  NAND_GATE U2973 ( .I1(n1973), .I2(donnee[25]), .O(n2024) );
  NAND_GATE U2974 ( .I1(\registres[2][25] ), .I2(n1974), .O(n2023) );
  NAND_GATE U2975 ( .I1(n2025), .I2(n2026), .O(n5713) );
  NAND_GATE U2976 ( .I1(n1973), .I2(donnee[26]), .O(n2026) );
  NAND_GATE U2977 ( .I1(\registres[2][26] ), .I2(n1974), .O(n2025) );
  NAND_GATE U2978 ( .I1(n2027), .I2(n2028), .O(n5714) );
  NAND_GATE U2979 ( .I1(n1973), .I2(donnee[27]), .O(n2028) );
  NAND_GATE U2980 ( .I1(\registres[2][27] ), .I2(n1974), .O(n2027) );
  NAND_GATE U2981 ( .I1(n2029), .I2(n2030), .O(n5715) );
  NAND_GATE U2982 ( .I1(n1973), .I2(donnee[28]), .O(n2030) );
  NAND_GATE U2983 ( .I1(\registres[2][28] ), .I2(n1974), .O(n2029) );
  NAND_GATE U2984 ( .I1(n2031), .I2(n2032), .O(n5716) );
  NAND_GATE U2985 ( .I1(n1973), .I2(donnee[29]), .O(n2032) );
  NAND_GATE U2986 ( .I1(\registres[2][29] ), .I2(n1974), .O(n2031) );
  NAND_GATE U2987 ( .I1(n2033), .I2(n2034), .O(n5717) );
  NAND_GATE U2988 ( .I1(n1973), .I2(donnee[30]), .O(n2034) );
  NAND_GATE U2989 ( .I1(\registres[2][30] ), .I2(n1974), .O(n2033) );
  NAND_GATE U2990 ( .I1(n2035), .I2(n2036), .O(n5718) );
  NAND_GATE U2991 ( .I1(n1973), .I2(donnee[31]), .O(n2036) );
  AND_GATE U2992 ( .I1(n2037), .I2(n1), .O(n1973) );
  NAND_GATE U2993 ( .I1(\registres[2][31] ), .I2(n1974), .O(n2035) );
  NOR_GATE U2994 ( .I1(n2037), .I2(reset), .O(n1974) );
  AND3_GATE U2995 ( .I1(n424), .I2(cmd_ecr), .I3(n1702), .O(n2037) );
  NOR3_GATE U2996 ( .I1(reg_dest[0]), .I2(reg_dest[2]), .I3(n3), .O(n424) );
  NAND_GATE U2997 ( .I1(n2038), .I2(n2039), .O(n5719) );
  NAND_GATE U2998 ( .I1(n2040), .I2(donnee[0]), .O(n2039) );
  NAND_GATE U2999 ( .I1(\registres[1][0] ), .I2(n2041), .O(n2038) );
  NAND_GATE U3000 ( .I1(n2042), .I2(n2043), .O(n5720) );
  NAND_GATE U3001 ( .I1(n2040), .I2(donnee[1]), .O(n2043) );
  NAND_GATE U3002 ( .I1(\registres[1][1] ), .I2(n2041), .O(n2042) );
  NAND_GATE U3003 ( .I1(n2044), .I2(n2045), .O(n5721) );
  NAND_GATE U3004 ( .I1(n2040), .I2(donnee[2]), .O(n2045) );
  NAND_GATE U3005 ( .I1(\registres[1][2] ), .I2(n2041), .O(n2044) );
  NAND_GATE U3006 ( .I1(n2046), .I2(n2047), .O(n5722) );
  NAND_GATE U3007 ( .I1(n2040), .I2(donnee[3]), .O(n2047) );
  NAND_GATE U3008 ( .I1(\registres[1][3] ), .I2(n2041), .O(n2046) );
  NAND_GATE U3009 ( .I1(n2048), .I2(n2049), .O(n5723) );
  NAND_GATE U3010 ( .I1(n2040), .I2(donnee[4]), .O(n2049) );
  NAND_GATE U3011 ( .I1(\registres[1][4] ), .I2(n2041), .O(n2048) );
  NAND_GATE U3012 ( .I1(n2050), .I2(n2051), .O(n5724) );
  NAND_GATE U3013 ( .I1(n2040), .I2(donnee[5]), .O(n2051) );
  NAND_GATE U3014 ( .I1(\registres[1][5] ), .I2(n2041), .O(n2050) );
  NAND_GATE U3015 ( .I1(n2052), .I2(n2053), .O(n5725) );
  NAND_GATE U3016 ( .I1(n2040), .I2(donnee[6]), .O(n2053) );
  NAND_GATE U3017 ( .I1(\registres[1][6] ), .I2(n2041), .O(n2052) );
  NAND_GATE U3018 ( .I1(n2054), .I2(n2055), .O(n5726) );
  NAND_GATE U3019 ( .I1(n2040), .I2(donnee[7]), .O(n2055) );
  NAND_GATE U3020 ( .I1(\registres[1][7] ), .I2(n2041), .O(n2054) );
  NAND_GATE U3021 ( .I1(n2056), .I2(n2057), .O(n5727) );
  NAND_GATE U3022 ( .I1(n2040), .I2(donnee[8]), .O(n2057) );
  NAND_GATE U3023 ( .I1(\registres[1][8] ), .I2(n2041), .O(n2056) );
  NAND_GATE U3024 ( .I1(n2058), .I2(n2059), .O(n5728) );
  NAND_GATE U3025 ( .I1(n2040), .I2(donnee[9]), .O(n2059) );
  NAND_GATE U3026 ( .I1(\registres[1][9] ), .I2(n2041), .O(n2058) );
  NAND_GATE U3027 ( .I1(n2060), .I2(n2061), .O(n5729) );
  NAND_GATE U3028 ( .I1(n2040), .I2(donnee[10]), .O(n2061) );
  NAND_GATE U3029 ( .I1(\registres[1][10] ), .I2(n2041), .O(n2060) );
  NAND_GATE U3030 ( .I1(n2062), .I2(n2063), .O(n5730) );
  NAND_GATE U3031 ( .I1(n2040), .I2(donnee[11]), .O(n2063) );
  NAND_GATE U3032 ( .I1(\registres[1][11] ), .I2(n2041), .O(n2062) );
  NAND_GATE U3033 ( .I1(n2064), .I2(n2065), .O(n5731) );
  NAND_GATE U3034 ( .I1(n2040), .I2(donnee[12]), .O(n2065) );
  NAND_GATE U3035 ( .I1(\registres[1][12] ), .I2(n2041), .O(n2064) );
  NAND_GATE U3036 ( .I1(n2066), .I2(n2067), .O(n5732) );
  NAND_GATE U3037 ( .I1(n2040), .I2(donnee[13]), .O(n2067) );
  NAND_GATE U3038 ( .I1(\registres[1][13] ), .I2(n2041), .O(n2066) );
  NAND_GATE U3039 ( .I1(n2068), .I2(n2069), .O(n5733) );
  NAND_GATE U3040 ( .I1(n2040), .I2(donnee[14]), .O(n2069) );
  NAND_GATE U3041 ( .I1(\registres[1][14] ), .I2(n2041), .O(n2068) );
  NAND_GATE U3042 ( .I1(n2070), .I2(n2071), .O(n5734) );
  NAND_GATE U3043 ( .I1(n2040), .I2(donnee[15]), .O(n2071) );
  NAND_GATE U3044 ( .I1(\registres[1][15] ), .I2(n2041), .O(n2070) );
  NAND_GATE U3045 ( .I1(n2072), .I2(n2073), .O(n5735) );
  NAND_GATE U3046 ( .I1(n2040), .I2(donnee[16]), .O(n2073) );
  NAND_GATE U3047 ( .I1(\registres[1][16] ), .I2(n2041), .O(n2072) );
  NAND_GATE U3048 ( .I1(n2074), .I2(n2075), .O(n5736) );
  NAND_GATE U3049 ( .I1(n2040), .I2(donnee[17]), .O(n2075) );
  NAND_GATE U3050 ( .I1(\registres[1][17] ), .I2(n2041), .O(n2074) );
  NAND_GATE U3051 ( .I1(n2076), .I2(n2077), .O(n5737) );
  NAND_GATE U3052 ( .I1(n2040), .I2(donnee[18]), .O(n2077) );
  NAND_GATE U3053 ( .I1(\registres[1][18] ), .I2(n2041), .O(n2076) );
  NAND_GATE U3054 ( .I1(n2078), .I2(n2079), .O(n5738) );
  NAND_GATE U3055 ( .I1(n2040), .I2(donnee[19]), .O(n2079) );
  NAND_GATE U3056 ( .I1(\registres[1][19] ), .I2(n2041), .O(n2078) );
  NAND_GATE U3057 ( .I1(n2080), .I2(n2081), .O(n5739) );
  NAND_GATE U3058 ( .I1(n2040), .I2(donnee[20]), .O(n2081) );
  NAND_GATE U3059 ( .I1(\registres[1][20] ), .I2(n2041), .O(n2080) );
  NAND_GATE U3060 ( .I1(n2082), .I2(n2083), .O(n5740) );
  NAND_GATE U3061 ( .I1(n2040), .I2(donnee[21]), .O(n2083) );
  NAND_GATE U3062 ( .I1(\registres[1][21] ), .I2(n2041), .O(n2082) );
  NAND_GATE U3063 ( .I1(n2084), .I2(n2085), .O(n5741) );
  NAND_GATE U3064 ( .I1(n2040), .I2(donnee[22]), .O(n2085) );
  NAND_GATE U3065 ( .I1(\registres[1][22] ), .I2(n2041), .O(n2084) );
  NAND_GATE U3066 ( .I1(n2086), .I2(n2087), .O(n5742) );
  NAND_GATE U3067 ( .I1(n2040), .I2(donnee[23]), .O(n2087) );
  NAND_GATE U3068 ( .I1(\registres[1][23] ), .I2(n2041), .O(n2086) );
  NAND_GATE U3069 ( .I1(n2088), .I2(n2089), .O(n5743) );
  NAND_GATE U3070 ( .I1(n2040), .I2(donnee[24]), .O(n2089) );
  NAND_GATE U3071 ( .I1(\registres[1][24] ), .I2(n2041), .O(n2088) );
  NAND_GATE U3072 ( .I1(n2090), .I2(n2091), .O(n5744) );
  NAND_GATE U3073 ( .I1(n2040), .I2(donnee[25]), .O(n2091) );
  NAND_GATE U3074 ( .I1(\registres[1][25] ), .I2(n2041), .O(n2090) );
  NAND_GATE U3075 ( .I1(n2092), .I2(n2093), .O(n5745) );
  NAND_GATE U3076 ( .I1(n2040), .I2(donnee[26]), .O(n2093) );
  NAND_GATE U3077 ( .I1(\registres[1][26] ), .I2(n2041), .O(n2092) );
  NAND_GATE U3078 ( .I1(n2094), .I2(n2095), .O(n5746) );
  NAND_GATE U3079 ( .I1(n2040), .I2(donnee[27]), .O(n2095) );
  NAND_GATE U3080 ( .I1(\registres[1][27] ), .I2(n2041), .O(n2094) );
  NAND_GATE U3081 ( .I1(n2096), .I2(n2097), .O(n5747) );
  NAND_GATE U3082 ( .I1(n2040), .I2(donnee[28]), .O(n2097) );
  NAND_GATE U3083 ( .I1(\registres[1][28] ), .I2(n2041), .O(n2096) );
  NAND_GATE U3084 ( .I1(n2098), .I2(n2099), .O(n5748) );
  NAND_GATE U3085 ( .I1(n2040), .I2(donnee[29]), .O(n2099) );
  NAND_GATE U3086 ( .I1(\registres[1][29] ), .I2(n2041), .O(n2098) );
  NAND_GATE U3087 ( .I1(n2100), .I2(n2101), .O(n5749) );
  NAND_GATE U3088 ( .I1(n2040), .I2(donnee[30]), .O(n2101) );
  NAND_GATE U3089 ( .I1(\registres[1][30] ), .I2(n2041), .O(n2100) );
  NAND_GATE U3090 ( .I1(n2102), .I2(n2103), .O(n5750) );
  NAND_GATE U3091 ( .I1(n2040), .I2(donnee[31]), .O(n2103) );
  AND_GATE U3092 ( .I1(n2104), .I2(n1), .O(n2040) );
  NAND_GATE U3093 ( .I1(\registres[1][31] ), .I2(n2041), .O(n2102) );
  NOR_GATE U3094 ( .I1(n2104), .I2(reset), .O(n2041) );
  AND3_GATE U3095 ( .I1(n492), .I2(cmd_ecr), .I3(n1702), .O(n2104) );
  NOR_GATE U3096 ( .I1(reg_dest[4]), .I2(reg_dest[3]), .O(n1702) );
  NOR3_GATE U3097 ( .I1(reg_dest[1]), .I2(reg_dest[2]), .I3(n4), .O(n492) );
  AND_GATE U3098 ( .I1(n2105), .I2(n2106), .O(data_src2[9]) );
  NAND4_GATE U3099 ( .I1(n2107), .I2(n2108), .I3(n2109), .I4(n2110), .O(n2106)
         );
  AND5_GATE U3100 ( .I1(n2111), .I2(n2112), .I3(n2113), .I4(n2114), .I5(n2115), 
        .O(n2110) );
  AND4_GATE U3101 ( .I1(n2116), .I2(n2117), .I3(n2118), .I4(n2119), .O(n2115)
         );
  NAND_GATE U3102 ( .I1(n2120), .I2(\registres[24][9] ), .O(n2119) );
  NAND_GATE U3103 ( .I1(n2121), .I2(\registres[25][9] ), .O(n2118) );
  NAND_GATE U3104 ( .I1(n2122), .I2(\registres[3][9] ), .O(n2117) );
  NAND_GATE U3105 ( .I1(n2123), .I2(\registres[26][9] ), .O(n2116) );
  NAND_GATE U3106 ( .I1(n2124), .I2(\registres[27][9] ), .O(n2114) );
  NAND_GATE U3107 ( .I1(n2125), .I2(\registres[10][9] ), .O(n2113) );
  NAND_GATE U3108 ( .I1(n2126), .I2(\registres[18][9] ), .O(n2112) );
  NAND_GATE U3109 ( .I1(n2127), .I2(\registres[5][9] ), .O(n2111) );
  AND5_GATE U3110 ( .I1(n2128), .I2(n2129), .I3(n2130), .I4(n2131), .I5(n2132), 
        .O(n2109) );
  AND4_GATE U3111 ( .I1(n2133), .I2(n2134), .I3(n2135), .I4(n2136), .O(n2132)
         );
  NAND_GATE U3112 ( .I1(n2137), .I2(\registres[28][9] ), .O(n2136) );
  NAND_GATE U3113 ( .I1(n2138), .I2(\registres[29][9] ), .O(n2135) );
  NAND_GATE U3114 ( .I1(n2139), .I2(\registres[12][9] ), .O(n2134) );
  NAND_GATE U3115 ( .I1(n2140), .I2(\registres[20][9] ), .O(n2133) );
  NAND_GATE U3116 ( .I1(n2141), .I2(\registres[1][9] ), .O(n2131) );
  NAND_GATE U3117 ( .I1(n2142), .I2(\registres[9][9] ), .O(n2130) );
  NAND_GATE U3118 ( .I1(n2143), .I2(\registres[11][9] ), .O(n2129) );
  NAND_GATE U3119 ( .I1(n2144), .I2(\registres[13][9] ), .O(n2128) );
  AND5_GATE U3120 ( .I1(n2145), .I2(n2146), .I3(n2147), .I4(n2148), .I5(n2149), 
        .O(n2108) );
  AND4_GATE U3121 ( .I1(n2150), .I2(n2151), .I3(n2152), .I4(n2153), .O(n2149)
         );
  NAND_GATE U3122 ( .I1(n2154), .I2(\registres[17][9] ), .O(n2153) );
  NAND_GATE U3123 ( .I1(n2155), .I2(\registres[19][9] ), .O(n2152) );
  NAND_GATE U3124 ( .I1(n2156), .I2(\registres[21][9] ), .O(n2151) );
  NAND_GATE U3125 ( .I1(n2157), .I2(\registres[6][9] ), .O(n2150) );
  NAND_GATE U3126 ( .I1(n2158), .I2(\registres[7][9] ), .O(n2148) );
  NAND_GATE U3127 ( .I1(n2159), .I2(\registres[30][9] ), .O(n2147) );
  NAND_GATE U3128 ( .I1(n2160), .I2(\registres[31][9] ), .O(n2146) );
  NAND_GATE U3129 ( .I1(n2161), .I2(\registres[14][9] ), .O(n2145) );
  AND4_GATE U3130 ( .I1(n2162), .I2(n2163), .I3(n2164), .I4(n2165), .O(n2107)
         );
  AND4_GATE U3131 ( .I1(n2166), .I2(n2167), .I3(n2168), .I4(n2169), .O(n2165)
         );
  NAND_GATE U3132 ( .I1(n2170), .I2(\registres[22][9] ), .O(n2169) );
  NAND_GATE U3133 ( .I1(n2171), .I2(\registres[15][9] ), .O(n2168) );
  NAND_GATE U3134 ( .I1(n2172), .I2(\registres[23][9] ), .O(n2167) );
  NAND_GATE U3135 ( .I1(n2173), .I2(\registres[4][9] ), .O(n2166) );
  NAND_GATE U3136 ( .I1(n2174), .I2(\registres[8][9] ), .O(n2164) );
  NAND_GATE U3137 ( .I1(n2175), .I2(\registres[2][9] ), .O(n2163) );
  NAND_GATE U3138 ( .I1(n2176), .I2(\registres[16][9] ), .O(n2162) );
  AND_GATE U3139 ( .I1(n2177), .I2(n2105), .O(data_src2[8]) );
  NAND4_GATE U3140 ( .I1(n2178), .I2(n2179), .I3(n2180), .I4(n2181), .O(n2177)
         );
  AND5_GATE U3141 ( .I1(n2182), .I2(n2183), .I3(n2184), .I4(n2185), .I5(n2186), 
        .O(n2181) );
  AND4_GATE U3142 ( .I1(n2187), .I2(n2188), .I3(n2189), .I4(n2190), .O(n2186)
         );
  NAND_GATE U3143 ( .I1(n2120), .I2(\registres[24][8] ), .O(n2190) );
  NAND_GATE U3144 ( .I1(n2121), .I2(\registres[25][8] ), .O(n2189) );
  NAND_GATE U3145 ( .I1(n2122), .I2(\registres[3][8] ), .O(n2188) );
  NAND_GATE U3146 ( .I1(n2123), .I2(\registres[26][8] ), .O(n2187) );
  NAND_GATE U3147 ( .I1(n2124), .I2(\registres[27][8] ), .O(n2185) );
  NAND_GATE U3148 ( .I1(n2125), .I2(\registres[10][8] ), .O(n2184) );
  NAND_GATE U3149 ( .I1(n2126), .I2(\registres[18][8] ), .O(n2183) );
  NAND_GATE U3150 ( .I1(n2127), .I2(\registres[5][8] ), .O(n2182) );
  AND5_GATE U3151 ( .I1(n2191), .I2(n2192), .I3(n2193), .I4(n2194), .I5(n2195), 
        .O(n2180) );
  AND4_GATE U3152 ( .I1(n2196), .I2(n2197), .I3(n2198), .I4(n2199), .O(n2195)
         );
  NAND_GATE U3153 ( .I1(n2137), .I2(\registres[28][8] ), .O(n2199) );
  NAND_GATE U3154 ( .I1(n2138), .I2(\registres[29][8] ), .O(n2198) );
  NAND_GATE U3155 ( .I1(n2139), .I2(\registres[12][8] ), .O(n2197) );
  NAND_GATE U3156 ( .I1(n2140), .I2(\registres[20][8] ), .O(n2196) );
  NAND_GATE U3157 ( .I1(n2141), .I2(\registres[1][8] ), .O(n2194) );
  NAND_GATE U3158 ( .I1(n2142), .I2(\registres[9][8] ), .O(n2193) );
  NAND_GATE U3159 ( .I1(n2143), .I2(\registres[11][8] ), .O(n2192) );
  NAND_GATE U3160 ( .I1(n2144), .I2(\registres[13][8] ), .O(n2191) );
  AND5_GATE U3161 ( .I1(n2200), .I2(n2201), .I3(n2202), .I4(n2203), .I5(n2204), 
        .O(n2179) );
  AND4_GATE U3162 ( .I1(n2205), .I2(n2206), .I3(n2207), .I4(n2208), .O(n2204)
         );
  NAND_GATE U3163 ( .I1(n2154), .I2(\registres[17][8] ), .O(n2208) );
  NAND_GATE U3164 ( .I1(n2155), .I2(\registres[19][8] ), .O(n2207) );
  NAND_GATE U3165 ( .I1(n2156), .I2(\registres[21][8] ), .O(n2206) );
  NAND_GATE U3166 ( .I1(n2157), .I2(\registres[6][8] ), .O(n2205) );
  NAND_GATE U3167 ( .I1(n2158), .I2(\registres[7][8] ), .O(n2203) );
  NAND_GATE U3168 ( .I1(n2159), .I2(\registres[30][8] ), .O(n2202) );
  NAND_GATE U3169 ( .I1(n2160), .I2(\registres[31][8] ), .O(n2201) );
  NAND_GATE U3170 ( .I1(n2161), .I2(\registres[14][8] ), .O(n2200) );
  AND4_GATE U3171 ( .I1(n2209), .I2(n2210), .I3(n2211), .I4(n2212), .O(n2178)
         );
  AND4_GATE U3172 ( .I1(n2213), .I2(n2214), .I3(n2215), .I4(n2216), .O(n2212)
         );
  NAND_GATE U3173 ( .I1(n2170), .I2(\registres[22][8] ), .O(n2216) );
  NAND_GATE U3174 ( .I1(n2171), .I2(\registres[15][8] ), .O(n2215) );
  NAND_GATE U3175 ( .I1(n2172), .I2(\registres[23][8] ), .O(n2214) );
  NAND_GATE U3176 ( .I1(n2173), .I2(\registres[4][8] ), .O(n2213) );
  NAND_GATE U3177 ( .I1(n2174), .I2(\registres[8][8] ), .O(n2211) );
  NAND_GATE U3178 ( .I1(n2175), .I2(\registres[2][8] ), .O(n2210) );
  NAND_GATE U3179 ( .I1(n2176), .I2(\registres[16][8] ), .O(n2209) );
  AND_GATE U3180 ( .I1(n2217), .I2(n2105), .O(data_src2[7]) );
  NAND4_GATE U3181 ( .I1(n2218), .I2(n2219), .I3(n2220), .I4(n2221), .O(n2217)
         );
  AND5_GATE U3182 ( .I1(n2222), .I2(n2223), .I3(n2224), .I4(n2225), .I5(n2226), 
        .O(n2221) );
  AND4_GATE U3183 ( .I1(n2227), .I2(n2228), .I3(n2229), .I4(n2230), .O(n2226)
         );
  NAND_GATE U3184 ( .I1(n2120), .I2(\registres[24][7] ), .O(n2230) );
  NAND_GATE U3185 ( .I1(n2121), .I2(\registres[25][7] ), .O(n2229) );
  NAND_GATE U3186 ( .I1(n2122), .I2(\registres[3][7] ), .O(n2228) );
  NAND_GATE U3187 ( .I1(n2123), .I2(\registres[26][7] ), .O(n2227) );
  NAND_GATE U3188 ( .I1(n2124), .I2(\registres[27][7] ), .O(n2225) );
  NAND_GATE U3189 ( .I1(n2125), .I2(\registres[10][7] ), .O(n2224) );
  NAND_GATE U3190 ( .I1(n2126), .I2(\registres[18][7] ), .O(n2223) );
  NAND_GATE U3191 ( .I1(n2127), .I2(\registres[5][7] ), .O(n2222) );
  AND5_GATE U3192 ( .I1(n2231), .I2(n2232), .I3(n2233), .I4(n2234), .I5(n2235), 
        .O(n2220) );
  AND4_GATE U3193 ( .I1(n2236), .I2(n2237), .I3(n2238), .I4(n2239), .O(n2235)
         );
  NAND_GATE U3194 ( .I1(n2137), .I2(\registres[28][7] ), .O(n2239) );
  NAND_GATE U3195 ( .I1(n2138), .I2(\registres[29][7] ), .O(n2238) );
  NAND_GATE U3196 ( .I1(n2139), .I2(\registres[12][7] ), .O(n2237) );
  NAND_GATE U3197 ( .I1(n2140), .I2(\registres[20][7] ), .O(n2236) );
  NAND_GATE U3198 ( .I1(n2141), .I2(\registres[1][7] ), .O(n2234) );
  NAND_GATE U3199 ( .I1(n2142), .I2(\registres[9][7] ), .O(n2233) );
  NAND_GATE U3200 ( .I1(n2143), .I2(\registres[11][7] ), .O(n2232) );
  NAND_GATE U3201 ( .I1(n2144), .I2(\registres[13][7] ), .O(n2231) );
  AND5_GATE U3202 ( .I1(n2240), .I2(n2241), .I3(n2242), .I4(n2243), .I5(n2244), 
        .O(n2219) );
  AND4_GATE U3203 ( .I1(n2245), .I2(n2246), .I3(n2247), .I4(n2248), .O(n2244)
         );
  NAND_GATE U3204 ( .I1(n2154), .I2(\registres[17][7] ), .O(n2248) );
  NAND_GATE U3205 ( .I1(n2155), .I2(\registres[19][7] ), .O(n2247) );
  NAND_GATE U3206 ( .I1(n2156), .I2(\registres[21][7] ), .O(n2246) );
  NAND_GATE U3207 ( .I1(n2157), .I2(\registres[6][7] ), .O(n2245) );
  NAND_GATE U3208 ( .I1(n2158), .I2(\registres[7][7] ), .O(n2243) );
  NAND_GATE U3209 ( .I1(n2159), .I2(\registres[30][7] ), .O(n2242) );
  NAND_GATE U3210 ( .I1(n2160), .I2(\registres[31][7] ), .O(n2241) );
  NAND_GATE U3211 ( .I1(n2161), .I2(\registres[14][7] ), .O(n2240) );
  AND4_GATE U3212 ( .I1(n2249), .I2(n2250), .I3(n2251), .I4(n2252), .O(n2218)
         );
  AND4_GATE U3213 ( .I1(n2253), .I2(n2254), .I3(n2255), .I4(n2256), .O(n2252)
         );
  NAND_GATE U3214 ( .I1(n2170), .I2(\registres[22][7] ), .O(n2256) );
  NAND_GATE U3215 ( .I1(n2171), .I2(\registres[15][7] ), .O(n2255) );
  NAND_GATE U3216 ( .I1(n2172), .I2(\registres[23][7] ), .O(n2254) );
  NAND_GATE U3217 ( .I1(n2173), .I2(\registres[4][7] ), .O(n2253) );
  NAND_GATE U3218 ( .I1(n2174), .I2(\registres[8][7] ), .O(n2251) );
  NAND_GATE U3219 ( .I1(n2175), .I2(\registres[2][7] ), .O(n2250) );
  NAND_GATE U3220 ( .I1(n2176), .I2(\registres[16][7] ), .O(n2249) );
  AND_GATE U3221 ( .I1(n2257), .I2(n2105), .O(data_src2[6]) );
  NAND4_GATE U3222 ( .I1(n2258), .I2(n2259), .I3(n2260), .I4(n2261), .O(n2257)
         );
  AND5_GATE U3223 ( .I1(n2262), .I2(n2263), .I3(n2264), .I4(n2265), .I5(n2266), 
        .O(n2261) );
  AND4_GATE U3224 ( .I1(n2267), .I2(n2268), .I3(n2269), .I4(n2270), .O(n2266)
         );
  NAND_GATE U3225 ( .I1(n2120), .I2(\registres[24][6] ), .O(n2270) );
  NAND_GATE U3226 ( .I1(n2121), .I2(\registres[25][6] ), .O(n2269) );
  NAND_GATE U3227 ( .I1(n2122), .I2(\registres[3][6] ), .O(n2268) );
  NAND_GATE U3228 ( .I1(n2123), .I2(\registres[26][6] ), .O(n2267) );
  NAND_GATE U3229 ( .I1(n2124), .I2(\registres[27][6] ), .O(n2265) );
  NAND_GATE U3230 ( .I1(n2125), .I2(\registres[10][6] ), .O(n2264) );
  NAND_GATE U3231 ( .I1(n2126), .I2(\registres[18][6] ), .O(n2263) );
  NAND_GATE U3232 ( .I1(n2127), .I2(\registres[5][6] ), .O(n2262) );
  AND5_GATE U3233 ( .I1(n2271), .I2(n2272), .I3(n2273), .I4(n2274), .I5(n2275), 
        .O(n2260) );
  AND4_GATE U3234 ( .I1(n2276), .I2(n2277), .I3(n2278), .I4(n2279), .O(n2275)
         );
  NAND_GATE U3235 ( .I1(n2137), .I2(\registres[28][6] ), .O(n2279) );
  NAND_GATE U3236 ( .I1(n2138), .I2(\registres[29][6] ), .O(n2278) );
  NAND_GATE U3237 ( .I1(n2139), .I2(\registres[12][6] ), .O(n2277) );
  NAND_GATE U3238 ( .I1(n2140), .I2(\registres[20][6] ), .O(n2276) );
  NAND_GATE U3239 ( .I1(n2141), .I2(\registres[1][6] ), .O(n2274) );
  NAND_GATE U3240 ( .I1(n2142), .I2(\registres[9][6] ), .O(n2273) );
  NAND_GATE U3241 ( .I1(n2143), .I2(\registres[11][6] ), .O(n2272) );
  NAND_GATE U3242 ( .I1(n2144), .I2(\registres[13][6] ), .O(n2271) );
  AND5_GATE U3243 ( .I1(n2280), .I2(n2281), .I3(n2282), .I4(n2283), .I5(n2284), 
        .O(n2259) );
  AND4_GATE U3244 ( .I1(n2285), .I2(n2286), .I3(n2287), .I4(n2288), .O(n2284)
         );
  NAND_GATE U3245 ( .I1(n2154), .I2(\registres[17][6] ), .O(n2288) );
  NAND_GATE U3246 ( .I1(n2155), .I2(\registres[19][6] ), .O(n2287) );
  NAND_GATE U3247 ( .I1(n2156), .I2(\registres[21][6] ), .O(n2286) );
  NAND_GATE U3248 ( .I1(n2157), .I2(\registres[6][6] ), .O(n2285) );
  NAND_GATE U3249 ( .I1(n2158), .I2(\registres[7][6] ), .O(n2283) );
  NAND_GATE U3250 ( .I1(n2159), .I2(\registres[30][6] ), .O(n2282) );
  NAND_GATE U3251 ( .I1(n2160), .I2(\registres[31][6] ), .O(n2281) );
  NAND_GATE U3252 ( .I1(n2161), .I2(\registres[14][6] ), .O(n2280) );
  AND4_GATE U3253 ( .I1(n2289), .I2(n2290), .I3(n2291), .I4(n2292), .O(n2258)
         );
  AND4_GATE U3254 ( .I1(n2293), .I2(n2294), .I3(n2295), .I4(n2296), .O(n2292)
         );
  NAND_GATE U3255 ( .I1(n2170), .I2(\registres[22][6] ), .O(n2296) );
  NAND_GATE U3256 ( .I1(n2171), .I2(\registres[15][6] ), .O(n2295) );
  NAND_GATE U3257 ( .I1(n2172), .I2(\registres[23][6] ), .O(n2294) );
  NAND_GATE U3258 ( .I1(n2173), .I2(\registres[4][6] ), .O(n2293) );
  NAND_GATE U3259 ( .I1(n2174), .I2(\registres[8][6] ), .O(n2291) );
  NAND_GATE U3260 ( .I1(n2175), .I2(\registres[2][6] ), .O(n2290) );
  NAND_GATE U3261 ( .I1(n2176), .I2(\registres[16][6] ), .O(n2289) );
  AND_GATE U3262 ( .I1(n2297), .I2(n2105), .O(data_src2[5]) );
  NAND4_GATE U3263 ( .I1(n2298), .I2(n2299), .I3(n2300), .I4(n2301), .O(n2297)
         );
  AND5_GATE U3264 ( .I1(n2302), .I2(n2303), .I3(n2304), .I4(n2305), .I5(n2306), 
        .O(n2301) );
  AND4_GATE U3265 ( .I1(n2307), .I2(n2308), .I3(n2309), .I4(n2310), .O(n2306)
         );
  NAND_GATE U3266 ( .I1(n2120), .I2(\registres[24][5] ), .O(n2310) );
  NAND_GATE U3267 ( .I1(n2121), .I2(\registres[25][5] ), .O(n2309) );
  NAND_GATE U3268 ( .I1(n2122), .I2(\registres[3][5] ), .O(n2308) );
  NAND_GATE U3269 ( .I1(n2123), .I2(\registres[26][5] ), .O(n2307) );
  NAND_GATE U3270 ( .I1(n2124), .I2(\registres[27][5] ), .O(n2305) );
  NAND_GATE U3271 ( .I1(n2125), .I2(\registres[10][5] ), .O(n2304) );
  NAND_GATE U3272 ( .I1(n2126), .I2(\registres[18][5] ), .O(n2303) );
  NAND_GATE U3273 ( .I1(n2127), .I2(\registres[5][5] ), .O(n2302) );
  AND5_GATE U3274 ( .I1(n2311), .I2(n2312), .I3(n2313), .I4(n2314), .I5(n2315), 
        .O(n2300) );
  AND4_GATE U3275 ( .I1(n2316), .I2(n2317), .I3(n2318), .I4(n2319), .O(n2315)
         );
  NAND_GATE U3276 ( .I1(n2137), .I2(\registres[28][5] ), .O(n2319) );
  NAND_GATE U3277 ( .I1(n2138), .I2(\registres[29][5] ), .O(n2318) );
  NAND_GATE U3278 ( .I1(n2139), .I2(\registres[12][5] ), .O(n2317) );
  NAND_GATE U3279 ( .I1(n2140), .I2(\registres[20][5] ), .O(n2316) );
  NAND_GATE U3280 ( .I1(n2141), .I2(\registres[1][5] ), .O(n2314) );
  NAND_GATE U3281 ( .I1(n2142), .I2(\registres[9][5] ), .O(n2313) );
  NAND_GATE U3282 ( .I1(n2143), .I2(\registres[11][5] ), .O(n2312) );
  NAND_GATE U3283 ( .I1(n2144), .I2(\registres[13][5] ), .O(n2311) );
  AND5_GATE U3284 ( .I1(n2320), .I2(n2321), .I3(n2322), .I4(n2323), .I5(n2324), 
        .O(n2299) );
  AND4_GATE U3285 ( .I1(n2325), .I2(n2326), .I3(n2327), .I4(n2328), .O(n2324)
         );
  NAND_GATE U3286 ( .I1(n2154), .I2(\registres[17][5] ), .O(n2328) );
  NAND_GATE U3287 ( .I1(n2155), .I2(\registres[19][5] ), .O(n2327) );
  NAND_GATE U3288 ( .I1(n2156), .I2(\registres[21][5] ), .O(n2326) );
  NAND_GATE U3289 ( .I1(n2157), .I2(\registres[6][5] ), .O(n2325) );
  NAND_GATE U3290 ( .I1(n2158), .I2(\registres[7][5] ), .O(n2323) );
  NAND_GATE U3291 ( .I1(n2159), .I2(\registres[30][5] ), .O(n2322) );
  NAND_GATE U3292 ( .I1(n2160), .I2(\registres[31][5] ), .O(n2321) );
  NAND_GATE U3293 ( .I1(n2161), .I2(\registres[14][5] ), .O(n2320) );
  AND4_GATE U3294 ( .I1(n2329), .I2(n2330), .I3(n2331), .I4(n2332), .O(n2298)
         );
  AND4_GATE U3295 ( .I1(n2333), .I2(n2334), .I3(n2335), .I4(n2336), .O(n2332)
         );
  NAND_GATE U3296 ( .I1(n2170), .I2(\registres[22][5] ), .O(n2336) );
  NAND_GATE U3297 ( .I1(n2171), .I2(\registres[15][5] ), .O(n2335) );
  NAND_GATE U3298 ( .I1(n2172), .I2(\registres[23][5] ), .O(n2334) );
  NAND_GATE U3299 ( .I1(n2173), .I2(\registres[4][5] ), .O(n2333) );
  NAND_GATE U3300 ( .I1(n2174), .I2(\registres[8][5] ), .O(n2331) );
  NAND_GATE U3301 ( .I1(n2175), .I2(\registres[2][5] ), .O(n2330) );
  NAND_GATE U3302 ( .I1(n2176), .I2(\registres[16][5] ), .O(n2329) );
  AND_GATE U3303 ( .I1(n2337), .I2(n2105), .O(data_src2[4]) );
  NAND4_GATE U3304 ( .I1(n2338), .I2(n2339), .I3(n2340), .I4(n2341), .O(n2337)
         );
  AND5_GATE U3305 ( .I1(n2342), .I2(n2343), .I3(n2344), .I4(n2345), .I5(n2346), 
        .O(n2341) );
  AND4_GATE U3306 ( .I1(n2347), .I2(n2348), .I3(n2349), .I4(n2350), .O(n2346)
         );
  NAND_GATE U3307 ( .I1(n2120), .I2(\registres[24][4] ), .O(n2350) );
  NAND_GATE U3308 ( .I1(n2121), .I2(\registres[25][4] ), .O(n2349) );
  NAND_GATE U3309 ( .I1(n2122), .I2(\registres[3][4] ), .O(n2348) );
  NAND_GATE U3310 ( .I1(n2123), .I2(\registres[26][4] ), .O(n2347) );
  NAND_GATE U3311 ( .I1(n2124), .I2(\registres[27][4] ), .O(n2345) );
  NAND_GATE U3312 ( .I1(n2125), .I2(\registres[10][4] ), .O(n2344) );
  NAND_GATE U3313 ( .I1(n2126), .I2(\registres[18][4] ), .O(n2343) );
  NAND_GATE U3314 ( .I1(n2127), .I2(\registres[5][4] ), .O(n2342) );
  AND5_GATE U3315 ( .I1(n2351), .I2(n2352), .I3(n2353), .I4(n2354), .I5(n2355), 
        .O(n2340) );
  AND4_GATE U3316 ( .I1(n2356), .I2(n2357), .I3(n2358), .I4(n2359), .O(n2355)
         );
  NAND_GATE U3317 ( .I1(n2137), .I2(\registres[28][4] ), .O(n2359) );
  NAND_GATE U3318 ( .I1(n2138), .I2(\registres[29][4] ), .O(n2358) );
  NAND_GATE U3319 ( .I1(n2139), .I2(\registres[12][4] ), .O(n2357) );
  NAND_GATE U3320 ( .I1(n2140), .I2(\registres[20][4] ), .O(n2356) );
  NAND_GATE U3321 ( .I1(n2141), .I2(\registres[1][4] ), .O(n2354) );
  NAND_GATE U3322 ( .I1(n2142), .I2(\registres[9][4] ), .O(n2353) );
  NAND_GATE U3323 ( .I1(n2143), .I2(\registres[11][4] ), .O(n2352) );
  NAND_GATE U3324 ( .I1(n2144), .I2(\registres[13][4] ), .O(n2351) );
  AND5_GATE U3325 ( .I1(n2360), .I2(n2361), .I3(n2362), .I4(n2363), .I5(n2364), 
        .O(n2339) );
  AND4_GATE U3326 ( .I1(n2365), .I2(n2366), .I3(n2367), .I4(n2368), .O(n2364)
         );
  NAND_GATE U3327 ( .I1(n2154), .I2(\registres[17][4] ), .O(n2368) );
  NAND_GATE U3328 ( .I1(n2155), .I2(\registres[19][4] ), .O(n2367) );
  NAND_GATE U3329 ( .I1(n2156), .I2(\registres[21][4] ), .O(n2366) );
  NAND_GATE U3330 ( .I1(n2157), .I2(\registres[6][4] ), .O(n2365) );
  NAND_GATE U3331 ( .I1(n2158), .I2(\registres[7][4] ), .O(n2363) );
  NAND_GATE U3332 ( .I1(n2159), .I2(\registres[30][4] ), .O(n2362) );
  NAND_GATE U3333 ( .I1(n2160), .I2(\registres[31][4] ), .O(n2361) );
  NAND_GATE U3334 ( .I1(n2161), .I2(\registres[14][4] ), .O(n2360) );
  AND4_GATE U3335 ( .I1(n2369), .I2(n2370), .I3(n2371), .I4(n2372), .O(n2338)
         );
  AND4_GATE U3336 ( .I1(n2373), .I2(n2374), .I3(n2375), .I4(n2376), .O(n2372)
         );
  NAND_GATE U3337 ( .I1(n2170), .I2(\registres[22][4] ), .O(n2376) );
  NAND_GATE U3338 ( .I1(n2171), .I2(\registres[15][4] ), .O(n2375) );
  NAND_GATE U3339 ( .I1(n2172), .I2(\registres[23][4] ), .O(n2374) );
  NAND_GATE U3340 ( .I1(n2173), .I2(\registres[4][4] ), .O(n2373) );
  NAND_GATE U3341 ( .I1(n2174), .I2(\registres[8][4] ), .O(n2371) );
  NAND_GATE U3342 ( .I1(n2175), .I2(\registres[2][4] ), .O(n2370) );
  NAND_GATE U3343 ( .I1(n2176), .I2(\registres[16][4] ), .O(n2369) );
  AND_GATE U3344 ( .I1(n2377), .I2(n2105), .O(data_src2[3]) );
  NAND4_GATE U3345 ( .I1(n2378), .I2(n2379), .I3(n2380), .I4(n2381), .O(n2377)
         );
  AND5_GATE U3346 ( .I1(n2382), .I2(n2383), .I3(n2384), .I4(n2385), .I5(n2386), 
        .O(n2381) );
  AND4_GATE U3347 ( .I1(n2387), .I2(n2388), .I3(n2389), .I4(n2390), .O(n2386)
         );
  NAND_GATE U3348 ( .I1(n2120), .I2(\registres[24][3] ), .O(n2390) );
  NAND_GATE U3349 ( .I1(n2121), .I2(\registres[25][3] ), .O(n2389) );
  NAND_GATE U3350 ( .I1(n2122), .I2(\registres[3][3] ), .O(n2388) );
  NAND_GATE U3351 ( .I1(n2123), .I2(\registres[26][3] ), .O(n2387) );
  NAND_GATE U3352 ( .I1(n2124), .I2(\registres[27][3] ), .O(n2385) );
  NAND_GATE U3353 ( .I1(n2125), .I2(\registres[10][3] ), .O(n2384) );
  NAND_GATE U3354 ( .I1(n2126), .I2(\registres[18][3] ), .O(n2383) );
  NAND_GATE U3355 ( .I1(n2127), .I2(\registres[5][3] ), .O(n2382) );
  AND5_GATE U3356 ( .I1(n2391), .I2(n2392), .I3(n2393), .I4(n2394), .I5(n2395), 
        .O(n2380) );
  AND4_GATE U3357 ( .I1(n2396), .I2(n2397), .I3(n2398), .I4(n2399), .O(n2395)
         );
  NAND_GATE U3358 ( .I1(n2137), .I2(\registres[28][3] ), .O(n2399) );
  NAND_GATE U3359 ( .I1(n2138), .I2(\registres[29][3] ), .O(n2398) );
  NAND_GATE U3360 ( .I1(n2139), .I2(\registres[12][3] ), .O(n2397) );
  NAND_GATE U3361 ( .I1(n2140), .I2(\registres[20][3] ), .O(n2396) );
  NAND_GATE U3362 ( .I1(n2141), .I2(\registres[1][3] ), .O(n2394) );
  NAND_GATE U3363 ( .I1(n2142), .I2(\registres[9][3] ), .O(n2393) );
  NAND_GATE U3364 ( .I1(n2143), .I2(\registres[11][3] ), .O(n2392) );
  NAND_GATE U3365 ( .I1(n2144), .I2(\registres[13][3] ), .O(n2391) );
  AND5_GATE U3366 ( .I1(n2400), .I2(n2401), .I3(n2402), .I4(n2403), .I5(n2404), 
        .O(n2379) );
  AND4_GATE U3367 ( .I1(n2405), .I2(n2406), .I3(n2407), .I4(n2408), .O(n2404)
         );
  NAND_GATE U3368 ( .I1(n2154), .I2(\registres[17][3] ), .O(n2408) );
  NAND_GATE U3369 ( .I1(n2155), .I2(\registres[19][3] ), .O(n2407) );
  NAND_GATE U3370 ( .I1(n2156), .I2(\registres[21][3] ), .O(n2406) );
  NAND_GATE U3371 ( .I1(n2157), .I2(\registres[6][3] ), .O(n2405) );
  NAND_GATE U3372 ( .I1(n2158), .I2(\registres[7][3] ), .O(n2403) );
  NAND_GATE U3373 ( .I1(n2159), .I2(\registres[30][3] ), .O(n2402) );
  NAND_GATE U3374 ( .I1(n2160), .I2(\registres[31][3] ), .O(n2401) );
  NAND_GATE U3375 ( .I1(n2161), .I2(\registres[14][3] ), .O(n2400) );
  AND4_GATE U3376 ( .I1(n2409), .I2(n2410), .I3(n2411), .I4(n2412), .O(n2378)
         );
  AND4_GATE U3377 ( .I1(n2413), .I2(n2414), .I3(n2415), .I4(n2416), .O(n2412)
         );
  NAND_GATE U3378 ( .I1(n2170), .I2(\registres[22][3] ), .O(n2416) );
  NAND_GATE U3379 ( .I1(n2171), .I2(\registres[15][3] ), .O(n2415) );
  NAND_GATE U3380 ( .I1(n2172), .I2(\registres[23][3] ), .O(n2414) );
  NAND_GATE U3381 ( .I1(n2173), .I2(\registres[4][3] ), .O(n2413) );
  NAND_GATE U3382 ( .I1(n2174), .I2(\registres[8][3] ), .O(n2411) );
  NAND_GATE U3383 ( .I1(n2175), .I2(\registres[2][3] ), .O(n2410) );
  NAND_GATE U3384 ( .I1(n2176), .I2(\registres[16][3] ), .O(n2409) );
  AND_GATE U3385 ( .I1(n2417), .I2(n2105), .O(data_src2[31]) );
  NAND4_GATE U3386 ( .I1(n2418), .I2(n2419), .I3(n2420), .I4(n2421), .O(n2417)
         );
  AND5_GATE U3387 ( .I1(n2422), .I2(n2423), .I3(n2424), .I4(n2425), .I5(n2426), 
        .O(n2421) );
  AND4_GATE U3388 ( .I1(n2427), .I2(n2428), .I3(n2429), .I4(n2430), .O(n2426)
         );
  NAND_GATE U3389 ( .I1(n2120), .I2(\registres[24][31] ), .O(n2430) );
  NAND_GATE U3390 ( .I1(n2121), .I2(\registres[25][31] ), .O(n2429) );
  NAND_GATE U3391 ( .I1(n2122), .I2(\registres[3][31] ), .O(n2428) );
  NAND_GATE U3392 ( .I1(n2123), .I2(\registres[26][31] ), .O(n2427) );
  NAND_GATE U3393 ( .I1(n2124), .I2(\registres[27][31] ), .O(n2425) );
  NAND_GATE U3394 ( .I1(n2125), .I2(\registres[10][31] ), .O(n2424) );
  NAND_GATE U3395 ( .I1(n2126), .I2(\registres[18][31] ), .O(n2423) );
  NAND_GATE U3396 ( .I1(n2127), .I2(\registres[5][31] ), .O(n2422) );
  AND5_GATE U3397 ( .I1(n2431), .I2(n2432), .I3(n2433), .I4(n2434), .I5(n2435), 
        .O(n2420) );
  AND4_GATE U3398 ( .I1(n2436), .I2(n2437), .I3(n2438), .I4(n2439), .O(n2435)
         );
  NAND_GATE U3399 ( .I1(n2137), .I2(\registres[28][31] ), .O(n2439) );
  NAND_GATE U3400 ( .I1(n2138), .I2(\registres[29][31] ), .O(n2438) );
  NAND_GATE U3401 ( .I1(n2139), .I2(\registres[12][31] ), .O(n2437) );
  NAND_GATE U3402 ( .I1(n2140), .I2(\registres[20][31] ), .O(n2436) );
  NAND_GATE U3403 ( .I1(n2141), .I2(\registres[1][31] ), .O(n2434) );
  NAND_GATE U3404 ( .I1(n2142), .I2(\registres[9][31] ), .O(n2433) );
  NAND_GATE U3405 ( .I1(n2143), .I2(\registres[11][31] ), .O(n2432) );
  NAND_GATE U3406 ( .I1(n2144), .I2(\registres[13][31] ), .O(n2431) );
  AND5_GATE U3407 ( .I1(n2440), .I2(n2441), .I3(n2442), .I4(n2443), .I5(n2444), 
        .O(n2419) );
  AND4_GATE U3408 ( .I1(n2445), .I2(n2446), .I3(n2447), .I4(n2448), .O(n2444)
         );
  NAND_GATE U3409 ( .I1(n2154), .I2(\registres[17][31] ), .O(n2448) );
  NAND_GATE U3410 ( .I1(n2155), .I2(\registres[19][31] ), .O(n2447) );
  NAND_GATE U3411 ( .I1(n2156), .I2(\registres[21][31] ), .O(n2446) );
  NAND_GATE U3412 ( .I1(n2157), .I2(\registres[6][31] ), .O(n2445) );
  NAND_GATE U3413 ( .I1(n2158), .I2(\registres[7][31] ), .O(n2443) );
  NAND_GATE U3414 ( .I1(n2159), .I2(\registres[30][31] ), .O(n2442) );
  NAND_GATE U3415 ( .I1(n2160), .I2(\registres[31][31] ), .O(n2441) );
  NAND_GATE U3416 ( .I1(n2161), .I2(\registres[14][31] ), .O(n2440) );
  AND4_GATE U3417 ( .I1(n2449), .I2(n2450), .I3(n2451), .I4(n2452), .O(n2418)
         );
  AND4_GATE U3418 ( .I1(n2453), .I2(n2454), .I3(n2455), .I4(n2456), .O(n2452)
         );
  NAND_GATE U3419 ( .I1(n2170), .I2(\registres[22][31] ), .O(n2456) );
  NAND_GATE U3420 ( .I1(n2171), .I2(\registres[15][31] ), .O(n2455) );
  NAND_GATE U3421 ( .I1(n2172), .I2(\registres[23][31] ), .O(n2454) );
  NAND_GATE U3422 ( .I1(n2173), .I2(\registres[4][31] ), .O(n2453) );
  NAND_GATE U3423 ( .I1(n2174), .I2(\registres[8][31] ), .O(n2451) );
  NAND_GATE U3424 ( .I1(n2175), .I2(\registres[2][31] ), .O(n2450) );
  NAND_GATE U3425 ( .I1(n2176), .I2(\registres[16][31] ), .O(n2449) );
  AND_GATE U3426 ( .I1(n2457), .I2(n2105), .O(data_src2[30]) );
  NAND4_GATE U3427 ( .I1(n2458), .I2(n2459), .I3(n2460), .I4(n2461), .O(n2457)
         );
  AND5_GATE U3428 ( .I1(n2462), .I2(n2463), .I3(n2464), .I4(n2465), .I5(n2466), 
        .O(n2461) );
  AND4_GATE U3429 ( .I1(n2467), .I2(n2468), .I3(n2469), .I4(n2470), .O(n2466)
         );
  NAND_GATE U3430 ( .I1(n2120), .I2(\registres[24][30] ), .O(n2470) );
  NAND_GATE U3431 ( .I1(n2121), .I2(\registres[25][30] ), .O(n2469) );
  NAND_GATE U3432 ( .I1(n2122), .I2(\registres[3][30] ), .O(n2468) );
  NAND_GATE U3433 ( .I1(n2123), .I2(\registres[26][30] ), .O(n2467) );
  NAND_GATE U3434 ( .I1(n2124), .I2(\registres[27][30] ), .O(n2465) );
  NAND_GATE U3435 ( .I1(n2125), .I2(\registres[10][30] ), .O(n2464) );
  NAND_GATE U3436 ( .I1(n2126), .I2(\registres[18][30] ), .O(n2463) );
  NAND_GATE U3437 ( .I1(n2127), .I2(\registres[5][30] ), .O(n2462) );
  AND5_GATE U3438 ( .I1(n2471), .I2(n2472), .I3(n2473), .I4(n2474), .I5(n2475), 
        .O(n2460) );
  AND4_GATE U3439 ( .I1(n2476), .I2(n2477), .I3(n2478), .I4(n2479), .O(n2475)
         );
  NAND_GATE U3440 ( .I1(n2137), .I2(\registres[28][30] ), .O(n2479) );
  NAND_GATE U3441 ( .I1(n2138), .I2(\registres[29][30] ), .O(n2478) );
  NAND_GATE U3442 ( .I1(n2139), .I2(\registres[12][30] ), .O(n2477) );
  NAND_GATE U3443 ( .I1(n2140), .I2(\registres[20][30] ), .O(n2476) );
  NAND_GATE U3444 ( .I1(n2141), .I2(\registres[1][30] ), .O(n2474) );
  NAND_GATE U3445 ( .I1(n2142), .I2(\registres[9][30] ), .O(n2473) );
  NAND_GATE U3446 ( .I1(n2143), .I2(\registres[11][30] ), .O(n2472) );
  NAND_GATE U3447 ( .I1(n2144), .I2(\registres[13][30] ), .O(n2471) );
  AND5_GATE U3448 ( .I1(n2480), .I2(n2481), .I3(n2482), .I4(n2483), .I5(n2484), 
        .O(n2459) );
  AND4_GATE U3449 ( .I1(n2485), .I2(n2486), .I3(n2487), .I4(n2488), .O(n2484)
         );
  NAND_GATE U3450 ( .I1(n2154), .I2(\registres[17][30] ), .O(n2488) );
  NAND_GATE U3451 ( .I1(n2155), .I2(\registres[19][30] ), .O(n2487) );
  NAND_GATE U3452 ( .I1(n2156), .I2(\registres[21][30] ), .O(n2486) );
  NAND_GATE U3453 ( .I1(n2157), .I2(\registres[6][30] ), .O(n2485) );
  NAND_GATE U3454 ( .I1(n2158), .I2(\registres[7][30] ), .O(n2483) );
  NAND_GATE U3455 ( .I1(n2159), .I2(\registres[30][30] ), .O(n2482) );
  NAND_GATE U3456 ( .I1(n2160), .I2(\registres[31][30] ), .O(n2481) );
  NAND_GATE U3457 ( .I1(n2161), .I2(\registres[14][30] ), .O(n2480) );
  AND4_GATE U3458 ( .I1(n2489), .I2(n2490), .I3(n2491), .I4(n2492), .O(n2458)
         );
  AND4_GATE U3459 ( .I1(n2493), .I2(n2494), .I3(n2495), .I4(n2496), .O(n2492)
         );
  NAND_GATE U3460 ( .I1(n2170), .I2(\registres[22][30] ), .O(n2496) );
  NAND_GATE U3461 ( .I1(n2171), .I2(\registres[15][30] ), .O(n2495) );
  NAND_GATE U3462 ( .I1(n2172), .I2(\registres[23][30] ), .O(n2494) );
  NAND_GATE U3463 ( .I1(n2173), .I2(\registres[4][30] ), .O(n2493) );
  NAND_GATE U3464 ( .I1(n2174), .I2(\registres[8][30] ), .O(n2491) );
  NAND_GATE U3465 ( .I1(n2175), .I2(\registres[2][30] ), .O(n2490) );
  NAND_GATE U3466 ( .I1(n2176), .I2(\registres[16][30] ), .O(n2489) );
  AND_GATE U3467 ( .I1(n2497), .I2(n2105), .O(data_src2[2]) );
  NAND4_GATE U3468 ( .I1(n2498), .I2(n2499), .I3(n2500), .I4(n2501), .O(n2497)
         );
  AND5_GATE U3469 ( .I1(n2502), .I2(n2503), .I3(n2504), .I4(n2505), .I5(n2506), 
        .O(n2501) );
  AND4_GATE U3470 ( .I1(n2507), .I2(n2508), .I3(n2509), .I4(n2510), .O(n2506)
         );
  NAND_GATE U3471 ( .I1(n2120), .I2(\registres[24][2] ), .O(n2510) );
  NAND_GATE U3472 ( .I1(n2121), .I2(\registres[25][2] ), .O(n2509) );
  NAND_GATE U3473 ( .I1(n2122), .I2(\registres[3][2] ), .O(n2508) );
  NAND_GATE U3474 ( .I1(n2123), .I2(\registres[26][2] ), .O(n2507) );
  NAND_GATE U3475 ( .I1(n2124), .I2(\registres[27][2] ), .O(n2505) );
  NAND_GATE U3476 ( .I1(n2125), .I2(\registres[10][2] ), .O(n2504) );
  NAND_GATE U3477 ( .I1(n2126), .I2(\registres[18][2] ), .O(n2503) );
  NAND_GATE U3478 ( .I1(n2127), .I2(\registres[5][2] ), .O(n2502) );
  AND5_GATE U3479 ( .I1(n2511), .I2(n2512), .I3(n2513), .I4(n2514), .I5(n2515), 
        .O(n2500) );
  AND4_GATE U3480 ( .I1(n2516), .I2(n2517), .I3(n2518), .I4(n2519), .O(n2515)
         );
  NAND_GATE U3481 ( .I1(n2137), .I2(\registres[28][2] ), .O(n2519) );
  NAND_GATE U3482 ( .I1(n2138), .I2(\registres[29][2] ), .O(n2518) );
  NAND_GATE U3483 ( .I1(n2139), .I2(\registres[12][2] ), .O(n2517) );
  NAND_GATE U3484 ( .I1(n2140), .I2(\registres[20][2] ), .O(n2516) );
  NAND_GATE U3485 ( .I1(n2141), .I2(\registres[1][2] ), .O(n2514) );
  NAND_GATE U3486 ( .I1(n2142), .I2(\registres[9][2] ), .O(n2513) );
  NAND_GATE U3487 ( .I1(n2143), .I2(\registres[11][2] ), .O(n2512) );
  NAND_GATE U3488 ( .I1(n2144), .I2(\registres[13][2] ), .O(n2511) );
  AND5_GATE U3489 ( .I1(n2520), .I2(n2521), .I3(n2522), .I4(n2523), .I5(n2524), 
        .O(n2499) );
  AND4_GATE U3490 ( .I1(n2525), .I2(n2526), .I3(n2527), .I4(n2528), .O(n2524)
         );
  NAND_GATE U3491 ( .I1(n2154), .I2(\registres[17][2] ), .O(n2528) );
  NAND_GATE U3492 ( .I1(n2155), .I2(\registres[19][2] ), .O(n2527) );
  NAND_GATE U3493 ( .I1(n2156), .I2(\registres[21][2] ), .O(n2526) );
  NAND_GATE U3494 ( .I1(n2157), .I2(\registres[6][2] ), .O(n2525) );
  NAND_GATE U3495 ( .I1(n2158), .I2(\registres[7][2] ), .O(n2523) );
  NAND_GATE U3496 ( .I1(n2159), .I2(\registres[30][2] ), .O(n2522) );
  NAND_GATE U3497 ( .I1(n2160), .I2(\registres[31][2] ), .O(n2521) );
  NAND_GATE U3498 ( .I1(n2161), .I2(\registres[14][2] ), .O(n2520) );
  AND4_GATE U3499 ( .I1(n2529), .I2(n2530), .I3(n2531), .I4(n2532), .O(n2498)
         );
  AND4_GATE U3500 ( .I1(n2533), .I2(n2534), .I3(n2535), .I4(n2536), .O(n2532)
         );
  NAND_GATE U3501 ( .I1(n2170), .I2(\registres[22][2] ), .O(n2536) );
  NAND_GATE U3502 ( .I1(n2171), .I2(\registres[15][2] ), .O(n2535) );
  NAND_GATE U3503 ( .I1(n2172), .I2(\registres[23][2] ), .O(n2534) );
  NAND_GATE U3504 ( .I1(n2173), .I2(\registres[4][2] ), .O(n2533) );
  NAND_GATE U3505 ( .I1(n2174), .I2(\registres[8][2] ), .O(n2531) );
  NAND_GATE U3506 ( .I1(n2175), .I2(\registres[2][2] ), .O(n2530) );
  NAND_GATE U3507 ( .I1(n2176), .I2(\registres[16][2] ), .O(n2529) );
  AND_GATE U3508 ( .I1(n2537), .I2(n2105), .O(data_src2[29]) );
  NAND4_GATE U3509 ( .I1(n2538), .I2(n2539), .I3(n2540), .I4(n2541), .O(n2537)
         );
  AND5_GATE U3510 ( .I1(n2542), .I2(n2543), .I3(n2544), .I4(n2545), .I5(n2546), 
        .O(n2541) );
  AND4_GATE U3511 ( .I1(n2547), .I2(n2548), .I3(n2549), .I4(n2550), .O(n2546)
         );
  NAND_GATE U3512 ( .I1(n2120), .I2(\registres[24][29] ), .O(n2550) );
  NAND_GATE U3513 ( .I1(n2121), .I2(\registres[25][29] ), .O(n2549) );
  NAND_GATE U3514 ( .I1(n2122), .I2(\registres[3][29] ), .O(n2548) );
  NAND_GATE U3515 ( .I1(n2123), .I2(\registres[26][29] ), .O(n2547) );
  NAND_GATE U3516 ( .I1(n2124), .I2(\registres[27][29] ), .O(n2545) );
  NAND_GATE U3517 ( .I1(n2125), .I2(\registres[10][29] ), .O(n2544) );
  NAND_GATE U3518 ( .I1(n2126), .I2(\registres[18][29] ), .O(n2543) );
  NAND_GATE U3519 ( .I1(n2127), .I2(\registres[5][29] ), .O(n2542) );
  AND5_GATE U3520 ( .I1(n2551), .I2(n2552), .I3(n2553), .I4(n2554), .I5(n2555), 
        .O(n2540) );
  AND4_GATE U3521 ( .I1(n2556), .I2(n2557), .I3(n2558), .I4(n2559), .O(n2555)
         );
  NAND_GATE U3522 ( .I1(n2137), .I2(\registres[28][29] ), .O(n2559) );
  NAND_GATE U3523 ( .I1(n2138), .I2(\registres[29][29] ), .O(n2558) );
  NAND_GATE U3524 ( .I1(n2139), .I2(\registres[12][29] ), .O(n2557) );
  NAND_GATE U3525 ( .I1(n2140), .I2(\registres[20][29] ), .O(n2556) );
  NAND_GATE U3526 ( .I1(n2141), .I2(\registres[1][29] ), .O(n2554) );
  NAND_GATE U3527 ( .I1(n2142), .I2(\registres[9][29] ), .O(n2553) );
  NAND_GATE U3528 ( .I1(n2143), .I2(\registres[11][29] ), .O(n2552) );
  NAND_GATE U3529 ( .I1(n2144), .I2(\registres[13][29] ), .O(n2551) );
  AND5_GATE U3530 ( .I1(n2560), .I2(n2561), .I3(n2562), .I4(n2563), .I5(n2564), 
        .O(n2539) );
  AND4_GATE U3531 ( .I1(n2565), .I2(n2566), .I3(n2567), .I4(n2568), .O(n2564)
         );
  NAND_GATE U3532 ( .I1(n2154), .I2(\registres[17][29] ), .O(n2568) );
  NAND_GATE U3533 ( .I1(n2155), .I2(\registres[19][29] ), .O(n2567) );
  NAND_GATE U3534 ( .I1(n2156), .I2(\registres[21][29] ), .O(n2566) );
  NAND_GATE U3535 ( .I1(n2157), .I2(\registres[6][29] ), .O(n2565) );
  NAND_GATE U3536 ( .I1(n2158), .I2(\registres[7][29] ), .O(n2563) );
  NAND_GATE U3537 ( .I1(n2159), .I2(\registres[30][29] ), .O(n2562) );
  NAND_GATE U3538 ( .I1(n2160), .I2(\registres[31][29] ), .O(n2561) );
  NAND_GATE U3539 ( .I1(n2161), .I2(\registres[14][29] ), .O(n2560) );
  AND4_GATE U3540 ( .I1(n2569), .I2(n2570), .I3(n2571), .I4(n2572), .O(n2538)
         );
  AND4_GATE U3541 ( .I1(n2573), .I2(n2574), .I3(n2575), .I4(n2576), .O(n2572)
         );
  NAND_GATE U3542 ( .I1(n2170), .I2(\registres[22][29] ), .O(n2576) );
  NAND_GATE U3543 ( .I1(n2171), .I2(\registres[15][29] ), .O(n2575) );
  NAND_GATE U3544 ( .I1(n2172), .I2(\registres[23][29] ), .O(n2574) );
  NAND_GATE U3545 ( .I1(n2173), .I2(\registres[4][29] ), .O(n2573) );
  NAND_GATE U3546 ( .I1(n2174), .I2(\registres[8][29] ), .O(n2571) );
  NAND_GATE U3547 ( .I1(n2175), .I2(\registres[2][29] ), .O(n2570) );
  NAND_GATE U3548 ( .I1(n2176), .I2(\registres[16][29] ), .O(n2569) );
  AND_GATE U3549 ( .I1(n2577), .I2(n2105), .O(data_src2[28]) );
  NAND4_GATE U3550 ( .I1(n2578), .I2(n2579), .I3(n2580), .I4(n2581), .O(n2577)
         );
  AND5_GATE U3551 ( .I1(n2582), .I2(n2583), .I3(n2584), .I4(n2585), .I5(n2586), 
        .O(n2581) );
  AND4_GATE U3552 ( .I1(n2587), .I2(n2588), .I3(n2589), .I4(n2590), .O(n2586)
         );
  NAND_GATE U3553 ( .I1(n2120), .I2(\registres[24][28] ), .O(n2590) );
  NAND_GATE U3554 ( .I1(n2121), .I2(\registres[25][28] ), .O(n2589) );
  NAND_GATE U3555 ( .I1(n2122), .I2(\registres[3][28] ), .O(n2588) );
  NAND_GATE U3556 ( .I1(n2123), .I2(\registres[26][28] ), .O(n2587) );
  NAND_GATE U3557 ( .I1(n2124), .I2(\registres[27][28] ), .O(n2585) );
  NAND_GATE U3558 ( .I1(n2125), .I2(\registres[10][28] ), .O(n2584) );
  NAND_GATE U3559 ( .I1(n2126), .I2(\registres[18][28] ), .O(n2583) );
  NAND_GATE U3560 ( .I1(n2127), .I2(\registres[5][28] ), .O(n2582) );
  AND5_GATE U3561 ( .I1(n2591), .I2(n2592), .I3(n2593), .I4(n2594), .I5(n2595), 
        .O(n2580) );
  AND4_GATE U3562 ( .I1(n2596), .I2(n2597), .I3(n2598), .I4(n2599), .O(n2595)
         );
  NAND_GATE U3563 ( .I1(n2137), .I2(\registres[28][28] ), .O(n2599) );
  NAND_GATE U3564 ( .I1(n2138), .I2(\registres[29][28] ), .O(n2598) );
  NAND_GATE U3565 ( .I1(n2139), .I2(\registres[12][28] ), .O(n2597) );
  NAND_GATE U3566 ( .I1(n2140), .I2(\registres[20][28] ), .O(n2596) );
  NAND_GATE U3567 ( .I1(n2141), .I2(\registres[1][28] ), .O(n2594) );
  NAND_GATE U3568 ( .I1(n2142), .I2(\registres[9][28] ), .O(n2593) );
  NAND_GATE U3569 ( .I1(n2143), .I2(\registres[11][28] ), .O(n2592) );
  NAND_GATE U3570 ( .I1(n2144), .I2(\registres[13][28] ), .O(n2591) );
  AND5_GATE U3571 ( .I1(n2600), .I2(n2601), .I3(n2602), .I4(n2603), .I5(n2604), 
        .O(n2579) );
  AND4_GATE U3572 ( .I1(n2605), .I2(n2606), .I3(n2607), .I4(n2608), .O(n2604)
         );
  NAND_GATE U3573 ( .I1(n2154), .I2(\registres[17][28] ), .O(n2608) );
  NAND_GATE U3574 ( .I1(n2155), .I2(\registres[19][28] ), .O(n2607) );
  NAND_GATE U3575 ( .I1(n2156), .I2(\registres[21][28] ), .O(n2606) );
  NAND_GATE U3576 ( .I1(n2157), .I2(\registres[6][28] ), .O(n2605) );
  NAND_GATE U3577 ( .I1(n2158), .I2(\registres[7][28] ), .O(n2603) );
  NAND_GATE U3578 ( .I1(n2159), .I2(\registres[30][28] ), .O(n2602) );
  NAND_GATE U3579 ( .I1(n2160), .I2(\registres[31][28] ), .O(n2601) );
  NAND_GATE U3580 ( .I1(n2161), .I2(\registres[14][28] ), .O(n2600) );
  AND4_GATE U3581 ( .I1(n2609), .I2(n2610), .I3(n2611), .I4(n2612), .O(n2578)
         );
  AND4_GATE U3582 ( .I1(n2613), .I2(n2614), .I3(n2615), .I4(n2616), .O(n2612)
         );
  NAND_GATE U3583 ( .I1(n2170), .I2(\registres[22][28] ), .O(n2616) );
  NAND_GATE U3584 ( .I1(n2171), .I2(\registres[15][28] ), .O(n2615) );
  NAND_GATE U3585 ( .I1(n2172), .I2(\registres[23][28] ), .O(n2614) );
  NAND_GATE U3586 ( .I1(n2173), .I2(\registres[4][28] ), .O(n2613) );
  NAND_GATE U3587 ( .I1(n2174), .I2(\registres[8][28] ), .O(n2611) );
  NAND_GATE U3588 ( .I1(n2175), .I2(\registres[2][28] ), .O(n2610) );
  NAND_GATE U3589 ( .I1(n2176), .I2(\registres[16][28] ), .O(n2609) );
  AND_GATE U3590 ( .I1(n2617), .I2(n2105), .O(data_src2[27]) );
  NAND4_GATE U3591 ( .I1(n2618), .I2(n2619), .I3(n2620), .I4(n2621), .O(n2617)
         );
  AND5_GATE U3592 ( .I1(n2622), .I2(n2623), .I3(n2624), .I4(n2625), .I5(n2626), 
        .O(n2621) );
  AND4_GATE U3593 ( .I1(n2627), .I2(n2628), .I3(n2629), .I4(n2630), .O(n2626)
         );
  NAND_GATE U3594 ( .I1(n2120), .I2(\registres[24][27] ), .O(n2630) );
  NAND_GATE U3595 ( .I1(n2121), .I2(\registres[25][27] ), .O(n2629) );
  NAND_GATE U3596 ( .I1(n2122), .I2(\registres[3][27] ), .O(n2628) );
  NAND_GATE U3597 ( .I1(n2123), .I2(\registres[26][27] ), .O(n2627) );
  NAND_GATE U3598 ( .I1(n2124), .I2(\registres[27][27] ), .O(n2625) );
  NAND_GATE U3599 ( .I1(n2125), .I2(\registres[10][27] ), .O(n2624) );
  NAND_GATE U3600 ( .I1(n2126), .I2(\registres[18][27] ), .O(n2623) );
  NAND_GATE U3601 ( .I1(n2127), .I2(\registres[5][27] ), .O(n2622) );
  AND5_GATE U3602 ( .I1(n2631), .I2(n2632), .I3(n2633), .I4(n2634), .I5(n2635), 
        .O(n2620) );
  AND4_GATE U3603 ( .I1(n2636), .I2(n2637), .I3(n2638), .I4(n2639), .O(n2635)
         );
  NAND_GATE U3604 ( .I1(n2137), .I2(\registres[28][27] ), .O(n2639) );
  NAND_GATE U3605 ( .I1(n2138), .I2(\registres[29][27] ), .O(n2638) );
  NAND_GATE U3606 ( .I1(n2139), .I2(\registres[12][27] ), .O(n2637) );
  NAND_GATE U3607 ( .I1(n2140), .I2(\registres[20][27] ), .O(n2636) );
  NAND_GATE U3608 ( .I1(n2141), .I2(\registres[1][27] ), .O(n2634) );
  NAND_GATE U3609 ( .I1(n2142), .I2(\registres[9][27] ), .O(n2633) );
  NAND_GATE U3610 ( .I1(n2143), .I2(\registres[11][27] ), .O(n2632) );
  NAND_GATE U3611 ( .I1(n2144), .I2(\registres[13][27] ), .O(n2631) );
  AND5_GATE U3612 ( .I1(n2640), .I2(n2641), .I3(n2642), .I4(n2643), .I5(n2644), 
        .O(n2619) );
  AND4_GATE U3613 ( .I1(n2645), .I2(n2646), .I3(n2647), .I4(n2648), .O(n2644)
         );
  NAND_GATE U3614 ( .I1(n2154), .I2(\registres[17][27] ), .O(n2648) );
  NAND_GATE U3615 ( .I1(n2155), .I2(\registres[19][27] ), .O(n2647) );
  NAND_GATE U3616 ( .I1(n2156), .I2(\registres[21][27] ), .O(n2646) );
  NAND_GATE U3617 ( .I1(n2157), .I2(\registres[6][27] ), .O(n2645) );
  NAND_GATE U3618 ( .I1(n2158), .I2(\registres[7][27] ), .O(n2643) );
  NAND_GATE U3619 ( .I1(n2159), .I2(\registres[30][27] ), .O(n2642) );
  NAND_GATE U3620 ( .I1(n2160), .I2(\registres[31][27] ), .O(n2641) );
  NAND_GATE U3621 ( .I1(n2161), .I2(\registres[14][27] ), .O(n2640) );
  AND4_GATE U3622 ( .I1(n2649), .I2(n2650), .I3(n2651), .I4(n2652), .O(n2618)
         );
  AND4_GATE U3623 ( .I1(n2653), .I2(n2654), .I3(n2655), .I4(n2656), .O(n2652)
         );
  NAND_GATE U3624 ( .I1(n2170), .I2(\registres[22][27] ), .O(n2656) );
  NAND_GATE U3625 ( .I1(n2171), .I2(\registres[15][27] ), .O(n2655) );
  NAND_GATE U3626 ( .I1(n2172), .I2(\registres[23][27] ), .O(n2654) );
  NAND_GATE U3627 ( .I1(n2173), .I2(\registres[4][27] ), .O(n2653) );
  NAND_GATE U3628 ( .I1(n2174), .I2(\registres[8][27] ), .O(n2651) );
  NAND_GATE U3629 ( .I1(n2175), .I2(\registres[2][27] ), .O(n2650) );
  NAND_GATE U3630 ( .I1(n2176), .I2(\registres[16][27] ), .O(n2649) );
  AND_GATE U3631 ( .I1(n2657), .I2(n2105), .O(data_src2[26]) );
  NAND4_GATE U3632 ( .I1(n2658), .I2(n2659), .I3(n2660), .I4(n2661), .O(n2657)
         );
  AND5_GATE U3633 ( .I1(n2662), .I2(n2663), .I3(n2664), .I4(n2665), .I5(n2666), 
        .O(n2661) );
  AND4_GATE U3634 ( .I1(n2667), .I2(n2668), .I3(n2669), .I4(n2670), .O(n2666)
         );
  NAND_GATE U3635 ( .I1(n2120), .I2(\registres[24][26] ), .O(n2670) );
  NAND_GATE U3636 ( .I1(n2121), .I2(\registres[25][26] ), .O(n2669) );
  NAND_GATE U3637 ( .I1(n2122), .I2(\registres[3][26] ), .O(n2668) );
  NAND_GATE U3638 ( .I1(n2123), .I2(\registres[26][26] ), .O(n2667) );
  NAND_GATE U3639 ( .I1(n2124), .I2(\registres[27][26] ), .O(n2665) );
  NAND_GATE U3640 ( .I1(n2125), .I2(\registres[10][26] ), .O(n2664) );
  NAND_GATE U3641 ( .I1(n2126), .I2(\registres[18][26] ), .O(n2663) );
  NAND_GATE U3642 ( .I1(n2127), .I2(\registres[5][26] ), .O(n2662) );
  AND5_GATE U3643 ( .I1(n2671), .I2(n2672), .I3(n2673), .I4(n2674), .I5(n2675), 
        .O(n2660) );
  AND4_GATE U3644 ( .I1(n2676), .I2(n2677), .I3(n2678), .I4(n2679), .O(n2675)
         );
  NAND_GATE U3645 ( .I1(n2137), .I2(\registres[28][26] ), .O(n2679) );
  NAND_GATE U3646 ( .I1(n2138), .I2(\registres[29][26] ), .O(n2678) );
  NAND_GATE U3647 ( .I1(n2139), .I2(\registres[12][26] ), .O(n2677) );
  NAND_GATE U3648 ( .I1(n2140), .I2(\registres[20][26] ), .O(n2676) );
  NAND_GATE U3649 ( .I1(n2141), .I2(\registres[1][26] ), .O(n2674) );
  NAND_GATE U3650 ( .I1(n2142), .I2(\registres[9][26] ), .O(n2673) );
  NAND_GATE U3651 ( .I1(n2143), .I2(\registres[11][26] ), .O(n2672) );
  NAND_GATE U3652 ( .I1(n2144), .I2(\registres[13][26] ), .O(n2671) );
  AND5_GATE U3653 ( .I1(n2680), .I2(n2681), .I3(n2682), .I4(n2683), .I5(n2684), 
        .O(n2659) );
  AND4_GATE U3654 ( .I1(n2685), .I2(n2686), .I3(n2687), .I4(n2688), .O(n2684)
         );
  NAND_GATE U3655 ( .I1(n2154), .I2(\registres[17][26] ), .O(n2688) );
  NAND_GATE U3656 ( .I1(n2155), .I2(\registres[19][26] ), .O(n2687) );
  NAND_GATE U3657 ( .I1(n2156), .I2(\registres[21][26] ), .O(n2686) );
  NAND_GATE U3658 ( .I1(n2157), .I2(\registres[6][26] ), .O(n2685) );
  NAND_GATE U3659 ( .I1(n2158), .I2(\registres[7][26] ), .O(n2683) );
  NAND_GATE U3660 ( .I1(n2159), .I2(\registres[30][26] ), .O(n2682) );
  NAND_GATE U3661 ( .I1(n2160), .I2(\registres[31][26] ), .O(n2681) );
  NAND_GATE U3662 ( .I1(n2161), .I2(\registres[14][26] ), .O(n2680) );
  AND4_GATE U3663 ( .I1(n2689), .I2(n2690), .I3(n2691), .I4(n2692), .O(n2658)
         );
  AND4_GATE U3664 ( .I1(n2693), .I2(n2694), .I3(n2695), .I4(n2696), .O(n2692)
         );
  NAND_GATE U3665 ( .I1(n2170), .I2(\registres[22][26] ), .O(n2696) );
  NAND_GATE U3666 ( .I1(n2171), .I2(\registres[15][26] ), .O(n2695) );
  NAND_GATE U3667 ( .I1(n2172), .I2(\registres[23][26] ), .O(n2694) );
  NAND_GATE U3668 ( .I1(n2173), .I2(\registres[4][26] ), .O(n2693) );
  NAND_GATE U3669 ( .I1(n2174), .I2(\registres[8][26] ), .O(n2691) );
  NAND_GATE U3670 ( .I1(n2175), .I2(\registres[2][26] ), .O(n2690) );
  NAND_GATE U3671 ( .I1(n2176), .I2(\registres[16][26] ), .O(n2689) );
  AND_GATE U3672 ( .I1(n2697), .I2(n2105), .O(data_src2[25]) );
  NAND4_GATE U3673 ( .I1(n2698), .I2(n2699), .I3(n2700), .I4(n2701), .O(n2697)
         );
  AND5_GATE U3674 ( .I1(n2702), .I2(n2703), .I3(n2704), .I4(n2705), .I5(n2706), 
        .O(n2701) );
  AND4_GATE U3675 ( .I1(n2707), .I2(n2708), .I3(n2709), .I4(n2710), .O(n2706)
         );
  NAND_GATE U3676 ( .I1(n2120), .I2(\registres[24][25] ), .O(n2710) );
  NAND_GATE U3677 ( .I1(n2121), .I2(\registres[25][25] ), .O(n2709) );
  NAND_GATE U3678 ( .I1(n2122), .I2(\registres[3][25] ), .O(n2708) );
  NAND_GATE U3679 ( .I1(n2123), .I2(\registres[26][25] ), .O(n2707) );
  NAND_GATE U3680 ( .I1(n2124), .I2(\registres[27][25] ), .O(n2705) );
  NAND_GATE U3681 ( .I1(n2125), .I2(\registres[10][25] ), .O(n2704) );
  NAND_GATE U3682 ( .I1(n2126), .I2(\registres[18][25] ), .O(n2703) );
  NAND_GATE U3683 ( .I1(n2127), .I2(\registres[5][25] ), .O(n2702) );
  AND5_GATE U3684 ( .I1(n2711), .I2(n2712), .I3(n2713), .I4(n2714), .I5(n2715), 
        .O(n2700) );
  AND4_GATE U3685 ( .I1(n2716), .I2(n2717), .I3(n2718), .I4(n2719), .O(n2715)
         );
  NAND_GATE U3686 ( .I1(n2137), .I2(\registres[28][25] ), .O(n2719) );
  NAND_GATE U3687 ( .I1(n2138), .I2(\registres[29][25] ), .O(n2718) );
  NAND_GATE U3688 ( .I1(n2139), .I2(\registres[12][25] ), .O(n2717) );
  NAND_GATE U3689 ( .I1(n2140), .I2(\registres[20][25] ), .O(n2716) );
  NAND_GATE U3690 ( .I1(n2141), .I2(\registres[1][25] ), .O(n2714) );
  NAND_GATE U3691 ( .I1(n2142), .I2(\registres[9][25] ), .O(n2713) );
  NAND_GATE U3692 ( .I1(n2143), .I2(\registres[11][25] ), .O(n2712) );
  NAND_GATE U3693 ( .I1(n2144), .I2(\registres[13][25] ), .O(n2711) );
  AND5_GATE U3694 ( .I1(n2720), .I2(n2721), .I3(n2722), .I4(n2723), .I5(n2724), 
        .O(n2699) );
  AND4_GATE U3695 ( .I1(n2725), .I2(n2726), .I3(n2727), .I4(n2728), .O(n2724)
         );
  NAND_GATE U3696 ( .I1(n2154), .I2(\registres[17][25] ), .O(n2728) );
  NAND_GATE U3697 ( .I1(n2155), .I2(\registres[19][25] ), .O(n2727) );
  NAND_GATE U3698 ( .I1(n2156), .I2(\registres[21][25] ), .O(n2726) );
  NAND_GATE U3699 ( .I1(n2157), .I2(\registres[6][25] ), .O(n2725) );
  NAND_GATE U3700 ( .I1(n2158), .I2(\registres[7][25] ), .O(n2723) );
  NAND_GATE U3701 ( .I1(n2159), .I2(\registres[30][25] ), .O(n2722) );
  NAND_GATE U3702 ( .I1(n2160), .I2(\registres[31][25] ), .O(n2721) );
  NAND_GATE U3703 ( .I1(n2161), .I2(\registres[14][25] ), .O(n2720) );
  AND4_GATE U3704 ( .I1(n2729), .I2(n2730), .I3(n2731), .I4(n2732), .O(n2698)
         );
  AND4_GATE U3705 ( .I1(n2733), .I2(n2734), .I3(n2735), .I4(n2736), .O(n2732)
         );
  NAND_GATE U3706 ( .I1(n2170), .I2(\registres[22][25] ), .O(n2736) );
  NAND_GATE U3707 ( .I1(n2171), .I2(\registres[15][25] ), .O(n2735) );
  NAND_GATE U3708 ( .I1(n2172), .I2(\registres[23][25] ), .O(n2734) );
  NAND_GATE U3709 ( .I1(n2173), .I2(\registres[4][25] ), .O(n2733) );
  NAND_GATE U3710 ( .I1(n2174), .I2(\registres[8][25] ), .O(n2731) );
  NAND_GATE U3711 ( .I1(n2175), .I2(\registres[2][25] ), .O(n2730) );
  NAND_GATE U3712 ( .I1(n2176), .I2(\registres[16][25] ), .O(n2729) );
  AND_GATE U3713 ( .I1(n2737), .I2(n2105), .O(data_src2[24]) );
  NAND4_GATE U3714 ( .I1(n2738), .I2(n2739), .I3(n2740), .I4(n2741), .O(n2737)
         );
  AND5_GATE U3715 ( .I1(n2742), .I2(n2743), .I3(n2744), .I4(n2745), .I5(n2746), 
        .O(n2741) );
  AND4_GATE U3716 ( .I1(n2747), .I2(n2748), .I3(n2749), .I4(n2750), .O(n2746)
         );
  NAND_GATE U3717 ( .I1(n2120), .I2(\registres[24][24] ), .O(n2750) );
  NAND_GATE U3718 ( .I1(n2121), .I2(\registres[25][24] ), .O(n2749) );
  NAND_GATE U3719 ( .I1(n2122), .I2(\registres[3][24] ), .O(n2748) );
  NAND_GATE U3720 ( .I1(n2123), .I2(\registres[26][24] ), .O(n2747) );
  NAND_GATE U3721 ( .I1(n2124), .I2(\registres[27][24] ), .O(n2745) );
  NAND_GATE U3722 ( .I1(n2125), .I2(\registres[10][24] ), .O(n2744) );
  NAND_GATE U3723 ( .I1(n2126), .I2(\registres[18][24] ), .O(n2743) );
  NAND_GATE U3724 ( .I1(n2127), .I2(\registres[5][24] ), .O(n2742) );
  AND5_GATE U3725 ( .I1(n2751), .I2(n2752), .I3(n2753), .I4(n2754), .I5(n2755), 
        .O(n2740) );
  AND4_GATE U3726 ( .I1(n2756), .I2(n2757), .I3(n2758), .I4(n2759), .O(n2755)
         );
  NAND_GATE U3727 ( .I1(n2137), .I2(\registres[28][24] ), .O(n2759) );
  NAND_GATE U3728 ( .I1(n2138), .I2(\registres[29][24] ), .O(n2758) );
  NAND_GATE U3729 ( .I1(n2139), .I2(\registres[12][24] ), .O(n2757) );
  NAND_GATE U3730 ( .I1(n2140), .I2(\registres[20][24] ), .O(n2756) );
  NAND_GATE U3731 ( .I1(n2141), .I2(\registres[1][24] ), .O(n2754) );
  NAND_GATE U3732 ( .I1(n2142), .I2(\registres[9][24] ), .O(n2753) );
  NAND_GATE U3733 ( .I1(n2143), .I2(\registres[11][24] ), .O(n2752) );
  NAND_GATE U3734 ( .I1(n2144), .I2(\registres[13][24] ), .O(n2751) );
  AND5_GATE U3735 ( .I1(n2760), .I2(n2761), .I3(n2762), .I4(n2763), .I5(n2764), 
        .O(n2739) );
  AND4_GATE U3736 ( .I1(n2765), .I2(n2766), .I3(n2767), .I4(n2768), .O(n2764)
         );
  NAND_GATE U3737 ( .I1(n2154), .I2(\registres[17][24] ), .O(n2768) );
  NAND_GATE U3738 ( .I1(n2155), .I2(\registres[19][24] ), .O(n2767) );
  NAND_GATE U3739 ( .I1(n2156), .I2(\registres[21][24] ), .O(n2766) );
  NAND_GATE U3740 ( .I1(n2157), .I2(\registres[6][24] ), .O(n2765) );
  NAND_GATE U3741 ( .I1(n2158), .I2(\registres[7][24] ), .O(n2763) );
  NAND_GATE U3742 ( .I1(n2159), .I2(\registres[30][24] ), .O(n2762) );
  NAND_GATE U3743 ( .I1(n2160), .I2(\registres[31][24] ), .O(n2761) );
  NAND_GATE U3744 ( .I1(n2161), .I2(\registres[14][24] ), .O(n2760) );
  AND4_GATE U3745 ( .I1(n2769), .I2(n2770), .I3(n2771), .I4(n2772), .O(n2738)
         );
  AND4_GATE U3746 ( .I1(n2773), .I2(n2774), .I3(n2775), .I4(n2776), .O(n2772)
         );
  NAND_GATE U3747 ( .I1(n2170), .I2(\registres[22][24] ), .O(n2776) );
  NAND_GATE U3748 ( .I1(n2171), .I2(\registres[15][24] ), .O(n2775) );
  NAND_GATE U3749 ( .I1(n2172), .I2(\registres[23][24] ), .O(n2774) );
  NAND_GATE U3750 ( .I1(n2173), .I2(\registres[4][24] ), .O(n2773) );
  NAND_GATE U3751 ( .I1(n2174), .I2(\registres[8][24] ), .O(n2771) );
  NAND_GATE U3752 ( .I1(n2175), .I2(\registres[2][24] ), .O(n2770) );
  NAND_GATE U3753 ( .I1(n2176), .I2(\registres[16][24] ), .O(n2769) );
  AND_GATE U3754 ( .I1(n2777), .I2(n2105), .O(data_src2[23]) );
  NAND4_GATE U3755 ( .I1(n2778), .I2(n2779), .I3(n2780), .I4(n2781), .O(n2777)
         );
  AND5_GATE U3756 ( .I1(n2782), .I2(n2783), .I3(n2784), .I4(n2785), .I5(n2786), 
        .O(n2781) );
  AND4_GATE U3757 ( .I1(n2787), .I2(n2788), .I3(n2789), .I4(n2790), .O(n2786)
         );
  NAND_GATE U3758 ( .I1(n2120), .I2(\registres[24][23] ), .O(n2790) );
  NAND_GATE U3759 ( .I1(n2121), .I2(\registres[25][23] ), .O(n2789) );
  NAND_GATE U3760 ( .I1(n2122), .I2(\registres[3][23] ), .O(n2788) );
  NAND_GATE U3761 ( .I1(n2123), .I2(\registres[26][23] ), .O(n2787) );
  NAND_GATE U3762 ( .I1(n2124), .I2(\registres[27][23] ), .O(n2785) );
  NAND_GATE U3763 ( .I1(n2125), .I2(\registres[10][23] ), .O(n2784) );
  NAND_GATE U3764 ( .I1(n2126), .I2(\registres[18][23] ), .O(n2783) );
  NAND_GATE U3765 ( .I1(n2127), .I2(\registres[5][23] ), .O(n2782) );
  AND5_GATE U3766 ( .I1(n2791), .I2(n2792), .I3(n2793), .I4(n2794), .I5(n2795), 
        .O(n2780) );
  AND4_GATE U3767 ( .I1(n2796), .I2(n2797), .I3(n2798), .I4(n2799), .O(n2795)
         );
  NAND_GATE U3768 ( .I1(n2137), .I2(\registres[28][23] ), .O(n2799) );
  NAND_GATE U3769 ( .I1(n2138), .I2(\registres[29][23] ), .O(n2798) );
  NAND_GATE U3770 ( .I1(n2139), .I2(\registres[12][23] ), .O(n2797) );
  NAND_GATE U3771 ( .I1(n2140), .I2(\registres[20][23] ), .O(n2796) );
  NAND_GATE U3772 ( .I1(n2141), .I2(\registres[1][23] ), .O(n2794) );
  NAND_GATE U3773 ( .I1(n2142), .I2(\registres[9][23] ), .O(n2793) );
  NAND_GATE U3774 ( .I1(n2143), .I2(\registres[11][23] ), .O(n2792) );
  NAND_GATE U3775 ( .I1(n2144), .I2(\registres[13][23] ), .O(n2791) );
  AND5_GATE U3776 ( .I1(n2800), .I2(n2801), .I3(n2802), .I4(n2803), .I5(n2804), 
        .O(n2779) );
  AND4_GATE U3777 ( .I1(n2805), .I2(n2806), .I3(n2807), .I4(n2808), .O(n2804)
         );
  NAND_GATE U3778 ( .I1(n2154), .I2(\registres[17][23] ), .O(n2808) );
  NAND_GATE U3779 ( .I1(n2155), .I2(\registres[19][23] ), .O(n2807) );
  NAND_GATE U3780 ( .I1(n2156), .I2(\registres[21][23] ), .O(n2806) );
  NAND_GATE U3781 ( .I1(n2157), .I2(\registres[6][23] ), .O(n2805) );
  NAND_GATE U3782 ( .I1(n2158), .I2(\registres[7][23] ), .O(n2803) );
  NAND_GATE U3783 ( .I1(n2159), .I2(\registres[30][23] ), .O(n2802) );
  NAND_GATE U3784 ( .I1(n2160), .I2(\registres[31][23] ), .O(n2801) );
  NAND_GATE U3785 ( .I1(n2161), .I2(\registres[14][23] ), .O(n2800) );
  AND4_GATE U3786 ( .I1(n2809), .I2(n2810), .I3(n2811), .I4(n2812), .O(n2778)
         );
  AND4_GATE U3787 ( .I1(n2813), .I2(n2814), .I3(n2815), .I4(n2816), .O(n2812)
         );
  NAND_GATE U3788 ( .I1(n2170), .I2(\registres[22][23] ), .O(n2816) );
  NAND_GATE U3789 ( .I1(n2171), .I2(\registres[15][23] ), .O(n2815) );
  NAND_GATE U3790 ( .I1(n2172), .I2(\registres[23][23] ), .O(n2814) );
  NAND_GATE U3791 ( .I1(n2173), .I2(\registres[4][23] ), .O(n2813) );
  NAND_GATE U3792 ( .I1(n2174), .I2(\registres[8][23] ), .O(n2811) );
  NAND_GATE U3793 ( .I1(n2175), .I2(\registres[2][23] ), .O(n2810) );
  NAND_GATE U3794 ( .I1(n2176), .I2(\registres[16][23] ), .O(n2809) );
  AND_GATE U3795 ( .I1(n2817), .I2(n2105), .O(data_src2[22]) );
  NAND4_GATE U3796 ( .I1(n2818), .I2(n2819), .I3(n2820), .I4(n2821), .O(n2817)
         );
  AND5_GATE U3797 ( .I1(n2822), .I2(n2823), .I3(n2824), .I4(n2825), .I5(n2826), 
        .O(n2821) );
  AND4_GATE U3798 ( .I1(n2827), .I2(n2828), .I3(n2829), .I4(n2830), .O(n2826)
         );
  NAND_GATE U3799 ( .I1(n2120), .I2(\registres[24][22] ), .O(n2830) );
  NAND_GATE U3800 ( .I1(n2121), .I2(\registres[25][22] ), .O(n2829) );
  NAND_GATE U3801 ( .I1(n2122), .I2(\registres[3][22] ), .O(n2828) );
  NAND_GATE U3802 ( .I1(n2123), .I2(\registres[26][22] ), .O(n2827) );
  NAND_GATE U3803 ( .I1(n2124), .I2(\registres[27][22] ), .O(n2825) );
  NAND_GATE U3804 ( .I1(n2125), .I2(\registres[10][22] ), .O(n2824) );
  NAND_GATE U3805 ( .I1(n2126), .I2(\registres[18][22] ), .O(n2823) );
  NAND_GATE U3806 ( .I1(n2127), .I2(\registres[5][22] ), .O(n2822) );
  AND5_GATE U3807 ( .I1(n2831), .I2(n2832), .I3(n2833), .I4(n2834), .I5(n2835), 
        .O(n2820) );
  AND4_GATE U3808 ( .I1(n2836), .I2(n2837), .I3(n2838), .I4(n2839), .O(n2835)
         );
  NAND_GATE U3809 ( .I1(n2137), .I2(\registres[28][22] ), .O(n2839) );
  NAND_GATE U3810 ( .I1(n2138), .I2(\registres[29][22] ), .O(n2838) );
  NAND_GATE U3811 ( .I1(n2139), .I2(\registres[12][22] ), .O(n2837) );
  NAND_GATE U3812 ( .I1(n2140), .I2(\registres[20][22] ), .O(n2836) );
  NAND_GATE U3813 ( .I1(n2141), .I2(\registres[1][22] ), .O(n2834) );
  NAND_GATE U3814 ( .I1(n2142), .I2(\registres[9][22] ), .O(n2833) );
  NAND_GATE U3815 ( .I1(n2143), .I2(\registres[11][22] ), .O(n2832) );
  NAND_GATE U3816 ( .I1(n2144), .I2(\registres[13][22] ), .O(n2831) );
  AND5_GATE U3817 ( .I1(n2840), .I2(n2841), .I3(n2842), .I4(n2843), .I5(n2844), 
        .O(n2819) );
  AND4_GATE U3818 ( .I1(n2845), .I2(n2846), .I3(n2847), .I4(n2848), .O(n2844)
         );
  NAND_GATE U3819 ( .I1(n2154), .I2(\registres[17][22] ), .O(n2848) );
  NAND_GATE U3820 ( .I1(n2155), .I2(\registres[19][22] ), .O(n2847) );
  NAND_GATE U3821 ( .I1(n2156), .I2(\registres[21][22] ), .O(n2846) );
  NAND_GATE U3822 ( .I1(n2157), .I2(\registres[6][22] ), .O(n2845) );
  NAND_GATE U3823 ( .I1(n2158), .I2(\registres[7][22] ), .O(n2843) );
  NAND_GATE U3824 ( .I1(n2159), .I2(\registres[30][22] ), .O(n2842) );
  NAND_GATE U3825 ( .I1(n2160), .I2(\registres[31][22] ), .O(n2841) );
  NAND_GATE U3826 ( .I1(n2161), .I2(\registres[14][22] ), .O(n2840) );
  AND4_GATE U3827 ( .I1(n2849), .I2(n2850), .I3(n2851), .I4(n2852), .O(n2818)
         );
  AND4_GATE U3828 ( .I1(n2853), .I2(n2854), .I3(n2855), .I4(n2856), .O(n2852)
         );
  NAND_GATE U3829 ( .I1(n2170), .I2(\registres[22][22] ), .O(n2856) );
  NAND_GATE U3830 ( .I1(n2171), .I2(\registres[15][22] ), .O(n2855) );
  NAND_GATE U3831 ( .I1(n2172), .I2(\registres[23][22] ), .O(n2854) );
  NAND_GATE U3832 ( .I1(n2173), .I2(\registres[4][22] ), .O(n2853) );
  NAND_GATE U3833 ( .I1(n2174), .I2(\registres[8][22] ), .O(n2851) );
  NAND_GATE U3834 ( .I1(n2175), .I2(\registres[2][22] ), .O(n2850) );
  NAND_GATE U3835 ( .I1(n2176), .I2(\registres[16][22] ), .O(n2849) );
  AND_GATE U3836 ( .I1(n2857), .I2(n2105), .O(data_src2[21]) );
  NAND4_GATE U3837 ( .I1(n2858), .I2(n2859), .I3(n2860), .I4(n2861), .O(n2857)
         );
  AND5_GATE U3838 ( .I1(n2862), .I2(n2863), .I3(n2864), .I4(n2865), .I5(n2866), 
        .O(n2861) );
  AND4_GATE U3839 ( .I1(n2867), .I2(n2868), .I3(n2869), .I4(n2870), .O(n2866)
         );
  NAND_GATE U3840 ( .I1(n2120), .I2(\registres[24][21] ), .O(n2870) );
  NAND_GATE U3841 ( .I1(n2121), .I2(\registres[25][21] ), .O(n2869) );
  NAND_GATE U3842 ( .I1(n2122), .I2(\registres[3][21] ), .O(n2868) );
  NAND_GATE U3843 ( .I1(n2123), .I2(\registres[26][21] ), .O(n2867) );
  NAND_GATE U3844 ( .I1(n2124), .I2(\registres[27][21] ), .O(n2865) );
  NAND_GATE U3845 ( .I1(n2125), .I2(\registres[10][21] ), .O(n2864) );
  NAND_GATE U3846 ( .I1(n2126), .I2(\registres[18][21] ), .O(n2863) );
  NAND_GATE U3847 ( .I1(n2127), .I2(\registres[5][21] ), .O(n2862) );
  AND5_GATE U3848 ( .I1(n2871), .I2(n2872), .I3(n2873), .I4(n2874), .I5(n2875), 
        .O(n2860) );
  AND4_GATE U3849 ( .I1(n2876), .I2(n2877), .I3(n2878), .I4(n2879), .O(n2875)
         );
  NAND_GATE U3850 ( .I1(n2137), .I2(\registres[28][21] ), .O(n2879) );
  NAND_GATE U3851 ( .I1(n2138), .I2(\registres[29][21] ), .O(n2878) );
  NAND_GATE U3852 ( .I1(n2139), .I2(\registres[12][21] ), .O(n2877) );
  NAND_GATE U3853 ( .I1(n2140), .I2(\registres[20][21] ), .O(n2876) );
  NAND_GATE U3854 ( .I1(n2141), .I2(\registres[1][21] ), .O(n2874) );
  NAND_GATE U3855 ( .I1(n2142), .I2(\registres[9][21] ), .O(n2873) );
  NAND_GATE U3856 ( .I1(n2143), .I2(\registres[11][21] ), .O(n2872) );
  NAND_GATE U3857 ( .I1(n2144), .I2(\registres[13][21] ), .O(n2871) );
  AND5_GATE U3858 ( .I1(n2880), .I2(n2881), .I3(n2882), .I4(n2883), .I5(n2884), 
        .O(n2859) );
  AND4_GATE U3859 ( .I1(n2885), .I2(n2886), .I3(n2887), .I4(n2888), .O(n2884)
         );
  NAND_GATE U3860 ( .I1(n2154), .I2(\registres[17][21] ), .O(n2888) );
  NAND_GATE U3861 ( .I1(n2155), .I2(\registres[19][21] ), .O(n2887) );
  NAND_GATE U3862 ( .I1(n2156), .I2(\registres[21][21] ), .O(n2886) );
  NAND_GATE U3863 ( .I1(n2157), .I2(\registres[6][21] ), .O(n2885) );
  NAND_GATE U3864 ( .I1(n2158), .I2(\registres[7][21] ), .O(n2883) );
  NAND_GATE U3865 ( .I1(n2159), .I2(\registres[30][21] ), .O(n2882) );
  NAND_GATE U3866 ( .I1(n2160), .I2(\registres[31][21] ), .O(n2881) );
  NAND_GATE U3867 ( .I1(n2161), .I2(\registres[14][21] ), .O(n2880) );
  AND4_GATE U3868 ( .I1(n2889), .I2(n2890), .I3(n2891), .I4(n2892), .O(n2858)
         );
  AND4_GATE U3869 ( .I1(n2893), .I2(n2894), .I3(n2895), .I4(n2896), .O(n2892)
         );
  NAND_GATE U3870 ( .I1(n2170), .I2(\registres[22][21] ), .O(n2896) );
  NAND_GATE U3871 ( .I1(n2171), .I2(\registres[15][21] ), .O(n2895) );
  NAND_GATE U3872 ( .I1(n2172), .I2(\registres[23][21] ), .O(n2894) );
  NAND_GATE U3873 ( .I1(n2173), .I2(\registres[4][21] ), .O(n2893) );
  NAND_GATE U3874 ( .I1(n2174), .I2(\registres[8][21] ), .O(n2891) );
  NAND_GATE U3875 ( .I1(n2175), .I2(\registres[2][21] ), .O(n2890) );
  NAND_GATE U3876 ( .I1(n2176), .I2(\registres[16][21] ), .O(n2889) );
  AND_GATE U3877 ( .I1(n2897), .I2(n2105), .O(data_src2[20]) );
  NAND4_GATE U3878 ( .I1(n2898), .I2(n2899), .I3(n2900), .I4(n2901), .O(n2897)
         );
  AND5_GATE U3879 ( .I1(n2902), .I2(n2903), .I3(n2904), .I4(n2905), .I5(n2906), 
        .O(n2901) );
  AND4_GATE U3880 ( .I1(n2907), .I2(n2908), .I3(n2909), .I4(n2910), .O(n2906)
         );
  NAND_GATE U3881 ( .I1(n2120), .I2(\registres[24][20] ), .O(n2910) );
  NAND_GATE U3882 ( .I1(n2121), .I2(\registres[25][20] ), .O(n2909) );
  NAND_GATE U3883 ( .I1(n2122), .I2(\registres[3][20] ), .O(n2908) );
  NAND_GATE U3884 ( .I1(n2123), .I2(\registres[26][20] ), .O(n2907) );
  NAND_GATE U3885 ( .I1(n2124), .I2(\registres[27][20] ), .O(n2905) );
  NAND_GATE U3886 ( .I1(n2125), .I2(\registres[10][20] ), .O(n2904) );
  NAND_GATE U3887 ( .I1(n2126), .I2(\registres[18][20] ), .O(n2903) );
  NAND_GATE U3888 ( .I1(n2127), .I2(\registres[5][20] ), .O(n2902) );
  AND5_GATE U3889 ( .I1(n2911), .I2(n2912), .I3(n2913), .I4(n2914), .I5(n2915), 
        .O(n2900) );
  AND4_GATE U3890 ( .I1(n2916), .I2(n2917), .I3(n2918), .I4(n2919), .O(n2915)
         );
  NAND_GATE U3891 ( .I1(n2137), .I2(\registres[28][20] ), .O(n2919) );
  NAND_GATE U3892 ( .I1(n2138), .I2(\registres[29][20] ), .O(n2918) );
  NAND_GATE U3893 ( .I1(n2139), .I2(\registres[12][20] ), .O(n2917) );
  NAND_GATE U3894 ( .I1(n2140), .I2(\registres[20][20] ), .O(n2916) );
  NAND_GATE U3895 ( .I1(n2141), .I2(\registres[1][20] ), .O(n2914) );
  NAND_GATE U3896 ( .I1(n2142), .I2(\registres[9][20] ), .O(n2913) );
  NAND_GATE U3897 ( .I1(n2143), .I2(\registres[11][20] ), .O(n2912) );
  NAND_GATE U3898 ( .I1(n2144), .I2(\registres[13][20] ), .O(n2911) );
  AND5_GATE U3899 ( .I1(n2920), .I2(n2921), .I3(n2922), .I4(n2923), .I5(n2924), 
        .O(n2899) );
  AND4_GATE U3900 ( .I1(n2925), .I2(n2926), .I3(n2927), .I4(n2928), .O(n2924)
         );
  NAND_GATE U3901 ( .I1(n2154), .I2(\registres[17][20] ), .O(n2928) );
  NAND_GATE U3902 ( .I1(n2155), .I2(\registres[19][20] ), .O(n2927) );
  NAND_GATE U3903 ( .I1(n2156), .I2(\registres[21][20] ), .O(n2926) );
  NAND_GATE U3904 ( .I1(n2157), .I2(\registres[6][20] ), .O(n2925) );
  NAND_GATE U3905 ( .I1(n2158), .I2(\registres[7][20] ), .O(n2923) );
  NAND_GATE U3906 ( .I1(n2159), .I2(\registres[30][20] ), .O(n2922) );
  NAND_GATE U3907 ( .I1(n2160), .I2(\registres[31][20] ), .O(n2921) );
  NAND_GATE U3908 ( .I1(n2161), .I2(\registres[14][20] ), .O(n2920) );
  AND4_GATE U3909 ( .I1(n2929), .I2(n2930), .I3(n2931), .I4(n2932), .O(n2898)
         );
  AND4_GATE U3910 ( .I1(n2933), .I2(n2934), .I3(n2935), .I4(n2936), .O(n2932)
         );
  NAND_GATE U3911 ( .I1(n2170), .I2(\registres[22][20] ), .O(n2936) );
  NAND_GATE U3912 ( .I1(n2171), .I2(\registres[15][20] ), .O(n2935) );
  NAND_GATE U3913 ( .I1(n2172), .I2(\registres[23][20] ), .O(n2934) );
  NAND_GATE U3914 ( .I1(n2173), .I2(\registres[4][20] ), .O(n2933) );
  NAND_GATE U3915 ( .I1(n2174), .I2(\registres[8][20] ), .O(n2931) );
  NAND_GATE U3916 ( .I1(n2175), .I2(\registres[2][20] ), .O(n2930) );
  NAND_GATE U3917 ( .I1(n2176), .I2(\registres[16][20] ), .O(n2929) );
  AND_GATE U3918 ( .I1(n2937), .I2(n2105), .O(data_src2[1]) );
  NAND4_GATE U3919 ( .I1(n2938), .I2(n2939), .I3(n2940), .I4(n2941), .O(n2937)
         );
  AND5_GATE U3920 ( .I1(n2942), .I2(n2943), .I3(n2944), .I4(n2945), .I5(n2946), 
        .O(n2941) );
  AND4_GATE U3921 ( .I1(n2947), .I2(n2948), .I3(n2949), .I4(n2950), .O(n2946)
         );
  NAND_GATE U3922 ( .I1(n2120), .I2(\registres[24][1] ), .O(n2950) );
  NAND_GATE U3923 ( .I1(n2121), .I2(\registres[25][1] ), .O(n2949) );
  NAND_GATE U3924 ( .I1(n2122), .I2(\registres[3][1] ), .O(n2948) );
  NAND_GATE U3925 ( .I1(n2123), .I2(\registres[26][1] ), .O(n2947) );
  NAND_GATE U3926 ( .I1(n2124), .I2(\registres[27][1] ), .O(n2945) );
  NAND_GATE U3927 ( .I1(n2125), .I2(\registres[10][1] ), .O(n2944) );
  NAND_GATE U3928 ( .I1(n2126), .I2(\registres[18][1] ), .O(n2943) );
  NAND_GATE U3929 ( .I1(n2127), .I2(\registres[5][1] ), .O(n2942) );
  AND5_GATE U3930 ( .I1(n2951), .I2(n2952), .I3(n2953), .I4(n2954), .I5(n2955), 
        .O(n2940) );
  AND4_GATE U3931 ( .I1(n2956), .I2(n2957), .I3(n2958), .I4(n2959), .O(n2955)
         );
  NAND_GATE U3932 ( .I1(n2137), .I2(\registres[28][1] ), .O(n2959) );
  NAND_GATE U3933 ( .I1(n2138), .I2(\registres[29][1] ), .O(n2958) );
  NAND_GATE U3934 ( .I1(n2139), .I2(\registres[12][1] ), .O(n2957) );
  NAND_GATE U3935 ( .I1(n2140), .I2(\registres[20][1] ), .O(n2956) );
  NAND_GATE U3936 ( .I1(n2141), .I2(\registres[1][1] ), .O(n2954) );
  NAND_GATE U3937 ( .I1(n2142), .I2(\registres[9][1] ), .O(n2953) );
  NAND_GATE U3938 ( .I1(n2143), .I2(\registres[11][1] ), .O(n2952) );
  NAND_GATE U3939 ( .I1(n2144), .I2(\registres[13][1] ), .O(n2951) );
  AND5_GATE U3940 ( .I1(n2960), .I2(n2961), .I3(n2962), .I4(n2963), .I5(n2964), 
        .O(n2939) );
  AND4_GATE U3941 ( .I1(n2965), .I2(n2966), .I3(n2967), .I4(n2968), .O(n2964)
         );
  NAND_GATE U3942 ( .I1(n2154), .I2(\registres[17][1] ), .O(n2968) );
  NAND_GATE U3943 ( .I1(n2155), .I2(\registres[19][1] ), .O(n2967) );
  NAND_GATE U3944 ( .I1(n2156), .I2(\registres[21][1] ), .O(n2966) );
  NAND_GATE U3945 ( .I1(n2157), .I2(\registres[6][1] ), .O(n2965) );
  NAND_GATE U3946 ( .I1(n2158), .I2(\registres[7][1] ), .O(n2963) );
  NAND_GATE U3947 ( .I1(n2159), .I2(\registres[30][1] ), .O(n2962) );
  NAND_GATE U3948 ( .I1(n2160), .I2(\registres[31][1] ), .O(n2961) );
  NAND_GATE U3949 ( .I1(n2161), .I2(\registres[14][1] ), .O(n2960) );
  AND4_GATE U3950 ( .I1(n2969), .I2(n2970), .I3(n2971), .I4(n2972), .O(n2938)
         );
  AND4_GATE U3951 ( .I1(n2973), .I2(n2974), .I3(n2975), .I4(n2976), .O(n2972)
         );
  NAND_GATE U3952 ( .I1(n2170), .I2(\registres[22][1] ), .O(n2976) );
  NAND_GATE U3953 ( .I1(n2171), .I2(\registres[15][1] ), .O(n2975) );
  NAND_GATE U3954 ( .I1(n2172), .I2(\registres[23][1] ), .O(n2974) );
  NAND_GATE U3955 ( .I1(n2173), .I2(\registres[4][1] ), .O(n2973) );
  NAND_GATE U3956 ( .I1(n2174), .I2(\registres[8][1] ), .O(n2971) );
  NAND_GATE U3957 ( .I1(n2175), .I2(\registres[2][1] ), .O(n2970) );
  NAND_GATE U3958 ( .I1(n2176), .I2(\registres[16][1] ), .O(n2969) );
  AND_GATE U3959 ( .I1(n2977), .I2(n2105), .O(data_src2[19]) );
  NAND4_GATE U3960 ( .I1(n2978), .I2(n2979), .I3(n2980), .I4(n2981), .O(n2977)
         );
  AND5_GATE U3961 ( .I1(n2982), .I2(n2983), .I3(n2984), .I4(n2985), .I5(n2986), 
        .O(n2981) );
  AND4_GATE U3962 ( .I1(n2987), .I2(n2988), .I3(n2989), .I4(n2990), .O(n2986)
         );
  NAND_GATE U3963 ( .I1(n2120), .I2(\registres[24][19] ), .O(n2990) );
  NAND_GATE U3964 ( .I1(n2121), .I2(\registres[25][19] ), .O(n2989) );
  NAND_GATE U3965 ( .I1(n2122), .I2(\registres[3][19] ), .O(n2988) );
  NAND_GATE U3966 ( .I1(n2123), .I2(\registres[26][19] ), .O(n2987) );
  NAND_GATE U3967 ( .I1(n2124), .I2(\registres[27][19] ), .O(n2985) );
  NAND_GATE U3968 ( .I1(n2125), .I2(\registres[10][19] ), .O(n2984) );
  NAND_GATE U3969 ( .I1(n2126), .I2(\registres[18][19] ), .O(n2983) );
  NAND_GATE U3970 ( .I1(n2127), .I2(\registres[5][19] ), .O(n2982) );
  AND5_GATE U3971 ( .I1(n2991), .I2(n2992), .I3(n2993), .I4(n2994), .I5(n2995), 
        .O(n2980) );
  AND4_GATE U3972 ( .I1(n2996), .I2(n2997), .I3(n2998), .I4(n2999), .O(n2995)
         );
  NAND_GATE U3973 ( .I1(n2137), .I2(\registres[28][19] ), .O(n2999) );
  NAND_GATE U3974 ( .I1(n2138), .I2(\registres[29][19] ), .O(n2998) );
  NAND_GATE U3975 ( .I1(n2139), .I2(\registres[12][19] ), .O(n2997) );
  NAND_GATE U3976 ( .I1(n2140), .I2(\registres[20][19] ), .O(n2996) );
  NAND_GATE U3977 ( .I1(n2141), .I2(\registres[1][19] ), .O(n2994) );
  NAND_GATE U3978 ( .I1(n2142), .I2(\registres[9][19] ), .O(n2993) );
  NAND_GATE U3979 ( .I1(n2143), .I2(\registres[11][19] ), .O(n2992) );
  NAND_GATE U3980 ( .I1(n2144), .I2(\registres[13][19] ), .O(n2991) );
  AND5_GATE U3981 ( .I1(n3000), .I2(n3001), .I3(n3002), .I4(n3003), .I5(n3004), 
        .O(n2979) );
  AND4_GATE U3982 ( .I1(n3005), .I2(n3006), .I3(n3007), .I4(n3008), .O(n3004)
         );
  NAND_GATE U3983 ( .I1(n2154), .I2(\registres[17][19] ), .O(n3008) );
  NAND_GATE U3984 ( .I1(n2155), .I2(\registres[19][19] ), .O(n3007) );
  NAND_GATE U3985 ( .I1(n2156), .I2(\registres[21][19] ), .O(n3006) );
  NAND_GATE U3986 ( .I1(n2157), .I2(\registres[6][19] ), .O(n3005) );
  NAND_GATE U3987 ( .I1(n2158), .I2(\registres[7][19] ), .O(n3003) );
  NAND_GATE U3988 ( .I1(n2159), .I2(\registres[30][19] ), .O(n3002) );
  NAND_GATE U3989 ( .I1(n2160), .I2(\registres[31][19] ), .O(n3001) );
  NAND_GATE U3990 ( .I1(n2161), .I2(\registres[14][19] ), .O(n3000) );
  AND4_GATE U3991 ( .I1(n3009), .I2(n3010), .I3(n3011), .I4(n3012), .O(n2978)
         );
  AND4_GATE U3992 ( .I1(n3013), .I2(n3014), .I3(n3015), .I4(n3016), .O(n3012)
         );
  NAND_GATE U3993 ( .I1(n2170), .I2(\registres[22][19] ), .O(n3016) );
  NAND_GATE U3994 ( .I1(n2171), .I2(\registres[15][19] ), .O(n3015) );
  NAND_GATE U3995 ( .I1(n2172), .I2(\registres[23][19] ), .O(n3014) );
  NAND_GATE U3996 ( .I1(n2173), .I2(\registres[4][19] ), .O(n3013) );
  NAND_GATE U3997 ( .I1(n2174), .I2(\registres[8][19] ), .O(n3011) );
  NAND_GATE U3998 ( .I1(n2175), .I2(\registres[2][19] ), .O(n3010) );
  NAND_GATE U3999 ( .I1(n2176), .I2(\registres[16][19] ), .O(n3009) );
  AND_GATE U4000 ( .I1(n3017), .I2(n2105), .O(data_src2[18]) );
  NAND4_GATE U4001 ( .I1(n3018), .I2(n3019), .I3(n3020), .I4(n3021), .O(n3017)
         );
  AND5_GATE U4002 ( .I1(n3022), .I2(n3023), .I3(n3024), .I4(n3025), .I5(n3026), 
        .O(n3021) );
  AND4_GATE U4003 ( .I1(n3027), .I2(n3028), .I3(n3029), .I4(n3030), .O(n3026)
         );
  NAND_GATE U4004 ( .I1(n2120), .I2(\registres[24][18] ), .O(n3030) );
  NAND_GATE U4005 ( .I1(n2121), .I2(\registres[25][18] ), .O(n3029) );
  NAND_GATE U4006 ( .I1(n2122), .I2(\registres[3][18] ), .O(n3028) );
  NAND_GATE U4007 ( .I1(n2123), .I2(\registres[26][18] ), .O(n3027) );
  NAND_GATE U4008 ( .I1(n2124), .I2(\registres[27][18] ), .O(n3025) );
  NAND_GATE U4009 ( .I1(n2125), .I2(\registres[10][18] ), .O(n3024) );
  NAND_GATE U4010 ( .I1(n2126), .I2(\registres[18][18] ), .O(n3023) );
  NAND_GATE U4011 ( .I1(n2127), .I2(\registres[5][18] ), .O(n3022) );
  AND5_GATE U4012 ( .I1(n3031), .I2(n3032), .I3(n3033), .I4(n3034), .I5(n3035), 
        .O(n3020) );
  AND4_GATE U4013 ( .I1(n3036), .I2(n3037), .I3(n3038), .I4(n3039), .O(n3035)
         );
  NAND_GATE U4014 ( .I1(n2137), .I2(\registres[28][18] ), .O(n3039) );
  NAND_GATE U4015 ( .I1(n2138), .I2(\registres[29][18] ), .O(n3038) );
  NAND_GATE U4016 ( .I1(n2139), .I2(\registres[12][18] ), .O(n3037) );
  NAND_GATE U4017 ( .I1(n2140), .I2(\registres[20][18] ), .O(n3036) );
  NAND_GATE U4018 ( .I1(n2141), .I2(\registres[1][18] ), .O(n3034) );
  NAND_GATE U4019 ( .I1(n2142), .I2(\registres[9][18] ), .O(n3033) );
  NAND_GATE U4020 ( .I1(n2143), .I2(\registres[11][18] ), .O(n3032) );
  NAND_GATE U4021 ( .I1(n2144), .I2(\registres[13][18] ), .O(n3031) );
  AND5_GATE U4022 ( .I1(n3040), .I2(n3041), .I3(n3042), .I4(n3043), .I5(n3044), 
        .O(n3019) );
  AND4_GATE U4023 ( .I1(n3045), .I2(n3046), .I3(n3047), .I4(n3048), .O(n3044)
         );
  NAND_GATE U4024 ( .I1(n2154), .I2(\registres[17][18] ), .O(n3048) );
  NAND_GATE U4025 ( .I1(n2155), .I2(\registres[19][18] ), .O(n3047) );
  NAND_GATE U4026 ( .I1(n2156), .I2(\registres[21][18] ), .O(n3046) );
  NAND_GATE U4027 ( .I1(n2157), .I2(\registres[6][18] ), .O(n3045) );
  NAND_GATE U4028 ( .I1(n2158), .I2(\registres[7][18] ), .O(n3043) );
  NAND_GATE U4029 ( .I1(n2159), .I2(\registres[30][18] ), .O(n3042) );
  NAND_GATE U4030 ( .I1(n2160), .I2(\registres[31][18] ), .O(n3041) );
  NAND_GATE U4031 ( .I1(n2161), .I2(\registres[14][18] ), .O(n3040) );
  AND4_GATE U4032 ( .I1(n3049), .I2(n3050), .I3(n3051), .I4(n3052), .O(n3018)
         );
  AND4_GATE U4033 ( .I1(n3053), .I2(n3054), .I3(n3055), .I4(n3056), .O(n3052)
         );
  NAND_GATE U4034 ( .I1(n2170), .I2(\registres[22][18] ), .O(n3056) );
  NAND_GATE U4035 ( .I1(n2171), .I2(\registres[15][18] ), .O(n3055) );
  NAND_GATE U4036 ( .I1(n2172), .I2(\registres[23][18] ), .O(n3054) );
  NAND_GATE U4037 ( .I1(n2173), .I2(\registres[4][18] ), .O(n3053) );
  NAND_GATE U4038 ( .I1(n2174), .I2(\registres[8][18] ), .O(n3051) );
  NAND_GATE U4039 ( .I1(n2175), .I2(\registres[2][18] ), .O(n3050) );
  NAND_GATE U4040 ( .I1(n2176), .I2(\registres[16][18] ), .O(n3049) );
  AND_GATE U4041 ( .I1(n3057), .I2(n2105), .O(data_src2[17]) );
  NAND4_GATE U4042 ( .I1(n3058), .I2(n3059), .I3(n3060), .I4(n3061), .O(n3057)
         );
  AND5_GATE U4043 ( .I1(n3062), .I2(n3063), .I3(n3064), .I4(n3065), .I5(n3066), 
        .O(n3061) );
  AND4_GATE U4044 ( .I1(n3067), .I2(n3068), .I3(n3069), .I4(n3070), .O(n3066)
         );
  NAND_GATE U4045 ( .I1(n2120), .I2(\registres[24][17] ), .O(n3070) );
  NAND_GATE U4046 ( .I1(n2121), .I2(\registres[25][17] ), .O(n3069) );
  NAND_GATE U4047 ( .I1(n2122), .I2(\registres[3][17] ), .O(n3068) );
  NAND_GATE U4048 ( .I1(n2123), .I2(\registres[26][17] ), .O(n3067) );
  NAND_GATE U4049 ( .I1(n2124), .I2(\registres[27][17] ), .O(n3065) );
  NAND_GATE U4050 ( .I1(n2125), .I2(\registres[10][17] ), .O(n3064) );
  NAND_GATE U4051 ( .I1(n2126), .I2(\registres[18][17] ), .O(n3063) );
  NAND_GATE U4052 ( .I1(n2127), .I2(\registres[5][17] ), .O(n3062) );
  AND5_GATE U4053 ( .I1(n3071), .I2(n3072), .I3(n3073), .I4(n3074), .I5(n3075), 
        .O(n3060) );
  AND4_GATE U4054 ( .I1(n3076), .I2(n3077), .I3(n3078), .I4(n3079), .O(n3075)
         );
  NAND_GATE U4055 ( .I1(n2137), .I2(\registres[28][17] ), .O(n3079) );
  NAND_GATE U4056 ( .I1(n2138), .I2(\registres[29][17] ), .O(n3078) );
  NAND_GATE U4057 ( .I1(n2139), .I2(\registres[12][17] ), .O(n3077) );
  NAND_GATE U4058 ( .I1(n2140), .I2(\registres[20][17] ), .O(n3076) );
  NAND_GATE U4059 ( .I1(n2141), .I2(\registres[1][17] ), .O(n3074) );
  NAND_GATE U4060 ( .I1(n2142), .I2(\registres[9][17] ), .O(n3073) );
  NAND_GATE U4061 ( .I1(n2143), .I2(\registres[11][17] ), .O(n3072) );
  NAND_GATE U4062 ( .I1(n2144), .I2(\registres[13][17] ), .O(n3071) );
  AND5_GATE U4063 ( .I1(n3080), .I2(n3081), .I3(n3082), .I4(n3083), .I5(n3084), 
        .O(n3059) );
  AND4_GATE U4064 ( .I1(n3085), .I2(n3086), .I3(n3087), .I4(n3088), .O(n3084)
         );
  NAND_GATE U4065 ( .I1(n2154), .I2(\registres[17][17] ), .O(n3088) );
  NAND_GATE U4066 ( .I1(n2155), .I2(\registres[19][17] ), .O(n3087) );
  NAND_GATE U4067 ( .I1(n2156), .I2(\registres[21][17] ), .O(n3086) );
  NAND_GATE U4068 ( .I1(n2157), .I2(\registres[6][17] ), .O(n3085) );
  NAND_GATE U4069 ( .I1(n2158), .I2(\registres[7][17] ), .O(n3083) );
  NAND_GATE U4070 ( .I1(n2159), .I2(\registres[30][17] ), .O(n3082) );
  NAND_GATE U4071 ( .I1(n2160), .I2(\registres[31][17] ), .O(n3081) );
  NAND_GATE U4072 ( .I1(n2161), .I2(\registres[14][17] ), .O(n3080) );
  AND4_GATE U4073 ( .I1(n3089), .I2(n3090), .I3(n3091), .I4(n3092), .O(n3058)
         );
  AND4_GATE U4074 ( .I1(n3093), .I2(n3094), .I3(n3095), .I4(n3096), .O(n3092)
         );
  NAND_GATE U4075 ( .I1(n2170), .I2(\registres[22][17] ), .O(n3096) );
  NAND_GATE U4076 ( .I1(n2171), .I2(\registres[15][17] ), .O(n3095) );
  NAND_GATE U4077 ( .I1(n2172), .I2(\registres[23][17] ), .O(n3094) );
  NAND_GATE U4078 ( .I1(n2173), .I2(\registres[4][17] ), .O(n3093) );
  NAND_GATE U4079 ( .I1(n2174), .I2(\registres[8][17] ), .O(n3091) );
  NAND_GATE U4080 ( .I1(n2175), .I2(\registres[2][17] ), .O(n3090) );
  NAND_GATE U4081 ( .I1(n2176), .I2(\registres[16][17] ), .O(n3089) );
  AND_GATE U4082 ( .I1(n3097), .I2(n2105), .O(data_src2[16]) );
  NAND4_GATE U4083 ( .I1(n3098), .I2(n3099), .I3(n3100), .I4(n3101), .O(n3097)
         );
  AND5_GATE U4084 ( .I1(n3102), .I2(n3103), .I3(n3104), .I4(n3105), .I5(n3106), 
        .O(n3101) );
  AND4_GATE U4085 ( .I1(n3107), .I2(n3108), .I3(n3109), .I4(n3110), .O(n3106)
         );
  NAND_GATE U4086 ( .I1(n2120), .I2(\registres[24][16] ), .O(n3110) );
  NAND_GATE U4087 ( .I1(n2121), .I2(\registres[25][16] ), .O(n3109) );
  NAND_GATE U4088 ( .I1(n2122), .I2(\registres[3][16] ), .O(n3108) );
  NAND_GATE U4089 ( .I1(n2123), .I2(\registres[26][16] ), .O(n3107) );
  NAND_GATE U4090 ( .I1(n2124), .I2(\registres[27][16] ), .O(n3105) );
  NAND_GATE U4091 ( .I1(n2125), .I2(\registres[10][16] ), .O(n3104) );
  NAND_GATE U4092 ( .I1(n2126), .I2(\registres[18][16] ), .O(n3103) );
  NAND_GATE U4093 ( .I1(n2127), .I2(\registres[5][16] ), .O(n3102) );
  AND5_GATE U4094 ( .I1(n3111), .I2(n3112), .I3(n3113), .I4(n3114), .I5(n3115), 
        .O(n3100) );
  AND4_GATE U4095 ( .I1(n3116), .I2(n3117), .I3(n3118), .I4(n3119), .O(n3115)
         );
  NAND_GATE U4096 ( .I1(n2137), .I2(\registres[28][16] ), .O(n3119) );
  NAND_GATE U4097 ( .I1(n2138), .I2(\registres[29][16] ), .O(n3118) );
  NAND_GATE U4098 ( .I1(n2139), .I2(\registres[12][16] ), .O(n3117) );
  NAND_GATE U4099 ( .I1(n2140), .I2(\registres[20][16] ), .O(n3116) );
  NAND_GATE U4100 ( .I1(n2141), .I2(\registres[1][16] ), .O(n3114) );
  NAND_GATE U4101 ( .I1(n2142), .I2(\registres[9][16] ), .O(n3113) );
  NAND_GATE U4102 ( .I1(n2143), .I2(\registres[11][16] ), .O(n3112) );
  NAND_GATE U4103 ( .I1(n2144), .I2(\registres[13][16] ), .O(n3111) );
  AND5_GATE U4104 ( .I1(n3120), .I2(n3121), .I3(n3122), .I4(n3123), .I5(n3124), 
        .O(n3099) );
  AND4_GATE U4105 ( .I1(n3125), .I2(n3126), .I3(n3127), .I4(n3128), .O(n3124)
         );
  NAND_GATE U4106 ( .I1(n2154), .I2(\registres[17][16] ), .O(n3128) );
  NAND_GATE U4107 ( .I1(n2155), .I2(\registres[19][16] ), .O(n3127) );
  NAND_GATE U4108 ( .I1(n2156), .I2(\registres[21][16] ), .O(n3126) );
  NAND_GATE U4109 ( .I1(n2157), .I2(\registres[6][16] ), .O(n3125) );
  NAND_GATE U4110 ( .I1(n2158), .I2(\registres[7][16] ), .O(n3123) );
  NAND_GATE U4111 ( .I1(n2159), .I2(\registres[30][16] ), .O(n3122) );
  NAND_GATE U4112 ( .I1(n2160), .I2(\registres[31][16] ), .O(n3121) );
  NAND_GATE U4113 ( .I1(n2161), .I2(\registres[14][16] ), .O(n3120) );
  AND4_GATE U4114 ( .I1(n3129), .I2(n3130), .I3(n3131), .I4(n3132), .O(n3098)
         );
  AND4_GATE U4115 ( .I1(n3133), .I2(n3134), .I3(n3135), .I4(n3136), .O(n3132)
         );
  NAND_GATE U4116 ( .I1(n2170), .I2(\registres[22][16] ), .O(n3136) );
  NAND_GATE U4117 ( .I1(n2171), .I2(\registres[15][16] ), .O(n3135) );
  NAND_GATE U4118 ( .I1(n2172), .I2(\registres[23][16] ), .O(n3134) );
  NAND_GATE U4119 ( .I1(n2173), .I2(\registres[4][16] ), .O(n3133) );
  NAND_GATE U4120 ( .I1(n2174), .I2(\registres[8][16] ), .O(n3131) );
  NAND_GATE U4121 ( .I1(n2175), .I2(\registres[2][16] ), .O(n3130) );
  NAND_GATE U4122 ( .I1(n2176), .I2(\registres[16][16] ), .O(n3129) );
  AND_GATE U4123 ( .I1(n3137), .I2(n2105), .O(data_src2[15]) );
  NAND4_GATE U4124 ( .I1(n3138), .I2(n3139), .I3(n3140), .I4(n3141), .O(n3137)
         );
  AND5_GATE U4125 ( .I1(n3142), .I2(n3143), .I3(n3144), .I4(n3145), .I5(n3146), 
        .O(n3141) );
  AND4_GATE U4126 ( .I1(n3147), .I2(n3148), .I3(n3149), .I4(n3150), .O(n3146)
         );
  NAND_GATE U4127 ( .I1(n2120), .I2(\registres[24][15] ), .O(n3150) );
  NAND_GATE U4128 ( .I1(n2121), .I2(\registres[25][15] ), .O(n3149) );
  NAND_GATE U4129 ( .I1(n2122), .I2(\registres[3][15] ), .O(n3148) );
  NAND_GATE U4130 ( .I1(n2123), .I2(\registres[26][15] ), .O(n3147) );
  NAND_GATE U4131 ( .I1(n2124), .I2(\registres[27][15] ), .O(n3145) );
  NAND_GATE U4132 ( .I1(n2125), .I2(\registres[10][15] ), .O(n3144) );
  NAND_GATE U4133 ( .I1(n2126), .I2(\registres[18][15] ), .O(n3143) );
  NAND_GATE U4134 ( .I1(n2127), .I2(\registres[5][15] ), .O(n3142) );
  AND5_GATE U4135 ( .I1(n3151), .I2(n3152), .I3(n3153), .I4(n3154), .I5(n3155), 
        .O(n3140) );
  AND4_GATE U4136 ( .I1(n3156), .I2(n3157), .I3(n3158), .I4(n3159), .O(n3155)
         );
  NAND_GATE U4137 ( .I1(n2137), .I2(\registres[28][15] ), .O(n3159) );
  NAND_GATE U4138 ( .I1(n2138), .I2(\registres[29][15] ), .O(n3158) );
  NAND_GATE U4139 ( .I1(n2139), .I2(\registres[12][15] ), .O(n3157) );
  NAND_GATE U4140 ( .I1(n2140), .I2(\registres[20][15] ), .O(n3156) );
  NAND_GATE U4141 ( .I1(n2141), .I2(\registres[1][15] ), .O(n3154) );
  NAND_GATE U4142 ( .I1(n2142), .I2(\registres[9][15] ), .O(n3153) );
  NAND_GATE U4143 ( .I1(n2143), .I2(\registres[11][15] ), .O(n3152) );
  NAND_GATE U4144 ( .I1(n2144), .I2(\registres[13][15] ), .O(n3151) );
  AND5_GATE U4145 ( .I1(n3160), .I2(n3161), .I3(n3162), .I4(n3163), .I5(n3164), 
        .O(n3139) );
  AND4_GATE U4146 ( .I1(n3165), .I2(n3166), .I3(n3167), .I4(n3168), .O(n3164)
         );
  NAND_GATE U4147 ( .I1(n2154), .I2(\registres[17][15] ), .O(n3168) );
  NAND_GATE U4148 ( .I1(n2155), .I2(\registres[19][15] ), .O(n3167) );
  NAND_GATE U4149 ( .I1(n2156), .I2(\registres[21][15] ), .O(n3166) );
  NAND_GATE U4150 ( .I1(n2157), .I2(\registres[6][15] ), .O(n3165) );
  NAND_GATE U4151 ( .I1(n2158), .I2(\registres[7][15] ), .O(n3163) );
  NAND_GATE U4152 ( .I1(n2159), .I2(\registres[30][15] ), .O(n3162) );
  NAND_GATE U4153 ( .I1(n2160), .I2(\registres[31][15] ), .O(n3161) );
  NAND_GATE U4154 ( .I1(n2161), .I2(\registres[14][15] ), .O(n3160) );
  AND4_GATE U4155 ( .I1(n3169), .I2(n3170), .I3(n3171), .I4(n3172), .O(n3138)
         );
  AND4_GATE U4156 ( .I1(n3173), .I2(n3174), .I3(n3175), .I4(n3176), .O(n3172)
         );
  NAND_GATE U4157 ( .I1(n2170), .I2(\registres[22][15] ), .O(n3176) );
  NAND_GATE U4158 ( .I1(n2171), .I2(\registres[15][15] ), .O(n3175) );
  NAND_GATE U4159 ( .I1(n2172), .I2(\registres[23][15] ), .O(n3174) );
  NAND_GATE U4160 ( .I1(n2173), .I2(\registres[4][15] ), .O(n3173) );
  NAND_GATE U4161 ( .I1(n2174), .I2(\registres[8][15] ), .O(n3171) );
  NAND_GATE U4162 ( .I1(n2175), .I2(\registres[2][15] ), .O(n3170) );
  NAND_GATE U4163 ( .I1(n2176), .I2(\registres[16][15] ), .O(n3169) );
  AND_GATE U4164 ( .I1(n3177), .I2(n2105), .O(data_src2[14]) );
  NAND4_GATE U4165 ( .I1(n3178), .I2(n3179), .I3(n3180), .I4(n3181), .O(n3177)
         );
  AND5_GATE U4166 ( .I1(n3182), .I2(n3183), .I3(n3184), .I4(n3185), .I5(n3186), 
        .O(n3181) );
  AND4_GATE U4167 ( .I1(n3187), .I2(n3188), .I3(n3189), .I4(n3190), .O(n3186)
         );
  NAND_GATE U4168 ( .I1(n2120), .I2(\registres[24][14] ), .O(n3190) );
  NAND_GATE U4169 ( .I1(n2121), .I2(\registres[25][14] ), .O(n3189) );
  NAND_GATE U4170 ( .I1(n2122), .I2(\registres[3][14] ), .O(n3188) );
  NAND_GATE U4171 ( .I1(n2123), .I2(\registres[26][14] ), .O(n3187) );
  NAND_GATE U4172 ( .I1(n2124), .I2(\registres[27][14] ), .O(n3185) );
  NAND_GATE U4173 ( .I1(n2125), .I2(\registres[10][14] ), .O(n3184) );
  NAND_GATE U4174 ( .I1(n2126), .I2(\registres[18][14] ), .O(n3183) );
  NAND_GATE U4175 ( .I1(n2127), .I2(\registres[5][14] ), .O(n3182) );
  AND5_GATE U4176 ( .I1(n3191), .I2(n3192), .I3(n3193), .I4(n3194), .I5(n3195), 
        .O(n3180) );
  AND4_GATE U4177 ( .I1(n3196), .I2(n3197), .I3(n3198), .I4(n3199), .O(n3195)
         );
  NAND_GATE U4178 ( .I1(n2137), .I2(\registres[28][14] ), .O(n3199) );
  NAND_GATE U4179 ( .I1(n2138), .I2(\registres[29][14] ), .O(n3198) );
  NAND_GATE U4180 ( .I1(n2139), .I2(\registres[12][14] ), .O(n3197) );
  NAND_GATE U4181 ( .I1(n2140), .I2(\registres[20][14] ), .O(n3196) );
  NAND_GATE U4182 ( .I1(n2141), .I2(\registres[1][14] ), .O(n3194) );
  NAND_GATE U4183 ( .I1(n2142), .I2(\registres[9][14] ), .O(n3193) );
  NAND_GATE U4184 ( .I1(n2143), .I2(\registres[11][14] ), .O(n3192) );
  NAND_GATE U4185 ( .I1(n2144), .I2(\registres[13][14] ), .O(n3191) );
  AND5_GATE U4186 ( .I1(n3200), .I2(n3201), .I3(n3202), .I4(n3203), .I5(n3204), 
        .O(n3179) );
  AND4_GATE U4187 ( .I1(n3205), .I2(n3206), .I3(n3207), .I4(n3208), .O(n3204)
         );
  NAND_GATE U4188 ( .I1(n2154), .I2(\registres[17][14] ), .O(n3208) );
  NAND_GATE U4189 ( .I1(n2155), .I2(\registres[19][14] ), .O(n3207) );
  NAND_GATE U4190 ( .I1(n2156), .I2(\registres[21][14] ), .O(n3206) );
  NAND_GATE U4191 ( .I1(n2157), .I2(\registres[6][14] ), .O(n3205) );
  NAND_GATE U4192 ( .I1(n2158), .I2(\registres[7][14] ), .O(n3203) );
  NAND_GATE U4193 ( .I1(n2159), .I2(\registres[30][14] ), .O(n3202) );
  NAND_GATE U4194 ( .I1(n2160), .I2(\registres[31][14] ), .O(n3201) );
  NAND_GATE U4195 ( .I1(n2161), .I2(\registres[14][14] ), .O(n3200) );
  AND4_GATE U4196 ( .I1(n3209), .I2(n3210), .I3(n3211), .I4(n3212), .O(n3178)
         );
  AND4_GATE U4197 ( .I1(n3213), .I2(n3214), .I3(n3215), .I4(n3216), .O(n3212)
         );
  NAND_GATE U4198 ( .I1(n2170), .I2(\registres[22][14] ), .O(n3216) );
  NAND_GATE U4199 ( .I1(n2171), .I2(\registres[15][14] ), .O(n3215) );
  NAND_GATE U4200 ( .I1(n2172), .I2(\registres[23][14] ), .O(n3214) );
  NAND_GATE U4201 ( .I1(n2173), .I2(\registres[4][14] ), .O(n3213) );
  NAND_GATE U4202 ( .I1(n2174), .I2(\registres[8][14] ), .O(n3211) );
  NAND_GATE U4203 ( .I1(n2175), .I2(\registres[2][14] ), .O(n3210) );
  NAND_GATE U4204 ( .I1(n2176), .I2(\registres[16][14] ), .O(n3209) );
  AND_GATE U4205 ( .I1(n3217), .I2(n2105), .O(data_src2[13]) );
  NAND4_GATE U4206 ( .I1(n3218), .I2(n3219), .I3(n3220), .I4(n3221), .O(n3217)
         );
  AND5_GATE U4207 ( .I1(n3222), .I2(n3223), .I3(n3224), .I4(n3225), .I5(n3226), 
        .O(n3221) );
  AND4_GATE U4208 ( .I1(n3227), .I2(n3228), .I3(n3229), .I4(n3230), .O(n3226)
         );
  NAND_GATE U4209 ( .I1(n2120), .I2(\registres[24][13] ), .O(n3230) );
  NAND_GATE U4210 ( .I1(n2121), .I2(\registres[25][13] ), .O(n3229) );
  NAND_GATE U4211 ( .I1(n2122), .I2(\registres[3][13] ), .O(n3228) );
  NAND_GATE U4212 ( .I1(n2123), .I2(\registres[26][13] ), .O(n3227) );
  NAND_GATE U4213 ( .I1(n2124), .I2(\registres[27][13] ), .O(n3225) );
  NAND_GATE U4214 ( .I1(n2125), .I2(\registres[10][13] ), .O(n3224) );
  NAND_GATE U4215 ( .I1(n2126), .I2(\registres[18][13] ), .O(n3223) );
  NAND_GATE U4216 ( .I1(n2127), .I2(\registres[5][13] ), .O(n3222) );
  AND5_GATE U4217 ( .I1(n3231), .I2(n3232), .I3(n3233), .I4(n3234), .I5(n3235), 
        .O(n3220) );
  AND4_GATE U4218 ( .I1(n3236), .I2(n3237), .I3(n3238), .I4(n3239), .O(n3235)
         );
  NAND_GATE U4219 ( .I1(n2137), .I2(\registres[28][13] ), .O(n3239) );
  NAND_GATE U4220 ( .I1(n2138), .I2(\registres[29][13] ), .O(n3238) );
  NAND_GATE U4221 ( .I1(n2139), .I2(\registres[12][13] ), .O(n3237) );
  NAND_GATE U4222 ( .I1(n2140), .I2(\registres[20][13] ), .O(n3236) );
  NAND_GATE U4223 ( .I1(n2141), .I2(\registres[1][13] ), .O(n3234) );
  NAND_GATE U4224 ( .I1(n2142), .I2(\registres[9][13] ), .O(n3233) );
  NAND_GATE U4225 ( .I1(n2143), .I2(\registres[11][13] ), .O(n3232) );
  NAND_GATE U4226 ( .I1(n2144), .I2(\registres[13][13] ), .O(n3231) );
  AND5_GATE U4227 ( .I1(n3240), .I2(n3241), .I3(n3242), .I4(n3243), .I5(n3244), 
        .O(n3219) );
  AND4_GATE U4228 ( .I1(n3245), .I2(n3246), .I3(n3247), .I4(n3248), .O(n3244)
         );
  NAND_GATE U4229 ( .I1(n2154), .I2(\registres[17][13] ), .O(n3248) );
  NAND_GATE U4230 ( .I1(n2155), .I2(\registres[19][13] ), .O(n3247) );
  NAND_GATE U4231 ( .I1(n2156), .I2(\registres[21][13] ), .O(n3246) );
  NAND_GATE U4232 ( .I1(n2157), .I2(\registres[6][13] ), .O(n3245) );
  NAND_GATE U4233 ( .I1(n2158), .I2(\registres[7][13] ), .O(n3243) );
  NAND_GATE U4234 ( .I1(n2159), .I2(\registres[30][13] ), .O(n3242) );
  NAND_GATE U4235 ( .I1(n2160), .I2(\registres[31][13] ), .O(n3241) );
  NAND_GATE U4236 ( .I1(n2161), .I2(\registres[14][13] ), .O(n3240) );
  AND4_GATE U4237 ( .I1(n3249), .I2(n3250), .I3(n3251), .I4(n3252), .O(n3218)
         );
  AND4_GATE U4238 ( .I1(n3253), .I2(n3254), .I3(n3255), .I4(n3256), .O(n3252)
         );
  NAND_GATE U4239 ( .I1(n2170), .I2(\registres[22][13] ), .O(n3256) );
  NAND_GATE U4240 ( .I1(n2171), .I2(\registres[15][13] ), .O(n3255) );
  NAND_GATE U4241 ( .I1(n2172), .I2(\registres[23][13] ), .O(n3254) );
  NAND_GATE U4242 ( .I1(n2173), .I2(\registres[4][13] ), .O(n3253) );
  NAND_GATE U4243 ( .I1(n2174), .I2(\registres[8][13] ), .O(n3251) );
  NAND_GATE U4244 ( .I1(n2175), .I2(\registres[2][13] ), .O(n3250) );
  NAND_GATE U4245 ( .I1(n2176), .I2(\registres[16][13] ), .O(n3249) );
  AND_GATE U4246 ( .I1(n3257), .I2(n2105), .O(data_src2[12]) );
  NAND4_GATE U4247 ( .I1(n3258), .I2(n3259), .I3(n3260), .I4(n3261), .O(n3257)
         );
  AND5_GATE U4248 ( .I1(n3262), .I2(n3263), .I3(n3264), .I4(n3265), .I5(n3266), 
        .O(n3261) );
  AND4_GATE U4249 ( .I1(n3267), .I2(n3268), .I3(n3269), .I4(n3270), .O(n3266)
         );
  NAND_GATE U4250 ( .I1(n2120), .I2(\registres[24][12] ), .O(n3270) );
  NAND_GATE U4251 ( .I1(n2121), .I2(\registres[25][12] ), .O(n3269) );
  NAND_GATE U4252 ( .I1(n2122), .I2(\registres[3][12] ), .O(n3268) );
  NAND_GATE U4253 ( .I1(n2123), .I2(\registres[26][12] ), .O(n3267) );
  NAND_GATE U4254 ( .I1(n2124), .I2(\registres[27][12] ), .O(n3265) );
  NAND_GATE U4255 ( .I1(n2125), .I2(\registres[10][12] ), .O(n3264) );
  NAND_GATE U4256 ( .I1(n2126), .I2(\registres[18][12] ), .O(n3263) );
  NAND_GATE U4257 ( .I1(n2127), .I2(\registres[5][12] ), .O(n3262) );
  AND5_GATE U4258 ( .I1(n3271), .I2(n3272), .I3(n3273), .I4(n3274), .I5(n3275), 
        .O(n3260) );
  AND4_GATE U4259 ( .I1(n3276), .I2(n3277), .I3(n3278), .I4(n3279), .O(n3275)
         );
  NAND_GATE U4260 ( .I1(n2137), .I2(\registres[28][12] ), .O(n3279) );
  NAND_GATE U4261 ( .I1(n2138), .I2(\registres[29][12] ), .O(n3278) );
  NAND_GATE U4262 ( .I1(n2139), .I2(\registres[12][12] ), .O(n3277) );
  NAND_GATE U4263 ( .I1(n2140), .I2(\registres[20][12] ), .O(n3276) );
  NAND_GATE U4264 ( .I1(n2141), .I2(\registres[1][12] ), .O(n3274) );
  NAND_GATE U4265 ( .I1(n2142), .I2(\registres[9][12] ), .O(n3273) );
  NAND_GATE U4266 ( .I1(n2143), .I2(\registres[11][12] ), .O(n3272) );
  NAND_GATE U4267 ( .I1(n2144), .I2(\registres[13][12] ), .O(n3271) );
  AND5_GATE U4268 ( .I1(n3280), .I2(n3281), .I3(n3282), .I4(n3283), .I5(n3284), 
        .O(n3259) );
  AND4_GATE U4269 ( .I1(n3285), .I2(n3286), .I3(n3287), .I4(n3288), .O(n3284)
         );
  NAND_GATE U4270 ( .I1(n2154), .I2(\registres[17][12] ), .O(n3288) );
  NAND_GATE U4271 ( .I1(n2155), .I2(\registres[19][12] ), .O(n3287) );
  NAND_GATE U4272 ( .I1(n2156), .I2(\registres[21][12] ), .O(n3286) );
  NAND_GATE U4273 ( .I1(n2157), .I2(\registres[6][12] ), .O(n3285) );
  NAND_GATE U4274 ( .I1(n2158), .I2(\registres[7][12] ), .O(n3283) );
  NAND_GATE U4275 ( .I1(n2159), .I2(\registres[30][12] ), .O(n3282) );
  NAND_GATE U4276 ( .I1(n2160), .I2(\registres[31][12] ), .O(n3281) );
  NAND_GATE U4277 ( .I1(n2161), .I2(\registres[14][12] ), .O(n3280) );
  AND4_GATE U4278 ( .I1(n3289), .I2(n3290), .I3(n3291), .I4(n3292), .O(n3258)
         );
  AND4_GATE U4279 ( .I1(n3293), .I2(n3294), .I3(n3295), .I4(n3296), .O(n3292)
         );
  NAND_GATE U4280 ( .I1(n2170), .I2(\registres[22][12] ), .O(n3296) );
  NAND_GATE U4281 ( .I1(n2171), .I2(\registres[15][12] ), .O(n3295) );
  NAND_GATE U4282 ( .I1(n2172), .I2(\registres[23][12] ), .O(n3294) );
  NAND_GATE U4283 ( .I1(n2173), .I2(\registres[4][12] ), .O(n3293) );
  NAND_GATE U4284 ( .I1(n2174), .I2(\registres[8][12] ), .O(n3291) );
  NAND_GATE U4285 ( .I1(n2175), .I2(\registres[2][12] ), .O(n3290) );
  NAND_GATE U4286 ( .I1(n2176), .I2(\registres[16][12] ), .O(n3289) );
  AND_GATE U4287 ( .I1(n3297), .I2(n2105), .O(data_src2[11]) );
  NAND4_GATE U4288 ( .I1(n3298), .I2(n3299), .I3(n3300), .I4(n3301), .O(n3297)
         );
  AND5_GATE U4289 ( .I1(n3302), .I2(n3303), .I3(n3304), .I4(n3305), .I5(n3306), 
        .O(n3301) );
  AND4_GATE U4290 ( .I1(n3307), .I2(n3308), .I3(n3309), .I4(n3310), .O(n3306)
         );
  NAND_GATE U4291 ( .I1(n2120), .I2(\registres[24][11] ), .O(n3310) );
  NAND_GATE U4292 ( .I1(n2121), .I2(\registres[25][11] ), .O(n3309) );
  NAND_GATE U4293 ( .I1(n2122), .I2(\registres[3][11] ), .O(n3308) );
  NAND_GATE U4294 ( .I1(n2123), .I2(\registres[26][11] ), .O(n3307) );
  NAND_GATE U4295 ( .I1(n2124), .I2(\registres[27][11] ), .O(n3305) );
  NAND_GATE U4296 ( .I1(n2125), .I2(\registres[10][11] ), .O(n3304) );
  NAND_GATE U4297 ( .I1(n2126), .I2(\registres[18][11] ), .O(n3303) );
  NAND_GATE U4298 ( .I1(n2127), .I2(\registres[5][11] ), .O(n3302) );
  AND5_GATE U4299 ( .I1(n3311), .I2(n3312), .I3(n3313), .I4(n3314), .I5(n3315), 
        .O(n3300) );
  AND4_GATE U4300 ( .I1(n3316), .I2(n3317), .I3(n3318), .I4(n3319), .O(n3315)
         );
  NAND_GATE U4301 ( .I1(n2137), .I2(\registres[28][11] ), .O(n3319) );
  NAND_GATE U4302 ( .I1(n2138), .I2(\registres[29][11] ), .O(n3318) );
  NAND_GATE U4303 ( .I1(n2139), .I2(\registres[12][11] ), .O(n3317) );
  NAND_GATE U4304 ( .I1(n2140), .I2(\registres[20][11] ), .O(n3316) );
  NAND_GATE U4305 ( .I1(n2141), .I2(\registres[1][11] ), .O(n3314) );
  NAND_GATE U4306 ( .I1(n2142), .I2(\registres[9][11] ), .O(n3313) );
  NAND_GATE U4307 ( .I1(n2143), .I2(\registres[11][11] ), .O(n3312) );
  NAND_GATE U4308 ( .I1(n2144), .I2(\registres[13][11] ), .O(n3311) );
  AND5_GATE U4309 ( .I1(n3320), .I2(n3321), .I3(n3322), .I4(n3323), .I5(n3324), 
        .O(n3299) );
  AND4_GATE U4310 ( .I1(n3325), .I2(n3326), .I3(n3327), .I4(n3328), .O(n3324)
         );
  NAND_GATE U4311 ( .I1(n2154), .I2(\registres[17][11] ), .O(n3328) );
  NAND_GATE U4312 ( .I1(n2155), .I2(\registres[19][11] ), .O(n3327) );
  NAND_GATE U4313 ( .I1(n2156), .I2(\registres[21][11] ), .O(n3326) );
  NAND_GATE U4314 ( .I1(n2157), .I2(\registres[6][11] ), .O(n3325) );
  NAND_GATE U4315 ( .I1(n2158), .I2(\registres[7][11] ), .O(n3323) );
  NAND_GATE U4316 ( .I1(n2159), .I2(\registres[30][11] ), .O(n3322) );
  NAND_GATE U4317 ( .I1(n2160), .I2(\registres[31][11] ), .O(n3321) );
  NAND_GATE U4318 ( .I1(n2161), .I2(\registres[14][11] ), .O(n3320) );
  AND4_GATE U4319 ( .I1(n3329), .I2(n3330), .I3(n3331), .I4(n3332), .O(n3298)
         );
  AND4_GATE U4320 ( .I1(n3333), .I2(n3334), .I3(n3335), .I4(n3336), .O(n3332)
         );
  NAND_GATE U4321 ( .I1(n2170), .I2(\registres[22][11] ), .O(n3336) );
  NAND_GATE U4322 ( .I1(n2171), .I2(\registres[15][11] ), .O(n3335) );
  NAND_GATE U4323 ( .I1(n2172), .I2(\registres[23][11] ), .O(n3334) );
  NAND_GATE U4324 ( .I1(n2173), .I2(\registres[4][11] ), .O(n3333) );
  NAND_GATE U4325 ( .I1(n2174), .I2(\registres[8][11] ), .O(n3331) );
  NAND_GATE U4326 ( .I1(n2175), .I2(\registres[2][11] ), .O(n3330) );
  NAND_GATE U4327 ( .I1(n2176), .I2(\registres[16][11] ), .O(n3329) );
  AND_GATE U4328 ( .I1(n3337), .I2(n2105), .O(data_src2[10]) );
  NAND4_GATE U4329 ( .I1(n3338), .I2(n3339), .I3(n3340), .I4(n3341), .O(n3337)
         );
  AND5_GATE U4330 ( .I1(n3342), .I2(n3343), .I3(n3344), .I4(n3345), .I5(n3346), 
        .O(n3341) );
  AND4_GATE U4331 ( .I1(n3347), .I2(n3348), .I3(n3349), .I4(n3350), .O(n3346)
         );
  NAND_GATE U4332 ( .I1(n2120), .I2(\registres[24][10] ), .O(n3350) );
  NAND_GATE U4333 ( .I1(n2121), .I2(\registres[25][10] ), .O(n3349) );
  NAND_GATE U4334 ( .I1(n2122), .I2(\registres[3][10] ), .O(n3348) );
  NAND_GATE U4335 ( .I1(n2123), .I2(\registres[26][10] ), .O(n3347) );
  NAND_GATE U4336 ( .I1(n2124), .I2(\registres[27][10] ), .O(n3345) );
  NAND_GATE U4337 ( .I1(n2125), .I2(\registres[10][10] ), .O(n3344) );
  NAND_GATE U4338 ( .I1(n2126), .I2(\registres[18][10] ), .O(n3343) );
  NAND_GATE U4339 ( .I1(n2127), .I2(\registres[5][10] ), .O(n3342) );
  AND5_GATE U4340 ( .I1(n3351), .I2(n3352), .I3(n3353), .I4(n3354), .I5(n3355), 
        .O(n3340) );
  AND4_GATE U4341 ( .I1(n3356), .I2(n3357), .I3(n3358), .I4(n3359), .O(n3355)
         );
  NAND_GATE U4342 ( .I1(n2137), .I2(\registres[28][10] ), .O(n3359) );
  NAND_GATE U4343 ( .I1(n2138), .I2(\registres[29][10] ), .O(n3358) );
  NAND_GATE U4344 ( .I1(n2139), .I2(\registres[12][10] ), .O(n3357) );
  NAND_GATE U4345 ( .I1(n2140), .I2(\registres[20][10] ), .O(n3356) );
  NAND_GATE U4346 ( .I1(n2141), .I2(\registres[1][10] ), .O(n3354) );
  NAND_GATE U4347 ( .I1(n2142), .I2(\registres[9][10] ), .O(n3353) );
  NAND_GATE U4348 ( .I1(n2143), .I2(\registres[11][10] ), .O(n3352) );
  NAND_GATE U4349 ( .I1(n2144), .I2(\registres[13][10] ), .O(n3351) );
  AND5_GATE U4350 ( .I1(n3360), .I2(n3361), .I3(n3362), .I4(n3363), .I5(n3364), 
        .O(n3339) );
  AND4_GATE U4351 ( .I1(n3365), .I2(n3366), .I3(n3367), .I4(n3368), .O(n3364)
         );
  NAND_GATE U4352 ( .I1(n2154), .I2(\registres[17][10] ), .O(n3368) );
  NAND_GATE U4353 ( .I1(n2155), .I2(\registres[19][10] ), .O(n3367) );
  NAND_GATE U4354 ( .I1(n2156), .I2(\registres[21][10] ), .O(n3366) );
  NAND_GATE U4355 ( .I1(n2157), .I2(\registres[6][10] ), .O(n3365) );
  NAND_GATE U4356 ( .I1(n2158), .I2(\registres[7][10] ), .O(n3363) );
  NAND_GATE U4357 ( .I1(n2159), .I2(\registres[30][10] ), .O(n3362) );
  NAND_GATE U4358 ( .I1(n2160), .I2(\registres[31][10] ), .O(n3361) );
  NAND_GATE U4359 ( .I1(n2161), .I2(\registres[14][10] ), .O(n3360) );
  AND4_GATE U4360 ( .I1(n3369), .I2(n3370), .I3(n3371), .I4(n3372), .O(n3338)
         );
  AND4_GATE U4361 ( .I1(n3373), .I2(n3374), .I3(n3375), .I4(n3376), .O(n3372)
         );
  NAND_GATE U4362 ( .I1(n2170), .I2(\registres[22][10] ), .O(n3376) );
  NAND_GATE U4363 ( .I1(n2171), .I2(\registres[15][10] ), .O(n3375) );
  NAND_GATE U4364 ( .I1(n2172), .I2(\registres[23][10] ), .O(n3374) );
  NAND_GATE U4365 ( .I1(n2173), .I2(\registres[4][10] ), .O(n3373) );
  NAND_GATE U4366 ( .I1(n2174), .I2(\registres[8][10] ), .O(n3371) );
  NAND_GATE U4367 ( .I1(n2175), .I2(\registres[2][10] ), .O(n3370) );
  NAND_GATE U4368 ( .I1(n2176), .I2(\registres[16][10] ), .O(n3369) );
  AND_GATE U4369 ( .I1(n3377), .I2(n2105), .O(data_src2[0]) );
  NAND_GATE U4370 ( .I1(n2174), .I2(n13), .O(n2105) );
  NAND4_GATE U4371 ( .I1(n3378), .I2(n3379), .I3(n3380), .I4(n3381), .O(n3377)
         );
  AND5_GATE U4372 ( .I1(n3382), .I2(n3383), .I3(n3384), .I4(n3385), .I5(n3386), 
        .O(n3381) );
  AND4_GATE U4373 ( .I1(n3387), .I2(n3388), .I3(n3389), .I4(n3390), .O(n3386)
         );
  NAND_GATE U4374 ( .I1(n2120), .I2(\registres[24][0] ), .O(n3390) );
  AND_GATE U4375 ( .I1(n3391), .I2(n3392), .O(n2120) );
  NAND_GATE U4376 ( .I1(n2121), .I2(\registres[25][0] ), .O(n3389) );
  AND_GATE U4377 ( .I1(n3393), .I2(n3391), .O(n2121) );
  NAND_GATE U4378 ( .I1(n2122), .I2(\registres[3][0] ), .O(n3388) );
  AND_GATE U4379 ( .I1(n3394), .I2(n3395), .O(n2122) );
  NAND_GATE U4380 ( .I1(n2123), .I2(\registres[26][0] ), .O(n3387) );
  AND_GATE U4381 ( .I1(n3394), .I2(n3392), .O(n2123) );
  NAND_GATE U4382 ( .I1(n2124), .I2(\registres[27][0] ), .O(n3385) );
  AND_GATE U4383 ( .I1(n3394), .I2(n3393), .O(n2124) );
  NAND_GATE U4384 ( .I1(n2125), .I2(\registres[10][0] ), .O(n3384) );
  AND_GATE U4385 ( .I1(n3396), .I2(n3394), .O(n2125) );
  NAND_GATE U4386 ( .I1(n2126), .I2(\registres[18][0] ), .O(n3383) );
  AND_GATE U4387 ( .I1(n3397), .I2(n3394), .O(n2126) );
  NAND_GATE U4388 ( .I1(n2127), .I2(\registres[5][0] ), .O(n3382) );
  AND_GATE U4389 ( .I1(n3398), .I2(n3395), .O(n2127) );
  AND5_GATE U4390 ( .I1(n3399), .I2(n3400), .I3(n3401), .I4(n3402), .I5(n3403), 
        .O(n3380) );
  AND4_GATE U4391 ( .I1(n3404), .I2(n3405), .I3(n3406), .I4(n3407), .O(n3403)
         );
  NAND_GATE U4392 ( .I1(n2137), .I2(\registres[28][0] ), .O(n3407) );
  AND_GATE U4393 ( .I1(n3398), .I2(n3392), .O(n2137) );
  NAND_GATE U4394 ( .I1(n2138), .I2(\registres[29][0] ), .O(n3406) );
  AND_GATE U4395 ( .I1(n3398), .I2(n3393), .O(n2138) );
  NAND_GATE U4396 ( .I1(n2139), .I2(\registres[12][0] ), .O(n3405) );
  AND_GATE U4397 ( .I1(n3398), .I2(n3396), .O(n2139) );
  NAND_GATE U4398 ( .I1(n2140), .I2(\registres[20][0] ), .O(n3404) );
  AND_GATE U4399 ( .I1(n3398), .I2(n3397), .O(n2140) );
  NAND_GATE U4400 ( .I1(n2141), .I2(\registres[1][0] ), .O(n3402) );
  AND_GATE U4401 ( .I1(n3408), .I2(n3391), .O(n2141) );
  NAND_GATE U4402 ( .I1(n2142), .I2(\registres[9][0] ), .O(n3401) );
  AND_GATE U4403 ( .I1(n3409), .I2(n3391), .O(n2142) );
  NAND_GATE U4404 ( .I1(n2143), .I2(\registres[11][0] ), .O(n3400) );
  AND_GATE U4405 ( .I1(n3409), .I2(n3394), .O(n2143) );
  NAND_GATE U4406 ( .I1(n2144), .I2(\registres[13][0] ), .O(n3399) );
  AND_GATE U4407 ( .I1(n3409), .I2(n3398), .O(n2144) );
  AND5_GATE U4408 ( .I1(n3410), .I2(n3411), .I3(n3412), .I4(n3413), .I5(n3414), 
        .O(n3379) );
  AND4_GATE U4409 ( .I1(n3415), .I2(n3416), .I3(n3417), .I4(n3418), .O(n3414)
         );
  NAND_GATE U4410 ( .I1(n2154), .I2(\registres[17][0] ), .O(n3418) );
  AND_GATE U4411 ( .I1(n3419), .I2(n3391), .O(n2154) );
  NAND_GATE U4412 ( .I1(n2155), .I2(\registres[19][0] ), .O(n3417) );
  AND_GATE U4413 ( .I1(n3419), .I2(n3394), .O(n2155) );
  NOR_GATE U4414 ( .I1(n11), .I2(reg_src2[2]), .O(n3394) );
  NAND_GATE U4415 ( .I1(n2156), .I2(\registres[21][0] ), .O(n3416) );
  AND_GATE U4416 ( .I1(n3419), .I2(n3398), .O(n2156) );
  NOR_GATE U4417 ( .I1(n12), .I2(reg_src2[1]), .O(n3398) );
  NAND_GATE U4418 ( .I1(n2157), .I2(\registres[6][0] ), .O(n3415) );
  AND_GATE U4419 ( .I1(n3420), .I2(n3421), .O(n2157) );
  NAND_GATE U4420 ( .I1(n2158), .I2(\registres[7][0] ), .O(n3413) );
  AND_GATE U4421 ( .I1(n3420), .I2(n3395), .O(n2158) );
  AND_GATE U4422 ( .I1(n3408), .I2(reg_src2[0]), .O(n3395) );
  NAND_GATE U4423 ( .I1(n2159), .I2(\registres[30][0] ), .O(n3412) );
  AND_GATE U4424 ( .I1(n3420), .I2(n3392), .O(n2159) );
  AND_GATE U4425 ( .I1(n3422), .I2(n10), .O(n3392) );
  NAND_GATE U4426 ( .I1(n2160), .I2(\registres[31][0] ), .O(n3411) );
  AND_GATE U4427 ( .I1(n3420), .I2(n3393), .O(n2160) );
  AND_GATE U4428 ( .I1(reg_src2[0]), .I2(n3422), .O(n3393) );
  NOR_GATE U4429 ( .I1(n14), .I2(n13), .O(n3422) );
  NAND_GATE U4430 ( .I1(n2161), .I2(\registres[14][0] ), .O(n3410) );
  AND_GATE U4431 ( .I1(n3420), .I2(n3396), .O(n2161) );
  NOR3_GATE U4432 ( .I1(reg_src2[0]), .I2(reg_src2[4]), .I3(n13), .O(n3396) );
  AND4_GATE U4433 ( .I1(n3423), .I2(n3424), .I3(n3425), .I4(n3426), .O(n3378)
         );
  AND4_GATE U4434 ( .I1(n3427), .I2(n3428), .I3(n3429), .I4(n3430), .O(n3426)
         );
  NAND_GATE U4435 ( .I1(n2170), .I2(\registres[22][0] ), .O(n3430) );
  AND_GATE U4436 ( .I1(n3420), .I2(n3397), .O(n2170) );
  NOR3_GATE U4437 ( .I1(reg_src2[0]), .I2(reg_src2[3]), .I3(n14), .O(n3397) );
  NAND_GATE U4438 ( .I1(n2171), .I2(\registres[15][0] ), .O(n3429) );
  AND_GATE U4439 ( .I1(n3420), .I2(n3409), .O(n2171) );
  NOR3_GATE U4440 ( .I1(n13), .I2(reg_src2[4]), .I3(n10), .O(n3409) );
  NAND_GATE U4441 ( .I1(n2172), .I2(\registres[23][0] ), .O(n3428) );
  AND_GATE U4442 ( .I1(n3420), .I2(n3419), .O(n2172) );
  NOR3_GATE U4443 ( .I1(n14), .I2(reg_src2[3]), .I3(n10), .O(n3419) );
  NOR_GATE U4444 ( .I1(n12), .I2(n11), .O(n3420) );
  NAND_GATE U4445 ( .I1(n2173), .I2(\registres[4][0] ), .O(n3427) );
  AND_GATE U4446 ( .I1(n3421), .I2(n11), .O(n2173) );
  NAND_GATE U4447 ( .I1(n2174), .I2(\registres[8][0] ), .O(n3425) );
  AND_GATE U4448 ( .I1(n3431), .I2(n14), .O(n2174) );
  NAND_GATE U4449 ( .I1(n2175), .I2(\registres[2][0] ), .O(n3424) );
  AND_GATE U4450 ( .I1(n3421), .I2(n12), .O(n2175) );
  AND_GATE U4451 ( .I1(n3408), .I2(n10), .O(n3421) );
  NOR_GATE U4452 ( .I1(reg_src2[4]), .I2(reg_src2[3]), .O(n3408) );
  NAND_GATE U4453 ( .I1(n2176), .I2(\registres[16][0] ), .O(n3423) );
  AND_GATE U4454 ( .I1(n3431), .I2(n13), .O(n2176) );
  AND_GATE U4455 ( .I1(n3391), .I2(n10), .O(n3431) );
  NOR_GATE U4456 ( .I1(reg_src2[2]), .I2(reg_src2[1]), .O(n3391) );
  AND_GATE U4457 ( .I1(n3432), .I2(n3433), .O(data_src1[9]) );
  NAND4_GATE U4458 ( .I1(n3434), .I2(n3435), .I3(n3436), .I4(n3437), .O(n3433)
         );
  AND5_GATE U4459 ( .I1(n3438), .I2(n3439), .I3(n3440), .I4(n3441), .I5(n3442), 
        .O(n3437) );
  AND4_GATE U4460 ( .I1(n3443), .I2(n3444), .I3(n3445), .I4(n3446), .O(n3442)
         );
  NAND_GATE U4461 ( .I1(n3447), .I2(\registres[24][9] ), .O(n3446) );
  NAND_GATE U4462 ( .I1(n3448), .I2(\registres[25][9] ), .O(n3445) );
  NAND_GATE U4463 ( .I1(n3449), .I2(\registres[3][9] ), .O(n3444) );
  NAND_GATE U4464 ( .I1(n3450), .I2(\registres[26][9] ), .O(n3443) );
  NAND_GATE U4465 ( .I1(n3451), .I2(\registres[27][9] ), .O(n3441) );
  NAND_GATE U4466 ( .I1(n3452), .I2(\registres[10][9] ), .O(n3440) );
  NAND_GATE U4467 ( .I1(n3453), .I2(\registres[18][9] ), .O(n3439) );
  NAND_GATE U4468 ( .I1(n3454), .I2(\registres[5][9] ), .O(n3438) );
  AND5_GATE U4469 ( .I1(n3455), .I2(n3456), .I3(n3457), .I4(n3458), .I5(n3459), 
        .O(n3436) );
  AND4_GATE U4470 ( .I1(n3460), .I2(n3461), .I3(n3462), .I4(n3463), .O(n3459)
         );
  NAND_GATE U4471 ( .I1(n3464), .I2(\registres[28][9] ), .O(n3463) );
  NAND_GATE U4472 ( .I1(n3465), .I2(\registres[29][9] ), .O(n3462) );
  NAND_GATE U4473 ( .I1(n3466), .I2(\registres[12][9] ), .O(n3461) );
  NAND_GATE U4474 ( .I1(n3467), .I2(\registres[20][9] ), .O(n3460) );
  NAND_GATE U4475 ( .I1(n3468), .I2(\registres[1][9] ), .O(n3458) );
  NAND_GATE U4476 ( .I1(n3469), .I2(\registres[9][9] ), .O(n3457) );
  NAND_GATE U4477 ( .I1(n3470), .I2(\registres[11][9] ), .O(n3456) );
  NAND_GATE U4478 ( .I1(n3471), .I2(\registres[13][9] ), .O(n3455) );
  AND5_GATE U4479 ( .I1(n3472), .I2(n3473), .I3(n3474), .I4(n3475), .I5(n3476), 
        .O(n3435) );
  AND4_GATE U4480 ( .I1(n3477), .I2(n3478), .I3(n3479), .I4(n3480), .O(n3476)
         );
  NAND_GATE U4481 ( .I1(n3481), .I2(\registres[17][9] ), .O(n3480) );
  NAND_GATE U4482 ( .I1(n3482), .I2(\registres[19][9] ), .O(n3479) );
  NAND_GATE U4483 ( .I1(n3483), .I2(\registres[21][9] ), .O(n3478) );
  NAND_GATE U4484 ( .I1(n3484), .I2(\registres[6][9] ), .O(n3477) );
  NAND_GATE U4485 ( .I1(n3485), .I2(\registres[7][9] ), .O(n3475) );
  NAND_GATE U4486 ( .I1(n3486), .I2(\registres[30][9] ), .O(n3474) );
  NAND_GATE U4487 ( .I1(n3487), .I2(\registres[31][9] ), .O(n3473) );
  NAND_GATE U4488 ( .I1(n3488), .I2(\registres[14][9] ), .O(n3472) );
  AND4_GATE U4489 ( .I1(n3489), .I2(n3490), .I3(n3491), .I4(n3492), .O(n3434)
         );
  AND4_GATE U4490 ( .I1(n3493), .I2(n3494), .I3(n3495), .I4(n3496), .O(n3492)
         );
  NAND_GATE U4491 ( .I1(n3497), .I2(\registres[22][9] ), .O(n3496) );
  NAND_GATE U4492 ( .I1(n3498), .I2(\registres[15][9] ), .O(n3495) );
  NAND_GATE U4493 ( .I1(n3499), .I2(\registres[23][9] ), .O(n3494) );
  NAND_GATE U4494 ( .I1(n3500), .I2(\registres[4][9] ), .O(n3493) );
  NAND_GATE U4495 ( .I1(n3501), .I2(\registres[8][9] ), .O(n3491) );
  NAND_GATE U4496 ( .I1(n3502), .I2(\registres[2][9] ), .O(n3490) );
  NAND_GATE U4497 ( .I1(n3503), .I2(\registres[16][9] ), .O(n3489) );
  AND_GATE U4498 ( .I1(n3504), .I2(n3432), .O(data_src1[8]) );
  NAND4_GATE U4499 ( .I1(n3505), .I2(n3506), .I3(n3507), .I4(n3508), .O(n3504)
         );
  AND5_GATE U4500 ( .I1(n3509), .I2(n3510), .I3(n3511), .I4(n3512), .I5(n3513), 
        .O(n3508) );
  AND4_GATE U4501 ( .I1(n3514), .I2(n3515), .I3(n3516), .I4(n3517), .O(n3513)
         );
  NAND_GATE U4502 ( .I1(n3447), .I2(\registres[24][8] ), .O(n3517) );
  NAND_GATE U4503 ( .I1(n3448), .I2(\registres[25][8] ), .O(n3516) );
  NAND_GATE U4504 ( .I1(n3449), .I2(\registres[3][8] ), .O(n3515) );
  NAND_GATE U4505 ( .I1(n3450), .I2(\registres[26][8] ), .O(n3514) );
  NAND_GATE U4506 ( .I1(n3451), .I2(\registres[27][8] ), .O(n3512) );
  NAND_GATE U4507 ( .I1(n3452), .I2(\registres[10][8] ), .O(n3511) );
  NAND_GATE U4508 ( .I1(n3453), .I2(\registres[18][8] ), .O(n3510) );
  NAND_GATE U4509 ( .I1(n3454), .I2(\registres[5][8] ), .O(n3509) );
  AND5_GATE U4510 ( .I1(n3518), .I2(n3519), .I3(n3520), .I4(n3521), .I5(n3522), 
        .O(n3507) );
  AND4_GATE U4511 ( .I1(n3523), .I2(n3524), .I3(n3525), .I4(n3526), .O(n3522)
         );
  NAND_GATE U4512 ( .I1(n3464), .I2(\registres[28][8] ), .O(n3526) );
  NAND_GATE U4513 ( .I1(n3465), .I2(\registres[29][8] ), .O(n3525) );
  NAND_GATE U4514 ( .I1(n3466), .I2(\registres[12][8] ), .O(n3524) );
  NAND_GATE U4515 ( .I1(n3467), .I2(\registres[20][8] ), .O(n3523) );
  NAND_GATE U4516 ( .I1(n3468), .I2(\registres[1][8] ), .O(n3521) );
  NAND_GATE U4517 ( .I1(n3469), .I2(\registres[9][8] ), .O(n3520) );
  NAND_GATE U4518 ( .I1(n3470), .I2(\registres[11][8] ), .O(n3519) );
  NAND_GATE U4519 ( .I1(n3471), .I2(\registres[13][8] ), .O(n3518) );
  AND5_GATE U4520 ( .I1(n3527), .I2(n3528), .I3(n3529), .I4(n3530), .I5(n3531), 
        .O(n3506) );
  AND4_GATE U4521 ( .I1(n3532), .I2(n3533), .I3(n3534), .I4(n3535), .O(n3531)
         );
  NAND_GATE U4522 ( .I1(n3481), .I2(\registres[17][8] ), .O(n3535) );
  NAND_GATE U4523 ( .I1(n3482), .I2(\registres[19][8] ), .O(n3534) );
  NAND_GATE U4524 ( .I1(n3483), .I2(\registres[21][8] ), .O(n3533) );
  NAND_GATE U4525 ( .I1(n3484), .I2(\registres[6][8] ), .O(n3532) );
  NAND_GATE U4526 ( .I1(n3485), .I2(\registres[7][8] ), .O(n3530) );
  NAND_GATE U4527 ( .I1(n3486), .I2(\registres[30][8] ), .O(n3529) );
  NAND_GATE U4528 ( .I1(n3487), .I2(\registres[31][8] ), .O(n3528) );
  NAND_GATE U4529 ( .I1(n3488), .I2(\registres[14][8] ), .O(n3527) );
  AND4_GATE U4530 ( .I1(n3536), .I2(n3537), .I3(n3538), .I4(n3539), .O(n3505)
         );
  AND4_GATE U4531 ( .I1(n3540), .I2(n3541), .I3(n3542), .I4(n3543), .O(n3539)
         );
  NAND_GATE U4532 ( .I1(n3497), .I2(\registres[22][8] ), .O(n3543) );
  NAND_GATE U4533 ( .I1(n3498), .I2(\registres[15][8] ), .O(n3542) );
  NAND_GATE U4534 ( .I1(n3499), .I2(\registres[23][8] ), .O(n3541) );
  NAND_GATE U4535 ( .I1(n3500), .I2(\registres[4][8] ), .O(n3540) );
  NAND_GATE U4536 ( .I1(n3501), .I2(\registres[8][8] ), .O(n3538) );
  NAND_GATE U4537 ( .I1(n3502), .I2(\registres[2][8] ), .O(n3537) );
  NAND_GATE U4538 ( .I1(n3503), .I2(\registres[16][8] ), .O(n3536) );
  AND_GATE U4539 ( .I1(n3544), .I2(n3432), .O(data_src1[7]) );
  NAND4_GATE U4540 ( .I1(n3545), .I2(n3546), .I3(n3547), .I4(n3548), .O(n3544)
         );
  AND5_GATE U4541 ( .I1(n3549), .I2(n3550), .I3(n3551), .I4(n3552), .I5(n3553), 
        .O(n3548) );
  AND4_GATE U4542 ( .I1(n3554), .I2(n3555), .I3(n3556), .I4(n3557), .O(n3553)
         );
  NAND_GATE U4543 ( .I1(n3447), .I2(\registres[24][7] ), .O(n3557) );
  NAND_GATE U4544 ( .I1(n3448), .I2(\registres[25][7] ), .O(n3556) );
  NAND_GATE U4545 ( .I1(n3449), .I2(\registres[3][7] ), .O(n3555) );
  NAND_GATE U4546 ( .I1(n3450), .I2(\registres[26][7] ), .O(n3554) );
  NAND_GATE U4547 ( .I1(n3451), .I2(\registres[27][7] ), .O(n3552) );
  NAND_GATE U4548 ( .I1(n3452), .I2(\registres[10][7] ), .O(n3551) );
  NAND_GATE U4549 ( .I1(n3453), .I2(\registres[18][7] ), .O(n3550) );
  NAND_GATE U4550 ( .I1(n3454), .I2(\registres[5][7] ), .O(n3549) );
  AND5_GATE U4551 ( .I1(n3558), .I2(n3559), .I3(n3560), .I4(n3561), .I5(n3562), 
        .O(n3547) );
  AND4_GATE U4552 ( .I1(n3563), .I2(n3564), .I3(n3565), .I4(n3566), .O(n3562)
         );
  NAND_GATE U4553 ( .I1(n3464), .I2(\registres[28][7] ), .O(n3566) );
  NAND_GATE U4554 ( .I1(n3465), .I2(\registres[29][7] ), .O(n3565) );
  NAND_GATE U4555 ( .I1(n3466), .I2(\registres[12][7] ), .O(n3564) );
  NAND_GATE U4556 ( .I1(n3467), .I2(\registres[20][7] ), .O(n3563) );
  NAND_GATE U4557 ( .I1(n3468), .I2(\registres[1][7] ), .O(n3561) );
  NAND_GATE U4558 ( .I1(n3469), .I2(\registres[9][7] ), .O(n3560) );
  NAND_GATE U4559 ( .I1(n3470), .I2(\registres[11][7] ), .O(n3559) );
  NAND_GATE U4560 ( .I1(n3471), .I2(\registres[13][7] ), .O(n3558) );
  AND5_GATE U4561 ( .I1(n3567), .I2(n3568), .I3(n3569), .I4(n3570), .I5(n3571), 
        .O(n3546) );
  AND4_GATE U4562 ( .I1(n3572), .I2(n3573), .I3(n3574), .I4(n3575), .O(n3571)
         );
  NAND_GATE U4563 ( .I1(n3481), .I2(\registres[17][7] ), .O(n3575) );
  NAND_GATE U4564 ( .I1(n3482), .I2(\registres[19][7] ), .O(n3574) );
  NAND_GATE U4565 ( .I1(n3483), .I2(\registres[21][7] ), .O(n3573) );
  NAND_GATE U4566 ( .I1(n3484), .I2(\registres[6][7] ), .O(n3572) );
  NAND_GATE U4567 ( .I1(n3485), .I2(\registres[7][7] ), .O(n3570) );
  NAND_GATE U4568 ( .I1(n3486), .I2(\registres[30][7] ), .O(n3569) );
  NAND_GATE U4569 ( .I1(n3487), .I2(\registres[31][7] ), .O(n3568) );
  NAND_GATE U4570 ( .I1(n3488), .I2(\registres[14][7] ), .O(n3567) );
  AND4_GATE U4571 ( .I1(n3576), .I2(n3577), .I3(n3578), .I4(n3579), .O(n3545)
         );
  AND4_GATE U4572 ( .I1(n3580), .I2(n3581), .I3(n3582), .I4(n3583), .O(n3579)
         );
  NAND_GATE U4573 ( .I1(n3497), .I2(\registres[22][7] ), .O(n3583) );
  NAND_GATE U4574 ( .I1(n3498), .I2(\registres[15][7] ), .O(n3582) );
  NAND_GATE U4575 ( .I1(n3499), .I2(\registres[23][7] ), .O(n3581) );
  NAND_GATE U4576 ( .I1(n3500), .I2(\registres[4][7] ), .O(n3580) );
  NAND_GATE U4577 ( .I1(n3501), .I2(\registres[8][7] ), .O(n3578) );
  NAND_GATE U4578 ( .I1(n3502), .I2(\registres[2][7] ), .O(n3577) );
  NAND_GATE U4579 ( .I1(n3503), .I2(\registres[16][7] ), .O(n3576) );
  AND_GATE U4580 ( .I1(n3584), .I2(n3432), .O(data_src1[6]) );
  NAND4_GATE U4581 ( .I1(n3585), .I2(n3586), .I3(n3587), .I4(n3588), .O(n3584)
         );
  AND5_GATE U4582 ( .I1(n3589), .I2(n3590), .I3(n3591), .I4(n3592), .I5(n3593), 
        .O(n3588) );
  AND4_GATE U4583 ( .I1(n3594), .I2(n3595), .I3(n3596), .I4(n3597), .O(n3593)
         );
  NAND_GATE U4584 ( .I1(n3447), .I2(\registres[24][6] ), .O(n3597) );
  NAND_GATE U4585 ( .I1(n3448), .I2(\registres[25][6] ), .O(n3596) );
  NAND_GATE U4586 ( .I1(n3449), .I2(\registres[3][6] ), .O(n3595) );
  NAND_GATE U4587 ( .I1(n3450), .I2(\registres[26][6] ), .O(n3594) );
  NAND_GATE U4588 ( .I1(n3451), .I2(\registres[27][6] ), .O(n3592) );
  NAND_GATE U4589 ( .I1(n3452), .I2(\registres[10][6] ), .O(n3591) );
  NAND_GATE U4590 ( .I1(n3453), .I2(\registres[18][6] ), .O(n3590) );
  NAND_GATE U4591 ( .I1(n3454), .I2(\registres[5][6] ), .O(n3589) );
  AND5_GATE U4592 ( .I1(n3598), .I2(n3599), .I3(n3600), .I4(n3601), .I5(n3602), 
        .O(n3587) );
  AND4_GATE U4593 ( .I1(n3603), .I2(n3604), .I3(n3605), .I4(n3606), .O(n3602)
         );
  NAND_GATE U4594 ( .I1(n3464), .I2(\registres[28][6] ), .O(n3606) );
  NAND_GATE U4595 ( .I1(n3465), .I2(\registres[29][6] ), .O(n3605) );
  NAND_GATE U4596 ( .I1(n3466), .I2(\registres[12][6] ), .O(n3604) );
  NAND_GATE U4597 ( .I1(n3467), .I2(\registres[20][6] ), .O(n3603) );
  NAND_GATE U4598 ( .I1(n3468), .I2(\registres[1][6] ), .O(n3601) );
  NAND_GATE U4599 ( .I1(n3469), .I2(\registres[9][6] ), .O(n3600) );
  NAND_GATE U4600 ( .I1(n3470), .I2(\registres[11][6] ), .O(n3599) );
  NAND_GATE U4601 ( .I1(n3471), .I2(\registres[13][6] ), .O(n3598) );
  AND5_GATE U4602 ( .I1(n3607), .I2(n3608), .I3(n3609), .I4(n3610), .I5(n3611), 
        .O(n3586) );
  AND4_GATE U4603 ( .I1(n3612), .I2(n3613), .I3(n3614), .I4(n3615), .O(n3611)
         );
  NAND_GATE U4604 ( .I1(n3481), .I2(\registres[17][6] ), .O(n3615) );
  NAND_GATE U4605 ( .I1(n3482), .I2(\registres[19][6] ), .O(n3614) );
  NAND_GATE U4606 ( .I1(n3483), .I2(\registres[21][6] ), .O(n3613) );
  NAND_GATE U4607 ( .I1(n3484), .I2(\registres[6][6] ), .O(n3612) );
  NAND_GATE U4608 ( .I1(n3485), .I2(\registres[7][6] ), .O(n3610) );
  NAND_GATE U4609 ( .I1(n3486), .I2(\registres[30][6] ), .O(n3609) );
  NAND_GATE U4610 ( .I1(n3487), .I2(\registres[31][6] ), .O(n3608) );
  NAND_GATE U4611 ( .I1(n3488), .I2(\registres[14][6] ), .O(n3607) );
  AND4_GATE U4612 ( .I1(n3616), .I2(n3617), .I3(n3618), .I4(n3619), .O(n3585)
         );
  AND4_GATE U4613 ( .I1(n3620), .I2(n3621), .I3(n3622), .I4(n3623), .O(n3619)
         );
  NAND_GATE U4614 ( .I1(n3497), .I2(\registres[22][6] ), .O(n3623) );
  NAND_GATE U4615 ( .I1(n3498), .I2(\registres[15][6] ), .O(n3622) );
  NAND_GATE U4616 ( .I1(n3499), .I2(\registres[23][6] ), .O(n3621) );
  NAND_GATE U4617 ( .I1(n3500), .I2(\registres[4][6] ), .O(n3620) );
  NAND_GATE U4618 ( .I1(n3501), .I2(\registres[8][6] ), .O(n3618) );
  NAND_GATE U4619 ( .I1(n3502), .I2(\registres[2][6] ), .O(n3617) );
  NAND_GATE U4620 ( .I1(n3503), .I2(\registres[16][6] ), .O(n3616) );
  AND_GATE U4621 ( .I1(n3624), .I2(n3432), .O(data_src1[5]) );
  NAND4_GATE U4622 ( .I1(n3625), .I2(n3626), .I3(n3627), .I4(n3628), .O(n3624)
         );
  AND5_GATE U4623 ( .I1(n3629), .I2(n3630), .I3(n3631), .I4(n3632), .I5(n3633), 
        .O(n3628) );
  AND4_GATE U4624 ( .I1(n3634), .I2(n3635), .I3(n3636), .I4(n3637), .O(n3633)
         );
  NAND_GATE U4625 ( .I1(n3447), .I2(\registres[24][5] ), .O(n3637) );
  NAND_GATE U4626 ( .I1(n3448), .I2(\registres[25][5] ), .O(n3636) );
  NAND_GATE U4627 ( .I1(n3449), .I2(\registres[3][5] ), .O(n3635) );
  NAND_GATE U4628 ( .I1(n3450), .I2(\registres[26][5] ), .O(n3634) );
  NAND_GATE U4629 ( .I1(n3451), .I2(\registres[27][5] ), .O(n3632) );
  NAND_GATE U4630 ( .I1(n3452), .I2(\registres[10][5] ), .O(n3631) );
  NAND_GATE U4631 ( .I1(n3453), .I2(\registres[18][5] ), .O(n3630) );
  NAND_GATE U4632 ( .I1(n3454), .I2(\registres[5][5] ), .O(n3629) );
  AND5_GATE U4633 ( .I1(n3638), .I2(n3639), .I3(n3640), .I4(n3641), .I5(n3642), 
        .O(n3627) );
  AND4_GATE U4634 ( .I1(n3643), .I2(n3644), .I3(n3645), .I4(n3646), .O(n3642)
         );
  NAND_GATE U4635 ( .I1(n3464), .I2(\registres[28][5] ), .O(n3646) );
  NAND_GATE U4636 ( .I1(n3465), .I2(\registres[29][5] ), .O(n3645) );
  NAND_GATE U4637 ( .I1(n3466), .I2(\registres[12][5] ), .O(n3644) );
  NAND_GATE U4638 ( .I1(n3467), .I2(\registres[20][5] ), .O(n3643) );
  NAND_GATE U4639 ( .I1(n3468), .I2(\registres[1][5] ), .O(n3641) );
  NAND_GATE U4640 ( .I1(n3469), .I2(\registres[9][5] ), .O(n3640) );
  NAND_GATE U4641 ( .I1(n3470), .I2(\registres[11][5] ), .O(n3639) );
  NAND_GATE U4642 ( .I1(n3471), .I2(\registres[13][5] ), .O(n3638) );
  AND5_GATE U4643 ( .I1(n3647), .I2(n3648), .I3(n3649), .I4(n3650), .I5(n3651), 
        .O(n3626) );
  AND4_GATE U4644 ( .I1(n3652), .I2(n3653), .I3(n3654), .I4(n3655), .O(n3651)
         );
  NAND_GATE U4645 ( .I1(n3481), .I2(\registres[17][5] ), .O(n3655) );
  NAND_GATE U4646 ( .I1(n3482), .I2(\registres[19][5] ), .O(n3654) );
  NAND_GATE U4647 ( .I1(n3483), .I2(\registres[21][5] ), .O(n3653) );
  NAND_GATE U4648 ( .I1(n3484), .I2(\registres[6][5] ), .O(n3652) );
  NAND_GATE U4649 ( .I1(n3485), .I2(\registres[7][5] ), .O(n3650) );
  NAND_GATE U4650 ( .I1(n3486), .I2(\registres[30][5] ), .O(n3649) );
  NAND_GATE U4651 ( .I1(n3487), .I2(\registres[31][5] ), .O(n3648) );
  NAND_GATE U4652 ( .I1(n3488), .I2(\registres[14][5] ), .O(n3647) );
  AND4_GATE U4653 ( .I1(n3656), .I2(n3657), .I3(n3658), .I4(n3659), .O(n3625)
         );
  AND4_GATE U4654 ( .I1(n3660), .I2(n3661), .I3(n3662), .I4(n3663), .O(n3659)
         );
  NAND_GATE U4655 ( .I1(n3497), .I2(\registres[22][5] ), .O(n3663) );
  NAND_GATE U4656 ( .I1(n3498), .I2(\registres[15][5] ), .O(n3662) );
  NAND_GATE U4657 ( .I1(n3499), .I2(\registres[23][5] ), .O(n3661) );
  NAND_GATE U4658 ( .I1(n3500), .I2(\registres[4][5] ), .O(n3660) );
  NAND_GATE U4659 ( .I1(n3501), .I2(\registres[8][5] ), .O(n3658) );
  NAND_GATE U4660 ( .I1(n3502), .I2(\registres[2][5] ), .O(n3657) );
  NAND_GATE U4661 ( .I1(n3503), .I2(\registres[16][5] ), .O(n3656) );
  AND_GATE U4662 ( .I1(n3664), .I2(n3432), .O(data_src1[4]) );
  NAND4_GATE U4663 ( .I1(n3665), .I2(n3666), .I3(n3667), .I4(n3668), .O(n3664)
         );
  AND5_GATE U4664 ( .I1(n3669), .I2(n3670), .I3(n3671), .I4(n3672), .I5(n3673), 
        .O(n3668) );
  AND4_GATE U4665 ( .I1(n3674), .I2(n3675), .I3(n3676), .I4(n3677), .O(n3673)
         );
  NAND_GATE U4666 ( .I1(n3447), .I2(\registres[24][4] ), .O(n3677) );
  NAND_GATE U4667 ( .I1(n3448), .I2(\registres[25][4] ), .O(n3676) );
  NAND_GATE U4668 ( .I1(n3449), .I2(\registres[3][4] ), .O(n3675) );
  NAND_GATE U4669 ( .I1(n3450), .I2(\registres[26][4] ), .O(n3674) );
  NAND_GATE U4670 ( .I1(n3451), .I2(\registres[27][4] ), .O(n3672) );
  NAND_GATE U4671 ( .I1(n3452), .I2(\registres[10][4] ), .O(n3671) );
  NAND_GATE U4672 ( .I1(n3453), .I2(\registres[18][4] ), .O(n3670) );
  NAND_GATE U4673 ( .I1(n3454), .I2(\registres[5][4] ), .O(n3669) );
  AND5_GATE U4674 ( .I1(n3678), .I2(n3679), .I3(n3680), .I4(n3681), .I5(n3682), 
        .O(n3667) );
  AND4_GATE U4675 ( .I1(n3683), .I2(n3684), .I3(n3685), .I4(n3686), .O(n3682)
         );
  NAND_GATE U4676 ( .I1(n3464), .I2(\registres[28][4] ), .O(n3686) );
  NAND_GATE U4677 ( .I1(n3465), .I2(\registres[29][4] ), .O(n3685) );
  NAND_GATE U4678 ( .I1(n3466), .I2(\registres[12][4] ), .O(n3684) );
  NAND_GATE U4679 ( .I1(n3467), .I2(\registres[20][4] ), .O(n3683) );
  NAND_GATE U4680 ( .I1(n3468), .I2(\registres[1][4] ), .O(n3681) );
  NAND_GATE U4681 ( .I1(n3469), .I2(\registres[9][4] ), .O(n3680) );
  NAND_GATE U4682 ( .I1(n3470), .I2(\registres[11][4] ), .O(n3679) );
  NAND_GATE U4683 ( .I1(n3471), .I2(\registres[13][4] ), .O(n3678) );
  AND5_GATE U4684 ( .I1(n3687), .I2(n3688), .I3(n3689), .I4(n3690), .I5(n3691), 
        .O(n3666) );
  AND4_GATE U4685 ( .I1(n3692), .I2(n3693), .I3(n3694), .I4(n3695), .O(n3691)
         );
  NAND_GATE U4686 ( .I1(n3481), .I2(\registres[17][4] ), .O(n3695) );
  NAND_GATE U4687 ( .I1(n3482), .I2(\registres[19][4] ), .O(n3694) );
  NAND_GATE U4688 ( .I1(n3483), .I2(\registres[21][4] ), .O(n3693) );
  NAND_GATE U4689 ( .I1(n3484), .I2(\registres[6][4] ), .O(n3692) );
  NAND_GATE U4690 ( .I1(n3485), .I2(\registres[7][4] ), .O(n3690) );
  NAND_GATE U4691 ( .I1(n3486), .I2(\registres[30][4] ), .O(n3689) );
  NAND_GATE U4692 ( .I1(n3487), .I2(\registres[31][4] ), .O(n3688) );
  NAND_GATE U4693 ( .I1(n3488), .I2(\registres[14][4] ), .O(n3687) );
  AND4_GATE U4694 ( .I1(n3696), .I2(n3697), .I3(n3698), .I4(n3699), .O(n3665)
         );
  AND4_GATE U4695 ( .I1(n3700), .I2(n3701), .I3(n3702), .I4(n3703), .O(n3699)
         );
  NAND_GATE U4696 ( .I1(n3497), .I2(\registres[22][4] ), .O(n3703) );
  NAND_GATE U4697 ( .I1(n3498), .I2(\registres[15][4] ), .O(n3702) );
  NAND_GATE U4698 ( .I1(n3499), .I2(\registres[23][4] ), .O(n3701) );
  NAND_GATE U4699 ( .I1(n3500), .I2(\registres[4][4] ), .O(n3700) );
  NAND_GATE U4700 ( .I1(n3501), .I2(\registres[8][4] ), .O(n3698) );
  NAND_GATE U4701 ( .I1(n3502), .I2(\registres[2][4] ), .O(n3697) );
  NAND_GATE U4702 ( .I1(n3503), .I2(\registres[16][4] ), .O(n3696) );
  AND_GATE U4703 ( .I1(n3704), .I2(n3432), .O(data_src1[3]) );
  NAND4_GATE U4704 ( .I1(n3705), .I2(n3706), .I3(n3707), .I4(n3708), .O(n3704)
         );
  AND5_GATE U4705 ( .I1(n3709), .I2(n3710), .I3(n3711), .I4(n3712), .I5(n3713), 
        .O(n3708) );
  AND4_GATE U4706 ( .I1(n3714), .I2(n3715), .I3(n3716), .I4(n3717), .O(n3713)
         );
  NAND_GATE U4707 ( .I1(n3447), .I2(\registres[24][3] ), .O(n3717) );
  NAND_GATE U4708 ( .I1(n3448), .I2(\registres[25][3] ), .O(n3716) );
  NAND_GATE U4709 ( .I1(n3449), .I2(\registres[3][3] ), .O(n3715) );
  NAND_GATE U4710 ( .I1(n3450), .I2(\registres[26][3] ), .O(n3714) );
  NAND_GATE U4711 ( .I1(n3451), .I2(\registres[27][3] ), .O(n3712) );
  NAND_GATE U4712 ( .I1(n3452), .I2(\registres[10][3] ), .O(n3711) );
  NAND_GATE U4713 ( .I1(n3453), .I2(\registres[18][3] ), .O(n3710) );
  NAND_GATE U4714 ( .I1(n3454), .I2(\registres[5][3] ), .O(n3709) );
  AND5_GATE U4715 ( .I1(n3718), .I2(n3719), .I3(n3720), .I4(n3721), .I5(n3722), 
        .O(n3707) );
  AND4_GATE U4716 ( .I1(n3723), .I2(n3724), .I3(n3725), .I4(n3726), .O(n3722)
         );
  NAND_GATE U4717 ( .I1(n3464), .I2(\registres[28][3] ), .O(n3726) );
  NAND_GATE U4718 ( .I1(n3465), .I2(\registres[29][3] ), .O(n3725) );
  NAND_GATE U4719 ( .I1(n3466), .I2(\registres[12][3] ), .O(n3724) );
  NAND_GATE U4720 ( .I1(n3467), .I2(\registres[20][3] ), .O(n3723) );
  NAND_GATE U4721 ( .I1(n3468), .I2(\registres[1][3] ), .O(n3721) );
  NAND_GATE U4722 ( .I1(n3469), .I2(\registres[9][3] ), .O(n3720) );
  NAND_GATE U4723 ( .I1(n3470), .I2(\registres[11][3] ), .O(n3719) );
  NAND_GATE U4724 ( .I1(n3471), .I2(\registres[13][3] ), .O(n3718) );
  AND5_GATE U4725 ( .I1(n3727), .I2(n3728), .I3(n3729), .I4(n3730), .I5(n3731), 
        .O(n3706) );
  AND4_GATE U4726 ( .I1(n3732), .I2(n3733), .I3(n3734), .I4(n3735), .O(n3731)
         );
  NAND_GATE U4727 ( .I1(n3481), .I2(\registres[17][3] ), .O(n3735) );
  NAND_GATE U4728 ( .I1(n3482), .I2(\registres[19][3] ), .O(n3734) );
  NAND_GATE U4729 ( .I1(n3483), .I2(\registres[21][3] ), .O(n3733) );
  NAND_GATE U4730 ( .I1(n3484), .I2(\registres[6][3] ), .O(n3732) );
  NAND_GATE U4731 ( .I1(n3485), .I2(\registres[7][3] ), .O(n3730) );
  NAND_GATE U4732 ( .I1(n3486), .I2(\registres[30][3] ), .O(n3729) );
  NAND_GATE U4733 ( .I1(n3487), .I2(\registres[31][3] ), .O(n3728) );
  NAND_GATE U4734 ( .I1(n3488), .I2(\registres[14][3] ), .O(n3727) );
  AND4_GATE U4735 ( .I1(n3736), .I2(n3737), .I3(n3738), .I4(n3739), .O(n3705)
         );
  AND4_GATE U4736 ( .I1(n3740), .I2(n3741), .I3(n3742), .I4(n3743), .O(n3739)
         );
  NAND_GATE U4737 ( .I1(n3497), .I2(\registres[22][3] ), .O(n3743) );
  NAND_GATE U4738 ( .I1(n3498), .I2(\registres[15][3] ), .O(n3742) );
  NAND_GATE U4739 ( .I1(n3499), .I2(\registres[23][3] ), .O(n3741) );
  NAND_GATE U4740 ( .I1(n3500), .I2(\registres[4][3] ), .O(n3740) );
  NAND_GATE U4741 ( .I1(n3501), .I2(\registres[8][3] ), .O(n3738) );
  NAND_GATE U4742 ( .I1(n3502), .I2(\registres[2][3] ), .O(n3737) );
  NAND_GATE U4743 ( .I1(n3503), .I2(\registres[16][3] ), .O(n3736) );
  AND_GATE U4744 ( .I1(n3744), .I2(n3432), .O(data_src1[31]) );
  NAND4_GATE U4745 ( .I1(n3745), .I2(n3746), .I3(n3747), .I4(n3748), .O(n3744)
         );
  AND5_GATE U4746 ( .I1(n3749), .I2(n3750), .I3(n3751), .I4(n3752), .I5(n3753), 
        .O(n3748) );
  AND4_GATE U4747 ( .I1(n3754), .I2(n3755), .I3(n3756), .I4(n3757), .O(n3753)
         );
  NAND_GATE U4748 ( .I1(n3447), .I2(\registres[24][31] ), .O(n3757) );
  NAND_GATE U4749 ( .I1(n3448), .I2(\registres[25][31] ), .O(n3756) );
  NAND_GATE U4750 ( .I1(n3449), .I2(\registres[3][31] ), .O(n3755) );
  NAND_GATE U4751 ( .I1(n3450), .I2(\registres[26][31] ), .O(n3754) );
  NAND_GATE U4752 ( .I1(n3451), .I2(\registres[27][31] ), .O(n3752) );
  NAND_GATE U4753 ( .I1(n3452), .I2(\registres[10][31] ), .O(n3751) );
  NAND_GATE U4754 ( .I1(n3453), .I2(\registres[18][31] ), .O(n3750) );
  NAND_GATE U4755 ( .I1(n3454), .I2(\registres[5][31] ), .O(n3749) );
  AND5_GATE U4756 ( .I1(n3758), .I2(n3759), .I3(n3760), .I4(n3761), .I5(n3762), 
        .O(n3747) );
  AND4_GATE U4757 ( .I1(n3763), .I2(n3764), .I3(n3765), .I4(n3766), .O(n3762)
         );
  NAND_GATE U4758 ( .I1(n3464), .I2(\registres[28][31] ), .O(n3766) );
  NAND_GATE U4759 ( .I1(n3465), .I2(\registres[29][31] ), .O(n3765) );
  NAND_GATE U4760 ( .I1(n3466), .I2(\registres[12][31] ), .O(n3764) );
  NAND_GATE U4761 ( .I1(n3467), .I2(\registres[20][31] ), .O(n3763) );
  NAND_GATE U4762 ( .I1(n3468), .I2(\registres[1][31] ), .O(n3761) );
  NAND_GATE U4763 ( .I1(n3469), .I2(\registres[9][31] ), .O(n3760) );
  NAND_GATE U4764 ( .I1(n3470), .I2(\registres[11][31] ), .O(n3759) );
  NAND_GATE U4765 ( .I1(n3471), .I2(\registres[13][31] ), .O(n3758) );
  AND5_GATE U4766 ( .I1(n3767), .I2(n3768), .I3(n3769), .I4(n3770), .I5(n3771), 
        .O(n3746) );
  AND4_GATE U4767 ( .I1(n3772), .I2(n3773), .I3(n3774), .I4(n3775), .O(n3771)
         );
  NAND_GATE U4768 ( .I1(n3481), .I2(\registres[17][31] ), .O(n3775) );
  NAND_GATE U4769 ( .I1(n3482), .I2(\registres[19][31] ), .O(n3774) );
  NAND_GATE U4770 ( .I1(n3483), .I2(\registres[21][31] ), .O(n3773) );
  NAND_GATE U4771 ( .I1(n3484), .I2(\registres[6][31] ), .O(n3772) );
  NAND_GATE U4772 ( .I1(n3485), .I2(\registres[7][31] ), .O(n3770) );
  NAND_GATE U4773 ( .I1(n3486), .I2(\registres[30][31] ), .O(n3769) );
  NAND_GATE U4774 ( .I1(n3487), .I2(\registres[31][31] ), .O(n3768) );
  NAND_GATE U4775 ( .I1(n3488), .I2(\registres[14][31] ), .O(n3767) );
  AND4_GATE U4776 ( .I1(n3776), .I2(n3777), .I3(n3778), .I4(n3779), .O(n3745)
         );
  AND4_GATE U4777 ( .I1(n3780), .I2(n3781), .I3(n3782), .I4(n3783), .O(n3779)
         );
  NAND_GATE U4778 ( .I1(n3497), .I2(\registres[22][31] ), .O(n3783) );
  NAND_GATE U4779 ( .I1(n3498), .I2(\registres[15][31] ), .O(n3782) );
  NAND_GATE U4780 ( .I1(n3499), .I2(\registres[23][31] ), .O(n3781) );
  NAND_GATE U4781 ( .I1(n3500), .I2(\registres[4][31] ), .O(n3780) );
  NAND_GATE U4782 ( .I1(n3501), .I2(\registres[8][31] ), .O(n3778) );
  NAND_GATE U4783 ( .I1(n3502), .I2(\registres[2][31] ), .O(n3777) );
  NAND_GATE U4784 ( .I1(n3503), .I2(\registres[16][31] ), .O(n3776) );
  AND_GATE U4785 ( .I1(n3784), .I2(n3432), .O(data_src1[30]) );
  NAND4_GATE U4786 ( .I1(n3785), .I2(n3786), .I3(n3787), .I4(n3788), .O(n3784)
         );
  AND5_GATE U4787 ( .I1(n3789), .I2(n3790), .I3(n3791), .I4(n3792), .I5(n3793), 
        .O(n3788) );
  AND4_GATE U4788 ( .I1(n3794), .I2(n3795), .I3(n3796), .I4(n3797), .O(n3793)
         );
  NAND_GATE U4789 ( .I1(n3447), .I2(\registres[24][30] ), .O(n3797) );
  NAND_GATE U4790 ( .I1(n3448), .I2(\registres[25][30] ), .O(n3796) );
  NAND_GATE U4791 ( .I1(n3449), .I2(\registres[3][30] ), .O(n3795) );
  NAND_GATE U4792 ( .I1(n3450), .I2(\registres[26][30] ), .O(n3794) );
  NAND_GATE U4793 ( .I1(n3451), .I2(\registres[27][30] ), .O(n3792) );
  NAND_GATE U4794 ( .I1(n3452), .I2(\registres[10][30] ), .O(n3791) );
  NAND_GATE U4795 ( .I1(n3453), .I2(\registres[18][30] ), .O(n3790) );
  NAND_GATE U4796 ( .I1(n3454), .I2(\registres[5][30] ), .O(n3789) );
  AND5_GATE U4797 ( .I1(n3798), .I2(n3799), .I3(n3800), .I4(n3801), .I5(n3802), 
        .O(n3787) );
  AND4_GATE U4798 ( .I1(n3803), .I2(n3804), .I3(n3805), .I4(n3806), .O(n3802)
         );
  NAND_GATE U4799 ( .I1(n3464), .I2(\registres[28][30] ), .O(n3806) );
  NAND_GATE U4800 ( .I1(n3465), .I2(\registres[29][30] ), .O(n3805) );
  NAND_GATE U4801 ( .I1(n3466), .I2(\registres[12][30] ), .O(n3804) );
  NAND_GATE U4802 ( .I1(n3467), .I2(\registres[20][30] ), .O(n3803) );
  NAND_GATE U4803 ( .I1(n3468), .I2(\registres[1][30] ), .O(n3801) );
  NAND_GATE U4804 ( .I1(n3469), .I2(\registres[9][30] ), .O(n3800) );
  NAND_GATE U4805 ( .I1(n3470), .I2(\registres[11][30] ), .O(n3799) );
  NAND_GATE U4806 ( .I1(n3471), .I2(\registres[13][30] ), .O(n3798) );
  AND5_GATE U4807 ( .I1(n3807), .I2(n3808), .I3(n3809), .I4(n3810), .I5(n3811), 
        .O(n3786) );
  AND4_GATE U4808 ( .I1(n3812), .I2(n3813), .I3(n3814), .I4(n3815), .O(n3811)
         );
  NAND_GATE U4809 ( .I1(n3481), .I2(\registres[17][30] ), .O(n3815) );
  NAND_GATE U4810 ( .I1(n3482), .I2(\registres[19][30] ), .O(n3814) );
  NAND_GATE U4811 ( .I1(n3483), .I2(\registres[21][30] ), .O(n3813) );
  NAND_GATE U4812 ( .I1(n3484), .I2(\registres[6][30] ), .O(n3812) );
  NAND_GATE U4813 ( .I1(n3485), .I2(\registres[7][30] ), .O(n3810) );
  NAND_GATE U4814 ( .I1(n3486), .I2(\registres[30][30] ), .O(n3809) );
  NAND_GATE U4815 ( .I1(n3487), .I2(\registres[31][30] ), .O(n3808) );
  NAND_GATE U4816 ( .I1(n3488), .I2(\registres[14][30] ), .O(n3807) );
  AND4_GATE U4817 ( .I1(n3816), .I2(n3817), .I3(n3818), .I4(n3819), .O(n3785)
         );
  AND4_GATE U4818 ( .I1(n3820), .I2(n3821), .I3(n3822), .I4(n3823), .O(n3819)
         );
  NAND_GATE U4819 ( .I1(n3497), .I2(\registres[22][30] ), .O(n3823) );
  NAND_GATE U4820 ( .I1(n3498), .I2(\registres[15][30] ), .O(n3822) );
  NAND_GATE U4821 ( .I1(n3499), .I2(\registres[23][30] ), .O(n3821) );
  NAND_GATE U4822 ( .I1(n3500), .I2(\registres[4][30] ), .O(n3820) );
  NAND_GATE U4823 ( .I1(n3501), .I2(\registres[8][30] ), .O(n3818) );
  NAND_GATE U4824 ( .I1(n3502), .I2(\registres[2][30] ), .O(n3817) );
  NAND_GATE U4825 ( .I1(n3503), .I2(\registres[16][30] ), .O(n3816) );
  AND_GATE U4826 ( .I1(n3824), .I2(n3432), .O(data_src1[2]) );
  NAND4_GATE U4827 ( .I1(n3825), .I2(n3826), .I3(n3827), .I4(n3828), .O(n3824)
         );
  AND5_GATE U4828 ( .I1(n3829), .I2(n3830), .I3(n3831), .I4(n3832), .I5(n3833), 
        .O(n3828) );
  AND4_GATE U4829 ( .I1(n3834), .I2(n3835), .I3(n3836), .I4(n3837), .O(n3833)
         );
  NAND_GATE U4830 ( .I1(n3447), .I2(\registres[24][2] ), .O(n3837) );
  NAND_GATE U4831 ( .I1(n3448), .I2(\registres[25][2] ), .O(n3836) );
  NAND_GATE U4832 ( .I1(n3449), .I2(\registres[3][2] ), .O(n3835) );
  NAND_GATE U4833 ( .I1(n3450), .I2(\registres[26][2] ), .O(n3834) );
  NAND_GATE U4834 ( .I1(n3451), .I2(\registres[27][2] ), .O(n3832) );
  NAND_GATE U4835 ( .I1(n3452), .I2(\registres[10][2] ), .O(n3831) );
  NAND_GATE U4836 ( .I1(n3453), .I2(\registres[18][2] ), .O(n3830) );
  NAND_GATE U4837 ( .I1(n3454), .I2(\registres[5][2] ), .O(n3829) );
  AND5_GATE U4838 ( .I1(n3838), .I2(n3839), .I3(n3840), .I4(n3841), .I5(n3842), 
        .O(n3827) );
  AND4_GATE U4839 ( .I1(n3843), .I2(n3844), .I3(n3845), .I4(n3846), .O(n3842)
         );
  NAND_GATE U4840 ( .I1(n3464), .I2(\registres[28][2] ), .O(n3846) );
  NAND_GATE U4841 ( .I1(n3465), .I2(\registres[29][2] ), .O(n3845) );
  NAND_GATE U4842 ( .I1(n3466), .I2(\registres[12][2] ), .O(n3844) );
  NAND_GATE U4843 ( .I1(n3467), .I2(\registres[20][2] ), .O(n3843) );
  NAND_GATE U4844 ( .I1(n3468), .I2(\registres[1][2] ), .O(n3841) );
  NAND_GATE U4845 ( .I1(n3469), .I2(\registres[9][2] ), .O(n3840) );
  NAND_GATE U4846 ( .I1(n3470), .I2(\registres[11][2] ), .O(n3839) );
  NAND_GATE U4847 ( .I1(n3471), .I2(\registres[13][2] ), .O(n3838) );
  AND5_GATE U4848 ( .I1(n3847), .I2(n3848), .I3(n3849), .I4(n3850), .I5(n3851), 
        .O(n3826) );
  AND4_GATE U4849 ( .I1(n3852), .I2(n3853), .I3(n3854), .I4(n3855), .O(n3851)
         );
  NAND_GATE U4850 ( .I1(n3481), .I2(\registres[17][2] ), .O(n3855) );
  NAND_GATE U4851 ( .I1(n3482), .I2(\registres[19][2] ), .O(n3854) );
  NAND_GATE U4852 ( .I1(n3483), .I2(\registres[21][2] ), .O(n3853) );
  NAND_GATE U4853 ( .I1(n3484), .I2(\registres[6][2] ), .O(n3852) );
  NAND_GATE U4854 ( .I1(n3485), .I2(\registres[7][2] ), .O(n3850) );
  NAND_GATE U4855 ( .I1(n3486), .I2(\registres[30][2] ), .O(n3849) );
  NAND_GATE U4856 ( .I1(n3487), .I2(\registres[31][2] ), .O(n3848) );
  NAND_GATE U4857 ( .I1(n3488), .I2(\registres[14][2] ), .O(n3847) );
  AND4_GATE U4858 ( .I1(n3856), .I2(n3857), .I3(n3858), .I4(n3859), .O(n3825)
         );
  AND4_GATE U4859 ( .I1(n3860), .I2(n3861), .I3(n3862), .I4(n3863), .O(n3859)
         );
  NAND_GATE U4860 ( .I1(n3497), .I2(\registres[22][2] ), .O(n3863) );
  NAND_GATE U4861 ( .I1(n3498), .I2(\registres[15][2] ), .O(n3862) );
  NAND_GATE U4862 ( .I1(n3499), .I2(\registres[23][2] ), .O(n3861) );
  NAND_GATE U4863 ( .I1(n3500), .I2(\registres[4][2] ), .O(n3860) );
  NAND_GATE U4864 ( .I1(n3501), .I2(\registres[8][2] ), .O(n3858) );
  NAND_GATE U4865 ( .I1(n3502), .I2(\registres[2][2] ), .O(n3857) );
  NAND_GATE U4866 ( .I1(n3503), .I2(\registres[16][2] ), .O(n3856) );
  AND_GATE U4867 ( .I1(n3864), .I2(n3432), .O(data_src1[29]) );
  NAND4_GATE U4868 ( .I1(n3865), .I2(n3866), .I3(n3867), .I4(n3868), .O(n3864)
         );
  AND5_GATE U4869 ( .I1(n3869), .I2(n3870), .I3(n3871), .I4(n3872), .I5(n3873), 
        .O(n3868) );
  AND4_GATE U4870 ( .I1(n3874), .I2(n3875), .I3(n3876), .I4(n3877), .O(n3873)
         );
  NAND_GATE U4871 ( .I1(n3447), .I2(\registres[24][29] ), .O(n3877) );
  NAND_GATE U4872 ( .I1(n3448), .I2(\registres[25][29] ), .O(n3876) );
  NAND_GATE U4873 ( .I1(n3449), .I2(\registres[3][29] ), .O(n3875) );
  NAND_GATE U4874 ( .I1(n3450), .I2(\registres[26][29] ), .O(n3874) );
  NAND_GATE U4875 ( .I1(n3451), .I2(\registres[27][29] ), .O(n3872) );
  NAND_GATE U4876 ( .I1(n3452), .I2(\registres[10][29] ), .O(n3871) );
  NAND_GATE U4877 ( .I1(n3453), .I2(\registres[18][29] ), .O(n3870) );
  NAND_GATE U4878 ( .I1(n3454), .I2(\registres[5][29] ), .O(n3869) );
  AND5_GATE U4879 ( .I1(n3878), .I2(n3879), .I3(n3880), .I4(n3881), .I5(n3882), 
        .O(n3867) );
  AND4_GATE U4880 ( .I1(n3883), .I2(n3884), .I3(n3885), .I4(n3886), .O(n3882)
         );
  NAND_GATE U4881 ( .I1(n3464), .I2(\registres[28][29] ), .O(n3886) );
  NAND_GATE U4882 ( .I1(n3465), .I2(\registres[29][29] ), .O(n3885) );
  NAND_GATE U4883 ( .I1(n3466), .I2(\registres[12][29] ), .O(n3884) );
  NAND_GATE U4884 ( .I1(n3467), .I2(\registres[20][29] ), .O(n3883) );
  NAND_GATE U4885 ( .I1(n3468), .I2(\registres[1][29] ), .O(n3881) );
  NAND_GATE U4886 ( .I1(n3469), .I2(\registres[9][29] ), .O(n3880) );
  NAND_GATE U4887 ( .I1(n3470), .I2(\registres[11][29] ), .O(n3879) );
  NAND_GATE U4888 ( .I1(n3471), .I2(\registres[13][29] ), .O(n3878) );
  AND5_GATE U4889 ( .I1(n3887), .I2(n3888), .I3(n3889), .I4(n3890), .I5(n3891), 
        .O(n3866) );
  AND4_GATE U4890 ( .I1(n3892), .I2(n3893), .I3(n3894), .I4(n3895), .O(n3891)
         );
  NAND_GATE U4891 ( .I1(n3481), .I2(\registres[17][29] ), .O(n3895) );
  NAND_GATE U4892 ( .I1(n3482), .I2(\registres[19][29] ), .O(n3894) );
  NAND_GATE U4893 ( .I1(n3483), .I2(\registres[21][29] ), .O(n3893) );
  NAND_GATE U4894 ( .I1(n3484), .I2(\registres[6][29] ), .O(n3892) );
  NAND_GATE U4895 ( .I1(n3485), .I2(\registres[7][29] ), .O(n3890) );
  NAND_GATE U4896 ( .I1(n3486), .I2(\registres[30][29] ), .O(n3889) );
  NAND_GATE U4897 ( .I1(n3487), .I2(\registres[31][29] ), .O(n3888) );
  NAND_GATE U4898 ( .I1(n3488), .I2(\registres[14][29] ), .O(n3887) );
  AND4_GATE U4899 ( .I1(n3896), .I2(n3897), .I3(n3898), .I4(n3899), .O(n3865)
         );
  AND4_GATE U4900 ( .I1(n3900), .I2(n3901), .I3(n3902), .I4(n3903), .O(n3899)
         );
  NAND_GATE U4901 ( .I1(n3497), .I2(\registres[22][29] ), .O(n3903) );
  NAND_GATE U4902 ( .I1(n3498), .I2(\registres[15][29] ), .O(n3902) );
  NAND_GATE U4903 ( .I1(n3499), .I2(\registres[23][29] ), .O(n3901) );
  NAND_GATE U4904 ( .I1(n3500), .I2(\registres[4][29] ), .O(n3900) );
  NAND_GATE U4905 ( .I1(n3501), .I2(\registres[8][29] ), .O(n3898) );
  NAND_GATE U4906 ( .I1(n3502), .I2(\registres[2][29] ), .O(n3897) );
  NAND_GATE U4907 ( .I1(n3503), .I2(\registres[16][29] ), .O(n3896) );
  AND_GATE U4908 ( .I1(n3904), .I2(n3432), .O(data_src1[28]) );
  NAND4_GATE U4909 ( .I1(n3905), .I2(n3906), .I3(n3907), .I4(n3908), .O(n3904)
         );
  AND5_GATE U4910 ( .I1(n3909), .I2(n3910), .I3(n3911), .I4(n3912), .I5(n3913), 
        .O(n3908) );
  AND4_GATE U4911 ( .I1(n3914), .I2(n3915), .I3(n3916), .I4(n3917), .O(n3913)
         );
  NAND_GATE U4912 ( .I1(n3447), .I2(\registres[24][28] ), .O(n3917) );
  NAND_GATE U4913 ( .I1(n3448), .I2(\registres[25][28] ), .O(n3916) );
  NAND_GATE U4914 ( .I1(n3449), .I2(\registres[3][28] ), .O(n3915) );
  NAND_GATE U4915 ( .I1(n3450), .I2(\registres[26][28] ), .O(n3914) );
  NAND_GATE U4916 ( .I1(n3451), .I2(\registres[27][28] ), .O(n3912) );
  NAND_GATE U4917 ( .I1(n3452), .I2(\registres[10][28] ), .O(n3911) );
  NAND_GATE U4918 ( .I1(n3453), .I2(\registres[18][28] ), .O(n3910) );
  NAND_GATE U4919 ( .I1(n3454), .I2(\registres[5][28] ), .O(n3909) );
  AND5_GATE U4920 ( .I1(n3918), .I2(n3919), .I3(n3920), .I4(n3921), .I5(n3922), 
        .O(n3907) );
  AND4_GATE U4921 ( .I1(n3923), .I2(n3924), .I3(n3925), .I4(n3926), .O(n3922)
         );
  NAND_GATE U4922 ( .I1(n3464), .I2(\registres[28][28] ), .O(n3926) );
  NAND_GATE U4923 ( .I1(n3465), .I2(\registres[29][28] ), .O(n3925) );
  NAND_GATE U4924 ( .I1(n3466), .I2(\registres[12][28] ), .O(n3924) );
  NAND_GATE U4925 ( .I1(n3467), .I2(\registres[20][28] ), .O(n3923) );
  NAND_GATE U4926 ( .I1(n3468), .I2(\registres[1][28] ), .O(n3921) );
  NAND_GATE U4927 ( .I1(n3469), .I2(\registres[9][28] ), .O(n3920) );
  NAND_GATE U4928 ( .I1(n3470), .I2(\registres[11][28] ), .O(n3919) );
  NAND_GATE U4929 ( .I1(n3471), .I2(\registres[13][28] ), .O(n3918) );
  AND5_GATE U4930 ( .I1(n3927), .I2(n3928), .I3(n3929), .I4(n3930), .I5(n3931), 
        .O(n3906) );
  AND4_GATE U4931 ( .I1(n3932), .I2(n3933), .I3(n3934), .I4(n3935), .O(n3931)
         );
  NAND_GATE U4932 ( .I1(n3481), .I2(\registres[17][28] ), .O(n3935) );
  NAND_GATE U4933 ( .I1(n3482), .I2(\registres[19][28] ), .O(n3934) );
  NAND_GATE U4934 ( .I1(n3483), .I2(\registres[21][28] ), .O(n3933) );
  NAND_GATE U4935 ( .I1(n3484), .I2(\registres[6][28] ), .O(n3932) );
  NAND_GATE U4936 ( .I1(n3485), .I2(\registres[7][28] ), .O(n3930) );
  NAND_GATE U4937 ( .I1(n3486), .I2(\registres[30][28] ), .O(n3929) );
  NAND_GATE U4938 ( .I1(n3487), .I2(\registres[31][28] ), .O(n3928) );
  NAND_GATE U4939 ( .I1(n3488), .I2(\registres[14][28] ), .O(n3927) );
  AND4_GATE U4940 ( .I1(n3936), .I2(n3937), .I3(n3938), .I4(n3939), .O(n3905)
         );
  AND4_GATE U4941 ( .I1(n3940), .I2(n3941), .I3(n3942), .I4(n3943), .O(n3939)
         );
  NAND_GATE U4942 ( .I1(n3497), .I2(\registres[22][28] ), .O(n3943) );
  NAND_GATE U4943 ( .I1(n3498), .I2(\registres[15][28] ), .O(n3942) );
  NAND_GATE U4944 ( .I1(n3499), .I2(\registres[23][28] ), .O(n3941) );
  NAND_GATE U4945 ( .I1(n3500), .I2(\registres[4][28] ), .O(n3940) );
  NAND_GATE U4946 ( .I1(n3501), .I2(\registres[8][28] ), .O(n3938) );
  NAND_GATE U4947 ( .I1(n3502), .I2(\registres[2][28] ), .O(n3937) );
  NAND_GATE U4948 ( .I1(n3503), .I2(\registres[16][28] ), .O(n3936) );
  AND_GATE U4949 ( .I1(n3944), .I2(n3432), .O(data_src1[27]) );
  NAND4_GATE U4950 ( .I1(n3945), .I2(n3946), .I3(n3947), .I4(n3948), .O(n3944)
         );
  AND5_GATE U4951 ( .I1(n3949), .I2(n3950), .I3(n3951), .I4(n3952), .I5(n3953), 
        .O(n3948) );
  AND4_GATE U4952 ( .I1(n3954), .I2(n3955), .I3(n3956), .I4(n3957), .O(n3953)
         );
  NAND_GATE U4953 ( .I1(n3447), .I2(\registres[24][27] ), .O(n3957) );
  NAND_GATE U4954 ( .I1(n3448), .I2(\registres[25][27] ), .O(n3956) );
  NAND_GATE U4955 ( .I1(n3449), .I2(\registres[3][27] ), .O(n3955) );
  NAND_GATE U4956 ( .I1(n3450), .I2(\registres[26][27] ), .O(n3954) );
  NAND_GATE U4957 ( .I1(n3451), .I2(\registres[27][27] ), .O(n3952) );
  NAND_GATE U4958 ( .I1(n3452), .I2(\registres[10][27] ), .O(n3951) );
  NAND_GATE U4959 ( .I1(n3453), .I2(\registres[18][27] ), .O(n3950) );
  NAND_GATE U4960 ( .I1(n3454), .I2(\registres[5][27] ), .O(n3949) );
  AND5_GATE U4961 ( .I1(n3958), .I2(n3959), .I3(n3960), .I4(n3961), .I5(n3962), 
        .O(n3947) );
  AND4_GATE U4962 ( .I1(n3963), .I2(n3964), .I3(n3965), .I4(n3966), .O(n3962)
         );
  NAND_GATE U4963 ( .I1(n3464), .I2(\registres[28][27] ), .O(n3966) );
  NAND_GATE U4964 ( .I1(n3465), .I2(\registres[29][27] ), .O(n3965) );
  NAND_GATE U4965 ( .I1(n3466), .I2(\registres[12][27] ), .O(n3964) );
  NAND_GATE U4966 ( .I1(n3467), .I2(\registres[20][27] ), .O(n3963) );
  NAND_GATE U4967 ( .I1(n3468), .I2(\registres[1][27] ), .O(n3961) );
  NAND_GATE U4968 ( .I1(n3469), .I2(\registres[9][27] ), .O(n3960) );
  NAND_GATE U4969 ( .I1(n3470), .I2(\registres[11][27] ), .O(n3959) );
  NAND_GATE U4970 ( .I1(n3471), .I2(\registres[13][27] ), .O(n3958) );
  AND5_GATE U4971 ( .I1(n3967), .I2(n3968), .I3(n3969), .I4(n3970), .I5(n3971), 
        .O(n3946) );
  AND4_GATE U4972 ( .I1(n3972), .I2(n3973), .I3(n3974), .I4(n3975), .O(n3971)
         );
  NAND_GATE U4973 ( .I1(n3481), .I2(\registres[17][27] ), .O(n3975) );
  NAND_GATE U4974 ( .I1(n3482), .I2(\registres[19][27] ), .O(n3974) );
  NAND_GATE U4975 ( .I1(n3483), .I2(\registres[21][27] ), .O(n3973) );
  NAND_GATE U4976 ( .I1(n3484), .I2(\registres[6][27] ), .O(n3972) );
  NAND_GATE U4977 ( .I1(n3485), .I2(\registres[7][27] ), .O(n3970) );
  NAND_GATE U4978 ( .I1(n3486), .I2(\registres[30][27] ), .O(n3969) );
  NAND_GATE U4979 ( .I1(n3487), .I2(\registres[31][27] ), .O(n3968) );
  NAND_GATE U4980 ( .I1(n3488), .I2(\registres[14][27] ), .O(n3967) );
  AND4_GATE U4981 ( .I1(n3976), .I2(n3977), .I3(n3978), .I4(n3979), .O(n3945)
         );
  AND4_GATE U4982 ( .I1(n3980), .I2(n3981), .I3(n3982), .I4(n3983), .O(n3979)
         );
  NAND_GATE U4983 ( .I1(n3497), .I2(\registres[22][27] ), .O(n3983) );
  NAND_GATE U4984 ( .I1(n3498), .I2(\registres[15][27] ), .O(n3982) );
  NAND_GATE U4985 ( .I1(n3499), .I2(\registres[23][27] ), .O(n3981) );
  NAND_GATE U4986 ( .I1(n3500), .I2(\registres[4][27] ), .O(n3980) );
  NAND_GATE U4987 ( .I1(n3501), .I2(\registres[8][27] ), .O(n3978) );
  NAND_GATE U4988 ( .I1(n3502), .I2(\registres[2][27] ), .O(n3977) );
  NAND_GATE U4989 ( .I1(n3503), .I2(\registres[16][27] ), .O(n3976) );
  AND_GATE U4990 ( .I1(n3984), .I2(n3432), .O(data_src1[26]) );
  NAND4_GATE U4991 ( .I1(n3985), .I2(n3986), .I3(n3987), .I4(n3988), .O(n3984)
         );
  AND5_GATE U4992 ( .I1(n3989), .I2(n3990), .I3(n3991), .I4(n3992), .I5(n3993), 
        .O(n3988) );
  AND4_GATE U4993 ( .I1(n3994), .I2(n3995), .I3(n3996), .I4(n3997), .O(n3993)
         );
  NAND_GATE U4994 ( .I1(n3447), .I2(\registres[24][26] ), .O(n3997) );
  NAND_GATE U4995 ( .I1(n3448), .I2(\registres[25][26] ), .O(n3996) );
  NAND_GATE U4996 ( .I1(n3449), .I2(\registres[3][26] ), .O(n3995) );
  NAND_GATE U4997 ( .I1(n3450), .I2(\registres[26][26] ), .O(n3994) );
  NAND_GATE U4998 ( .I1(n3451), .I2(\registres[27][26] ), .O(n3992) );
  NAND_GATE U4999 ( .I1(n3452), .I2(\registres[10][26] ), .O(n3991) );
  NAND_GATE U5000 ( .I1(n3453), .I2(\registres[18][26] ), .O(n3990) );
  NAND_GATE U5001 ( .I1(n3454), .I2(\registres[5][26] ), .O(n3989) );
  AND5_GATE U5002 ( .I1(n3998), .I2(n3999), .I3(n4000), .I4(n4001), .I5(n4002), 
        .O(n3987) );
  AND4_GATE U5003 ( .I1(n4003), .I2(n4004), .I3(n4005), .I4(n4006), .O(n4002)
         );
  NAND_GATE U5004 ( .I1(n3464), .I2(\registres[28][26] ), .O(n4006) );
  NAND_GATE U5005 ( .I1(n3465), .I2(\registres[29][26] ), .O(n4005) );
  NAND_GATE U5006 ( .I1(n3466), .I2(\registres[12][26] ), .O(n4004) );
  NAND_GATE U5007 ( .I1(n3467), .I2(\registres[20][26] ), .O(n4003) );
  NAND_GATE U5008 ( .I1(n3468), .I2(\registres[1][26] ), .O(n4001) );
  NAND_GATE U5009 ( .I1(n3469), .I2(\registres[9][26] ), .O(n4000) );
  NAND_GATE U5010 ( .I1(n3470), .I2(\registres[11][26] ), .O(n3999) );
  NAND_GATE U5011 ( .I1(n3471), .I2(\registres[13][26] ), .O(n3998) );
  AND5_GATE U5012 ( .I1(n4007), .I2(n4008), .I3(n4009), .I4(n4010), .I5(n4011), 
        .O(n3986) );
  AND4_GATE U5013 ( .I1(n4012), .I2(n4013), .I3(n4014), .I4(n4015), .O(n4011)
         );
  NAND_GATE U5014 ( .I1(n3481), .I2(\registres[17][26] ), .O(n4015) );
  NAND_GATE U5015 ( .I1(n3482), .I2(\registres[19][26] ), .O(n4014) );
  NAND_GATE U5016 ( .I1(n3483), .I2(\registres[21][26] ), .O(n4013) );
  NAND_GATE U5017 ( .I1(n3484), .I2(\registres[6][26] ), .O(n4012) );
  NAND_GATE U5018 ( .I1(n3485), .I2(\registres[7][26] ), .O(n4010) );
  NAND_GATE U5019 ( .I1(n3486), .I2(\registres[30][26] ), .O(n4009) );
  NAND_GATE U5020 ( .I1(n3487), .I2(\registres[31][26] ), .O(n4008) );
  NAND_GATE U5021 ( .I1(n3488), .I2(\registres[14][26] ), .O(n4007) );
  AND4_GATE U5022 ( .I1(n4016), .I2(n4017), .I3(n4018), .I4(n4019), .O(n3985)
         );
  AND4_GATE U5023 ( .I1(n4020), .I2(n4021), .I3(n4022), .I4(n4023), .O(n4019)
         );
  NAND_GATE U5024 ( .I1(n3497), .I2(\registres[22][26] ), .O(n4023) );
  NAND_GATE U5025 ( .I1(n3498), .I2(\registres[15][26] ), .O(n4022) );
  NAND_GATE U5026 ( .I1(n3499), .I2(\registres[23][26] ), .O(n4021) );
  NAND_GATE U5027 ( .I1(n3500), .I2(\registres[4][26] ), .O(n4020) );
  NAND_GATE U5028 ( .I1(n3501), .I2(\registres[8][26] ), .O(n4018) );
  NAND_GATE U5029 ( .I1(n3502), .I2(\registres[2][26] ), .O(n4017) );
  NAND_GATE U5030 ( .I1(n3503), .I2(\registres[16][26] ), .O(n4016) );
  AND_GATE U5031 ( .I1(n4024), .I2(n3432), .O(data_src1[25]) );
  NAND4_GATE U5032 ( .I1(n4025), .I2(n4026), .I3(n4027), .I4(n4028), .O(n4024)
         );
  AND5_GATE U5033 ( .I1(n4029), .I2(n4030), .I3(n4031), .I4(n4032), .I5(n4033), 
        .O(n4028) );
  AND4_GATE U5034 ( .I1(n4034), .I2(n4035), .I3(n4036), .I4(n4037), .O(n4033)
         );
  NAND_GATE U5035 ( .I1(n3447), .I2(\registres[24][25] ), .O(n4037) );
  NAND_GATE U5036 ( .I1(n3448), .I2(\registres[25][25] ), .O(n4036) );
  NAND_GATE U5037 ( .I1(n3449), .I2(\registres[3][25] ), .O(n4035) );
  NAND_GATE U5038 ( .I1(n3450), .I2(\registres[26][25] ), .O(n4034) );
  NAND_GATE U5039 ( .I1(n3451), .I2(\registres[27][25] ), .O(n4032) );
  NAND_GATE U5040 ( .I1(n3452), .I2(\registres[10][25] ), .O(n4031) );
  NAND_GATE U5041 ( .I1(n3453), .I2(\registres[18][25] ), .O(n4030) );
  NAND_GATE U5042 ( .I1(n3454), .I2(\registres[5][25] ), .O(n4029) );
  AND5_GATE U5043 ( .I1(n4038), .I2(n4039), .I3(n4040), .I4(n4041), .I5(n4042), 
        .O(n4027) );
  AND4_GATE U5044 ( .I1(n4043), .I2(n4044), .I3(n4045), .I4(n4046), .O(n4042)
         );
  NAND_GATE U5045 ( .I1(n3464), .I2(\registres[28][25] ), .O(n4046) );
  NAND_GATE U5046 ( .I1(n3465), .I2(\registres[29][25] ), .O(n4045) );
  NAND_GATE U5047 ( .I1(n3466), .I2(\registres[12][25] ), .O(n4044) );
  NAND_GATE U5048 ( .I1(n3467), .I2(\registres[20][25] ), .O(n4043) );
  NAND_GATE U5049 ( .I1(n3468), .I2(\registres[1][25] ), .O(n4041) );
  NAND_GATE U5050 ( .I1(n3469), .I2(\registres[9][25] ), .O(n4040) );
  NAND_GATE U5051 ( .I1(n3470), .I2(\registres[11][25] ), .O(n4039) );
  NAND_GATE U5052 ( .I1(n3471), .I2(\registres[13][25] ), .O(n4038) );
  AND5_GATE U5053 ( .I1(n4047), .I2(n4048), .I3(n4049), .I4(n4050), .I5(n4051), 
        .O(n4026) );
  AND4_GATE U5054 ( .I1(n4052), .I2(n4053), .I3(n4054), .I4(n4055), .O(n4051)
         );
  NAND_GATE U5055 ( .I1(n3481), .I2(\registres[17][25] ), .O(n4055) );
  NAND_GATE U5056 ( .I1(n3482), .I2(\registres[19][25] ), .O(n4054) );
  NAND_GATE U5057 ( .I1(n3483), .I2(\registres[21][25] ), .O(n4053) );
  NAND_GATE U5058 ( .I1(n3484), .I2(\registres[6][25] ), .O(n4052) );
  NAND_GATE U5059 ( .I1(n3485), .I2(\registres[7][25] ), .O(n4050) );
  NAND_GATE U5060 ( .I1(n3486), .I2(\registres[30][25] ), .O(n4049) );
  NAND_GATE U5061 ( .I1(n3487), .I2(\registres[31][25] ), .O(n4048) );
  NAND_GATE U5062 ( .I1(n3488), .I2(\registres[14][25] ), .O(n4047) );
  AND4_GATE U5063 ( .I1(n4056), .I2(n4057), .I3(n4058), .I4(n4059), .O(n4025)
         );
  AND4_GATE U5064 ( .I1(n4060), .I2(n4061), .I3(n4062), .I4(n4063), .O(n4059)
         );
  NAND_GATE U5065 ( .I1(n3497), .I2(\registres[22][25] ), .O(n4063) );
  NAND_GATE U5066 ( .I1(n3498), .I2(\registres[15][25] ), .O(n4062) );
  NAND_GATE U5067 ( .I1(n3499), .I2(\registres[23][25] ), .O(n4061) );
  NAND_GATE U5068 ( .I1(n3500), .I2(\registres[4][25] ), .O(n4060) );
  NAND_GATE U5069 ( .I1(n3501), .I2(\registres[8][25] ), .O(n4058) );
  NAND_GATE U5070 ( .I1(n3502), .I2(\registres[2][25] ), .O(n4057) );
  NAND_GATE U5071 ( .I1(n3503), .I2(\registres[16][25] ), .O(n4056) );
  AND_GATE U5072 ( .I1(n4064), .I2(n3432), .O(data_src1[24]) );
  NAND4_GATE U5073 ( .I1(n4065), .I2(n4066), .I3(n4067), .I4(n4068), .O(n4064)
         );
  AND5_GATE U5074 ( .I1(n4069), .I2(n4070), .I3(n4071), .I4(n4072), .I5(n4073), 
        .O(n4068) );
  AND4_GATE U5075 ( .I1(n4074), .I2(n4075), .I3(n4076), .I4(n4077), .O(n4073)
         );
  NAND_GATE U5076 ( .I1(n3447), .I2(\registres[24][24] ), .O(n4077) );
  NAND_GATE U5077 ( .I1(n3448), .I2(\registres[25][24] ), .O(n4076) );
  NAND_GATE U5078 ( .I1(n3449), .I2(\registres[3][24] ), .O(n4075) );
  NAND_GATE U5079 ( .I1(n3450), .I2(\registres[26][24] ), .O(n4074) );
  NAND_GATE U5080 ( .I1(n3451), .I2(\registres[27][24] ), .O(n4072) );
  NAND_GATE U5081 ( .I1(n3452), .I2(\registres[10][24] ), .O(n4071) );
  NAND_GATE U5082 ( .I1(n3453), .I2(\registres[18][24] ), .O(n4070) );
  NAND_GATE U5083 ( .I1(n3454), .I2(\registres[5][24] ), .O(n4069) );
  AND5_GATE U5084 ( .I1(n4078), .I2(n4079), .I3(n4080), .I4(n4081), .I5(n4082), 
        .O(n4067) );
  AND4_GATE U5085 ( .I1(n4083), .I2(n4084), .I3(n4085), .I4(n4086), .O(n4082)
         );
  NAND_GATE U5086 ( .I1(n3464), .I2(\registres[28][24] ), .O(n4086) );
  NAND_GATE U5087 ( .I1(n3465), .I2(\registres[29][24] ), .O(n4085) );
  NAND_GATE U5088 ( .I1(n3466), .I2(\registres[12][24] ), .O(n4084) );
  NAND_GATE U5089 ( .I1(n3467), .I2(\registres[20][24] ), .O(n4083) );
  NAND_GATE U5090 ( .I1(n3468), .I2(\registres[1][24] ), .O(n4081) );
  NAND_GATE U5091 ( .I1(n3469), .I2(\registres[9][24] ), .O(n4080) );
  NAND_GATE U5092 ( .I1(n3470), .I2(\registres[11][24] ), .O(n4079) );
  NAND_GATE U5093 ( .I1(n3471), .I2(\registres[13][24] ), .O(n4078) );
  AND5_GATE U5094 ( .I1(n4087), .I2(n4088), .I3(n4089), .I4(n4090), .I5(n4091), 
        .O(n4066) );
  AND4_GATE U5095 ( .I1(n4092), .I2(n4093), .I3(n4094), .I4(n4095), .O(n4091)
         );
  NAND_GATE U5096 ( .I1(n3481), .I2(\registres[17][24] ), .O(n4095) );
  NAND_GATE U5097 ( .I1(n3482), .I2(\registres[19][24] ), .O(n4094) );
  NAND_GATE U5098 ( .I1(n3483), .I2(\registres[21][24] ), .O(n4093) );
  NAND_GATE U5099 ( .I1(n3484), .I2(\registres[6][24] ), .O(n4092) );
  NAND_GATE U5100 ( .I1(n3485), .I2(\registres[7][24] ), .O(n4090) );
  NAND_GATE U5101 ( .I1(n3486), .I2(\registres[30][24] ), .O(n4089) );
  NAND_GATE U5102 ( .I1(n3487), .I2(\registres[31][24] ), .O(n4088) );
  NAND_GATE U5103 ( .I1(n3488), .I2(\registres[14][24] ), .O(n4087) );
  AND4_GATE U5104 ( .I1(n4096), .I2(n4097), .I3(n4098), .I4(n4099), .O(n4065)
         );
  AND4_GATE U5105 ( .I1(n4100), .I2(n4101), .I3(n4102), .I4(n4103), .O(n4099)
         );
  NAND_GATE U5106 ( .I1(n3497), .I2(\registres[22][24] ), .O(n4103) );
  NAND_GATE U5107 ( .I1(n3498), .I2(\registres[15][24] ), .O(n4102) );
  NAND_GATE U5108 ( .I1(n3499), .I2(\registres[23][24] ), .O(n4101) );
  NAND_GATE U5109 ( .I1(n3500), .I2(\registres[4][24] ), .O(n4100) );
  NAND_GATE U5110 ( .I1(n3501), .I2(\registres[8][24] ), .O(n4098) );
  NAND_GATE U5111 ( .I1(n3502), .I2(\registres[2][24] ), .O(n4097) );
  NAND_GATE U5112 ( .I1(n3503), .I2(\registres[16][24] ), .O(n4096) );
  AND_GATE U5113 ( .I1(n4104), .I2(n3432), .O(data_src1[23]) );
  NAND4_GATE U5114 ( .I1(n4105), .I2(n4106), .I3(n4107), .I4(n4108), .O(n4104)
         );
  AND5_GATE U5115 ( .I1(n4109), .I2(n4110), .I3(n4111), .I4(n4112), .I5(n4113), 
        .O(n4108) );
  AND4_GATE U5116 ( .I1(n4114), .I2(n4115), .I3(n4116), .I4(n4117), .O(n4113)
         );
  NAND_GATE U5117 ( .I1(n3447), .I2(\registres[24][23] ), .O(n4117) );
  NAND_GATE U5118 ( .I1(n3448), .I2(\registres[25][23] ), .O(n4116) );
  NAND_GATE U5119 ( .I1(n3449), .I2(\registres[3][23] ), .O(n4115) );
  NAND_GATE U5120 ( .I1(n3450), .I2(\registres[26][23] ), .O(n4114) );
  NAND_GATE U5121 ( .I1(n3451), .I2(\registres[27][23] ), .O(n4112) );
  NAND_GATE U5122 ( .I1(n3452), .I2(\registres[10][23] ), .O(n4111) );
  NAND_GATE U5123 ( .I1(n3453), .I2(\registres[18][23] ), .O(n4110) );
  NAND_GATE U5124 ( .I1(n3454), .I2(\registres[5][23] ), .O(n4109) );
  AND5_GATE U5125 ( .I1(n4118), .I2(n4119), .I3(n4120), .I4(n4121), .I5(n4122), 
        .O(n4107) );
  AND4_GATE U5126 ( .I1(n4123), .I2(n4124), .I3(n4125), .I4(n4126), .O(n4122)
         );
  NAND_GATE U5127 ( .I1(n3464), .I2(\registres[28][23] ), .O(n4126) );
  NAND_GATE U5128 ( .I1(n3465), .I2(\registres[29][23] ), .O(n4125) );
  NAND_GATE U5129 ( .I1(n3466), .I2(\registres[12][23] ), .O(n4124) );
  NAND_GATE U5130 ( .I1(n3467), .I2(\registres[20][23] ), .O(n4123) );
  NAND_GATE U5131 ( .I1(n3468), .I2(\registres[1][23] ), .O(n4121) );
  NAND_GATE U5132 ( .I1(n3469), .I2(\registres[9][23] ), .O(n4120) );
  NAND_GATE U5133 ( .I1(n3470), .I2(\registres[11][23] ), .O(n4119) );
  NAND_GATE U5134 ( .I1(n3471), .I2(\registres[13][23] ), .O(n4118) );
  AND5_GATE U5135 ( .I1(n4127), .I2(n4128), .I3(n4129), .I4(n4130), .I5(n4131), 
        .O(n4106) );
  AND4_GATE U5136 ( .I1(n4132), .I2(n4133), .I3(n4134), .I4(n4135), .O(n4131)
         );
  NAND_GATE U5137 ( .I1(n3481), .I2(\registres[17][23] ), .O(n4135) );
  NAND_GATE U5138 ( .I1(n3482), .I2(\registres[19][23] ), .O(n4134) );
  NAND_GATE U5139 ( .I1(n3483), .I2(\registres[21][23] ), .O(n4133) );
  NAND_GATE U5140 ( .I1(n3484), .I2(\registres[6][23] ), .O(n4132) );
  NAND_GATE U5141 ( .I1(n3485), .I2(\registres[7][23] ), .O(n4130) );
  NAND_GATE U5142 ( .I1(n3486), .I2(\registres[30][23] ), .O(n4129) );
  NAND_GATE U5143 ( .I1(n3487), .I2(\registres[31][23] ), .O(n4128) );
  NAND_GATE U5144 ( .I1(n3488), .I2(\registres[14][23] ), .O(n4127) );
  AND4_GATE U5145 ( .I1(n4136), .I2(n4137), .I3(n4138), .I4(n4139), .O(n4105)
         );
  AND4_GATE U5146 ( .I1(n4140), .I2(n4141), .I3(n4142), .I4(n4143), .O(n4139)
         );
  NAND_GATE U5147 ( .I1(n3497), .I2(\registres[22][23] ), .O(n4143) );
  NAND_GATE U5148 ( .I1(n3498), .I2(\registres[15][23] ), .O(n4142) );
  NAND_GATE U5149 ( .I1(n3499), .I2(\registres[23][23] ), .O(n4141) );
  NAND_GATE U5150 ( .I1(n3500), .I2(\registres[4][23] ), .O(n4140) );
  NAND_GATE U5151 ( .I1(n3501), .I2(\registres[8][23] ), .O(n4138) );
  NAND_GATE U5152 ( .I1(n3502), .I2(\registres[2][23] ), .O(n4137) );
  NAND_GATE U5153 ( .I1(n3503), .I2(\registres[16][23] ), .O(n4136) );
  AND_GATE U5154 ( .I1(n4144), .I2(n3432), .O(data_src1[22]) );
  NAND4_GATE U5155 ( .I1(n4145), .I2(n4146), .I3(n4147), .I4(n4148), .O(n4144)
         );
  AND5_GATE U5156 ( .I1(n4149), .I2(n4150), .I3(n4151), .I4(n4152), .I5(n4153), 
        .O(n4148) );
  AND4_GATE U5157 ( .I1(n4154), .I2(n4155), .I3(n4156), .I4(n4157), .O(n4153)
         );
  NAND_GATE U5158 ( .I1(n3447), .I2(\registres[24][22] ), .O(n4157) );
  NAND_GATE U5159 ( .I1(n3448), .I2(\registres[25][22] ), .O(n4156) );
  NAND_GATE U5160 ( .I1(n3449), .I2(\registres[3][22] ), .O(n4155) );
  NAND_GATE U5161 ( .I1(n3450), .I2(\registres[26][22] ), .O(n4154) );
  NAND_GATE U5162 ( .I1(n3451), .I2(\registres[27][22] ), .O(n4152) );
  NAND_GATE U5163 ( .I1(n3452), .I2(\registres[10][22] ), .O(n4151) );
  NAND_GATE U5164 ( .I1(n3453), .I2(\registres[18][22] ), .O(n4150) );
  NAND_GATE U5165 ( .I1(n3454), .I2(\registres[5][22] ), .O(n4149) );
  AND5_GATE U5166 ( .I1(n4158), .I2(n4159), .I3(n4160), .I4(n4161), .I5(n4162), 
        .O(n4147) );
  AND4_GATE U5167 ( .I1(n4163), .I2(n4164), .I3(n4165), .I4(n4166), .O(n4162)
         );
  NAND_GATE U5168 ( .I1(n3464), .I2(\registres[28][22] ), .O(n4166) );
  NAND_GATE U5169 ( .I1(n3465), .I2(\registres[29][22] ), .O(n4165) );
  NAND_GATE U5170 ( .I1(n3466), .I2(\registres[12][22] ), .O(n4164) );
  NAND_GATE U5171 ( .I1(n3467), .I2(\registres[20][22] ), .O(n4163) );
  NAND_GATE U5172 ( .I1(n3468), .I2(\registres[1][22] ), .O(n4161) );
  NAND_GATE U5173 ( .I1(n3469), .I2(\registres[9][22] ), .O(n4160) );
  NAND_GATE U5174 ( .I1(n3470), .I2(\registres[11][22] ), .O(n4159) );
  NAND_GATE U5175 ( .I1(n3471), .I2(\registres[13][22] ), .O(n4158) );
  AND5_GATE U5176 ( .I1(n4167), .I2(n4168), .I3(n4169), .I4(n4170), .I5(n4171), 
        .O(n4146) );
  AND4_GATE U5177 ( .I1(n4172), .I2(n4173), .I3(n4174), .I4(n4175), .O(n4171)
         );
  NAND_GATE U5178 ( .I1(n3481), .I2(\registres[17][22] ), .O(n4175) );
  NAND_GATE U5179 ( .I1(n3482), .I2(\registres[19][22] ), .O(n4174) );
  NAND_GATE U5180 ( .I1(n3483), .I2(\registres[21][22] ), .O(n4173) );
  NAND_GATE U5181 ( .I1(n3484), .I2(\registres[6][22] ), .O(n4172) );
  NAND_GATE U5182 ( .I1(n3485), .I2(\registres[7][22] ), .O(n4170) );
  NAND_GATE U5183 ( .I1(n3486), .I2(\registres[30][22] ), .O(n4169) );
  NAND_GATE U5184 ( .I1(n3487), .I2(\registres[31][22] ), .O(n4168) );
  NAND_GATE U5185 ( .I1(n3488), .I2(\registres[14][22] ), .O(n4167) );
  AND4_GATE U5186 ( .I1(n4176), .I2(n4177), .I3(n4178), .I4(n4179), .O(n4145)
         );
  AND4_GATE U5187 ( .I1(n4180), .I2(n4181), .I3(n4182), .I4(n4183), .O(n4179)
         );
  NAND_GATE U5188 ( .I1(n3497), .I2(\registres[22][22] ), .O(n4183) );
  NAND_GATE U5189 ( .I1(n3498), .I2(\registres[15][22] ), .O(n4182) );
  NAND_GATE U5190 ( .I1(n3499), .I2(\registres[23][22] ), .O(n4181) );
  NAND_GATE U5191 ( .I1(n3500), .I2(\registres[4][22] ), .O(n4180) );
  NAND_GATE U5192 ( .I1(n3501), .I2(\registres[8][22] ), .O(n4178) );
  NAND_GATE U5193 ( .I1(n3502), .I2(\registres[2][22] ), .O(n4177) );
  NAND_GATE U5194 ( .I1(n3503), .I2(\registres[16][22] ), .O(n4176) );
  AND_GATE U5195 ( .I1(n4184), .I2(n3432), .O(data_src1[21]) );
  NAND4_GATE U5196 ( .I1(n4185), .I2(n4186), .I3(n4187), .I4(n4188), .O(n4184)
         );
  AND5_GATE U5197 ( .I1(n4189), .I2(n4190), .I3(n4191), .I4(n4192), .I5(n4193), 
        .O(n4188) );
  AND4_GATE U5198 ( .I1(n4194), .I2(n4195), .I3(n4196), .I4(n4197), .O(n4193)
         );
  NAND_GATE U5199 ( .I1(n3447), .I2(\registres[24][21] ), .O(n4197) );
  NAND_GATE U5200 ( .I1(n3448), .I2(\registres[25][21] ), .O(n4196) );
  NAND_GATE U5201 ( .I1(n3449), .I2(\registres[3][21] ), .O(n4195) );
  NAND_GATE U5202 ( .I1(n3450), .I2(\registres[26][21] ), .O(n4194) );
  NAND_GATE U5203 ( .I1(n3451), .I2(\registres[27][21] ), .O(n4192) );
  NAND_GATE U5204 ( .I1(n3452), .I2(\registres[10][21] ), .O(n4191) );
  NAND_GATE U5205 ( .I1(n3453), .I2(\registres[18][21] ), .O(n4190) );
  NAND_GATE U5206 ( .I1(n3454), .I2(\registres[5][21] ), .O(n4189) );
  AND5_GATE U5207 ( .I1(n4198), .I2(n4199), .I3(n4200), .I4(n4201), .I5(n4202), 
        .O(n4187) );
  AND4_GATE U5208 ( .I1(n4203), .I2(n4204), .I3(n4205), .I4(n4206), .O(n4202)
         );
  NAND_GATE U5209 ( .I1(n3464), .I2(\registres[28][21] ), .O(n4206) );
  NAND_GATE U5210 ( .I1(n3465), .I2(\registres[29][21] ), .O(n4205) );
  NAND_GATE U5211 ( .I1(n3466), .I2(\registres[12][21] ), .O(n4204) );
  NAND_GATE U5212 ( .I1(n3467), .I2(\registres[20][21] ), .O(n4203) );
  NAND_GATE U5213 ( .I1(n3468), .I2(\registres[1][21] ), .O(n4201) );
  NAND_GATE U5214 ( .I1(n3469), .I2(\registres[9][21] ), .O(n4200) );
  NAND_GATE U5215 ( .I1(n3470), .I2(\registres[11][21] ), .O(n4199) );
  NAND_GATE U5216 ( .I1(n3471), .I2(\registres[13][21] ), .O(n4198) );
  AND5_GATE U5217 ( .I1(n4207), .I2(n4208), .I3(n4209), .I4(n4210), .I5(n4211), 
        .O(n4186) );
  AND4_GATE U5218 ( .I1(n4212), .I2(n4213), .I3(n4214), .I4(n4215), .O(n4211)
         );
  NAND_GATE U5219 ( .I1(n3481), .I2(\registres[17][21] ), .O(n4215) );
  NAND_GATE U5220 ( .I1(n3482), .I2(\registres[19][21] ), .O(n4214) );
  NAND_GATE U5221 ( .I1(n3483), .I2(\registres[21][21] ), .O(n4213) );
  NAND_GATE U5222 ( .I1(n3484), .I2(\registres[6][21] ), .O(n4212) );
  NAND_GATE U5223 ( .I1(n3485), .I2(\registres[7][21] ), .O(n4210) );
  NAND_GATE U5224 ( .I1(n3486), .I2(\registres[30][21] ), .O(n4209) );
  NAND_GATE U5225 ( .I1(n3487), .I2(\registres[31][21] ), .O(n4208) );
  NAND_GATE U5226 ( .I1(n3488), .I2(\registres[14][21] ), .O(n4207) );
  AND4_GATE U5227 ( .I1(n4216), .I2(n4217), .I3(n4218), .I4(n4219), .O(n4185)
         );
  AND4_GATE U5228 ( .I1(n4220), .I2(n4221), .I3(n4222), .I4(n4223), .O(n4219)
         );
  NAND_GATE U5229 ( .I1(n3497), .I2(\registres[22][21] ), .O(n4223) );
  NAND_GATE U5230 ( .I1(n3498), .I2(\registres[15][21] ), .O(n4222) );
  NAND_GATE U5231 ( .I1(n3499), .I2(\registres[23][21] ), .O(n4221) );
  NAND_GATE U5232 ( .I1(n3500), .I2(\registres[4][21] ), .O(n4220) );
  NAND_GATE U5233 ( .I1(n3501), .I2(\registres[8][21] ), .O(n4218) );
  NAND_GATE U5234 ( .I1(n3502), .I2(\registres[2][21] ), .O(n4217) );
  NAND_GATE U5235 ( .I1(n3503), .I2(\registres[16][21] ), .O(n4216) );
  AND_GATE U5236 ( .I1(n4224), .I2(n3432), .O(data_src1[20]) );
  NAND4_GATE U5237 ( .I1(n4225), .I2(n4226), .I3(n4227), .I4(n4228), .O(n4224)
         );
  AND5_GATE U5238 ( .I1(n4229), .I2(n4230), .I3(n4231), .I4(n4232), .I5(n4233), 
        .O(n4228) );
  AND4_GATE U5239 ( .I1(n4234), .I2(n4235), .I3(n4236), .I4(n4237), .O(n4233)
         );
  NAND_GATE U5240 ( .I1(n3447), .I2(\registres[24][20] ), .O(n4237) );
  NAND_GATE U5241 ( .I1(n3448), .I2(\registres[25][20] ), .O(n4236) );
  NAND_GATE U5242 ( .I1(n3449), .I2(\registres[3][20] ), .O(n4235) );
  NAND_GATE U5243 ( .I1(n3450), .I2(\registres[26][20] ), .O(n4234) );
  NAND_GATE U5244 ( .I1(n3451), .I2(\registres[27][20] ), .O(n4232) );
  NAND_GATE U5245 ( .I1(n3452), .I2(\registres[10][20] ), .O(n4231) );
  NAND_GATE U5246 ( .I1(n3453), .I2(\registres[18][20] ), .O(n4230) );
  NAND_GATE U5247 ( .I1(n3454), .I2(\registres[5][20] ), .O(n4229) );
  AND5_GATE U5248 ( .I1(n4238), .I2(n4239), .I3(n4240), .I4(n4241), .I5(n4242), 
        .O(n4227) );
  AND4_GATE U5249 ( .I1(n4243), .I2(n4244), .I3(n4245), .I4(n4246), .O(n4242)
         );
  NAND_GATE U5250 ( .I1(n3464), .I2(\registres[28][20] ), .O(n4246) );
  NAND_GATE U5251 ( .I1(n3465), .I2(\registres[29][20] ), .O(n4245) );
  NAND_GATE U5252 ( .I1(n3466), .I2(\registres[12][20] ), .O(n4244) );
  NAND_GATE U5253 ( .I1(n3467), .I2(\registres[20][20] ), .O(n4243) );
  NAND_GATE U5254 ( .I1(n3468), .I2(\registres[1][20] ), .O(n4241) );
  NAND_GATE U5255 ( .I1(n3469), .I2(\registres[9][20] ), .O(n4240) );
  NAND_GATE U5256 ( .I1(n3470), .I2(\registres[11][20] ), .O(n4239) );
  NAND_GATE U5257 ( .I1(n3471), .I2(\registres[13][20] ), .O(n4238) );
  AND5_GATE U5258 ( .I1(n4247), .I2(n4248), .I3(n4249), .I4(n4250), .I5(n4251), 
        .O(n4226) );
  AND4_GATE U5259 ( .I1(n4252), .I2(n4253), .I3(n4254), .I4(n4255), .O(n4251)
         );
  NAND_GATE U5260 ( .I1(n3481), .I2(\registres[17][20] ), .O(n4255) );
  NAND_GATE U5261 ( .I1(n3482), .I2(\registres[19][20] ), .O(n4254) );
  NAND_GATE U5262 ( .I1(n3483), .I2(\registres[21][20] ), .O(n4253) );
  NAND_GATE U5263 ( .I1(n3484), .I2(\registres[6][20] ), .O(n4252) );
  NAND_GATE U5264 ( .I1(n3485), .I2(\registres[7][20] ), .O(n4250) );
  NAND_GATE U5265 ( .I1(n3486), .I2(\registres[30][20] ), .O(n4249) );
  NAND_GATE U5266 ( .I1(n3487), .I2(\registres[31][20] ), .O(n4248) );
  NAND_GATE U5267 ( .I1(n3488), .I2(\registres[14][20] ), .O(n4247) );
  AND4_GATE U5268 ( .I1(n4256), .I2(n4257), .I3(n4258), .I4(n4259), .O(n4225)
         );
  AND4_GATE U5269 ( .I1(n4260), .I2(n4261), .I3(n4262), .I4(n4263), .O(n4259)
         );
  NAND_GATE U5270 ( .I1(n3497), .I2(\registres[22][20] ), .O(n4263) );
  NAND_GATE U5271 ( .I1(n3498), .I2(\registres[15][20] ), .O(n4262) );
  NAND_GATE U5272 ( .I1(n3499), .I2(\registres[23][20] ), .O(n4261) );
  NAND_GATE U5273 ( .I1(n3500), .I2(\registres[4][20] ), .O(n4260) );
  NAND_GATE U5274 ( .I1(n3501), .I2(\registres[8][20] ), .O(n4258) );
  NAND_GATE U5275 ( .I1(n3502), .I2(\registres[2][20] ), .O(n4257) );
  NAND_GATE U5276 ( .I1(n3503), .I2(\registres[16][20] ), .O(n4256) );
  AND_GATE U5277 ( .I1(n4264), .I2(n3432), .O(data_src1[1]) );
  NAND4_GATE U5278 ( .I1(n4265), .I2(n4266), .I3(n4267), .I4(n4268), .O(n4264)
         );
  AND5_GATE U5279 ( .I1(n4269), .I2(n4270), .I3(n4271), .I4(n4272), .I5(n4273), 
        .O(n4268) );
  AND4_GATE U5280 ( .I1(n4274), .I2(n4275), .I3(n4276), .I4(n4277), .O(n4273)
         );
  NAND_GATE U5281 ( .I1(n3447), .I2(\registres[24][1] ), .O(n4277) );
  NAND_GATE U5282 ( .I1(n3448), .I2(\registres[25][1] ), .O(n4276) );
  NAND_GATE U5283 ( .I1(n3449), .I2(\registres[3][1] ), .O(n4275) );
  NAND_GATE U5284 ( .I1(n3450), .I2(\registres[26][1] ), .O(n4274) );
  NAND_GATE U5285 ( .I1(n3451), .I2(\registres[27][1] ), .O(n4272) );
  NAND_GATE U5286 ( .I1(n3452), .I2(\registres[10][1] ), .O(n4271) );
  NAND_GATE U5287 ( .I1(n3453), .I2(\registres[18][1] ), .O(n4270) );
  NAND_GATE U5288 ( .I1(n3454), .I2(\registres[5][1] ), .O(n4269) );
  AND5_GATE U5289 ( .I1(n4278), .I2(n4279), .I3(n4280), .I4(n4281), .I5(n4282), 
        .O(n4267) );
  AND4_GATE U5290 ( .I1(n4283), .I2(n4284), .I3(n4285), .I4(n4286), .O(n4282)
         );
  NAND_GATE U5291 ( .I1(n3464), .I2(\registres[28][1] ), .O(n4286) );
  NAND_GATE U5292 ( .I1(n3465), .I2(\registres[29][1] ), .O(n4285) );
  NAND_GATE U5293 ( .I1(n3466), .I2(\registres[12][1] ), .O(n4284) );
  NAND_GATE U5294 ( .I1(n3467), .I2(\registres[20][1] ), .O(n4283) );
  NAND_GATE U5295 ( .I1(n3468), .I2(\registres[1][1] ), .O(n4281) );
  NAND_GATE U5296 ( .I1(n3469), .I2(\registres[9][1] ), .O(n4280) );
  NAND_GATE U5297 ( .I1(n3470), .I2(\registres[11][1] ), .O(n4279) );
  NAND_GATE U5298 ( .I1(n3471), .I2(\registres[13][1] ), .O(n4278) );
  AND5_GATE U5299 ( .I1(n4287), .I2(n4288), .I3(n4289), .I4(n4290), .I5(n4291), 
        .O(n4266) );
  AND4_GATE U5300 ( .I1(n4292), .I2(n4293), .I3(n4294), .I4(n4295), .O(n4291)
         );
  NAND_GATE U5301 ( .I1(n3481), .I2(\registres[17][1] ), .O(n4295) );
  NAND_GATE U5302 ( .I1(n3482), .I2(\registres[19][1] ), .O(n4294) );
  NAND_GATE U5303 ( .I1(n3483), .I2(\registres[21][1] ), .O(n4293) );
  NAND_GATE U5304 ( .I1(n3484), .I2(\registres[6][1] ), .O(n4292) );
  NAND_GATE U5305 ( .I1(n3485), .I2(\registres[7][1] ), .O(n4290) );
  NAND_GATE U5306 ( .I1(n3486), .I2(\registres[30][1] ), .O(n4289) );
  NAND_GATE U5307 ( .I1(n3487), .I2(\registres[31][1] ), .O(n4288) );
  NAND_GATE U5308 ( .I1(n3488), .I2(\registres[14][1] ), .O(n4287) );
  AND4_GATE U5309 ( .I1(n4296), .I2(n4297), .I3(n4298), .I4(n4299), .O(n4265)
         );
  AND4_GATE U5310 ( .I1(n4300), .I2(n4301), .I3(n4302), .I4(n4303), .O(n4299)
         );
  NAND_GATE U5311 ( .I1(n3497), .I2(\registres[22][1] ), .O(n4303) );
  NAND_GATE U5312 ( .I1(n3498), .I2(\registres[15][1] ), .O(n4302) );
  NAND_GATE U5313 ( .I1(n3499), .I2(\registres[23][1] ), .O(n4301) );
  NAND_GATE U5314 ( .I1(n3500), .I2(\registres[4][1] ), .O(n4300) );
  NAND_GATE U5315 ( .I1(n3501), .I2(\registres[8][1] ), .O(n4298) );
  NAND_GATE U5316 ( .I1(n3502), .I2(\registres[2][1] ), .O(n4297) );
  NAND_GATE U5317 ( .I1(n3503), .I2(\registres[16][1] ), .O(n4296) );
  AND_GATE U5318 ( .I1(n4304), .I2(n3432), .O(data_src1[19]) );
  NAND4_GATE U5319 ( .I1(n4305), .I2(n4306), .I3(n4307), .I4(n4308), .O(n4304)
         );
  AND5_GATE U5320 ( .I1(n4309), .I2(n4310), .I3(n4311), .I4(n4312), .I5(n4313), 
        .O(n4308) );
  AND4_GATE U5321 ( .I1(n4314), .I2(n4315), .I3(n4316), .I4(n4317), .O(n4313)
         );
  NAND_GATE U5322 ( .I1(n3447), .I2(\registres[24][19] ), .O(n4317) );
  NAND_GATE U5323 ( .I1(n3448), .I2(\registres[25][19] ), .O(n4316) );
  NAND_GATE U5324 ( .I1(n3449), .I2(\registres[3][19] ), .O(n4315) );
  NAND_GATE U5325 ( .I1(n3450), .I2(\registres[26][19] ), .O(n4314) );
  NAND_GATE U5326 ( .I1(n3451), .I2(\registres[27][19] ), .O(n4312) );
  NAND_GATE U5327 ( .I1(n3452), .I2(\registres[10][19] ), .O(n4311) );
  NAND_GATE U5328 ( .I1(n3453), .I2(\registres[18][19] ), .O(n4310) );
  NAND_GATE U5329 ( .I1(n3454), .I2(\registres[5][19] ), .O(n4309) );
  AND5_GATE U5330 ( .I1(n4318), .I2(n4319), .I3(n4320), .I4(n4321), .I5(n4322), 
        .O(n4307) );
  AND4_GATE U5331 ( .I1(n4323), .I2(n4324), .I3(n4325), .I4(n4326), .O(n4322)
         );
  NAND_GATE U5332 ( .I1(n3464), .I2(\registres[28][19] ), .O(n4326) );
  NAND_GATE U5333 ( .I1(n3465), .I2(\registres[29][19] ), .O(n4325) );
  NAND_GATE U5334 ( .I1(n3466), .I2(\registres[12][19] ), .O(n4324) );
  NAND_GATE U5335 ( .I1(n3467), .I2(\registres[20][19] ), .O(n4323) );
  NAND_GATE U5336 ( .I1(n3468), .I2(\registres[1][19] ), .O(n4321) );
  NAND_GATE U5337 ( .I1(n3469), .I2(\registres[9][19] ), .O(n4320) );
  NAND_GATE U5338 ( .I1(n3470), .I2(\registres[11][19] ), .O(n4319) );
  NAND_GATE U5339 ( .I1(n3471), .I2(\registres[13][19] ), .O(n4318) );
  AND5_GATE U5340 ( .I1(n4327), .I2(n4328), .I3(n4329), .I4(n4330), .I5(n4331), 
        .O(n4306) );
  AND4_GATE U5341 ( .I1(n4332), .I2(n4333), .I3(n4334), .I4(n4335), .O(n4331)
         );
  NAND_GATE U5342 ( .I1(n3481), .I2(\registres[17][19] ), .O(n4335) );
  NAND_GATE U5343 ( .I1(n3482), .I2(\registres[19][19] ), .O(n4334) );
  NAND_GATE U5344 ( .I1(n3483), .I2(\registres[21][19] ), .O(n4333) );
  NAND_GATE U5345 ( .I1(n3484), .I2(\registres[6][19] ), .O(n4332) );
  NAND_GATE U5346 ( .I1(n3485), .I2(\registres[7][19] ), .O(n4330) );
  NAND_GATE U5347 ( .I1(n3486), .I2(\registres[30][19] ), .O(n4329) );
  NAND_GATE U5348 ( .I1(n3487), .I2(\registres[31][19] ), .O(n4328) );
  NAND_GATE U5349 ( .I1(n3488), .I2(\registres[14][19] ), .O(n4327) );
  AND4_GATE U5350 ( .I1(n4336), .I2(n4337), .I3(n4338), .I4(n4339), .O(n4305)
         );
  AND4_GATE U5351 ( .I1(n4340), .I2(n4341), .I3(n4342), .I4(n4343), .O(n4339)
         );
  NAND_GATE U5352 ( .I1(n3497), .I2(\registres[22][19] ), .O(n4343) );
  NAND_GATE U5353 ( .I1(n3498), .I2(\registres[15][19] ), .O(n4342) );
  NAND_GATE U5354 ( .I1(n3499), .I2(\registres[23][19] ), .O(n4341) );
  NAND_GATE U5355 ( .I1(n3500), .I2(\registres[4][19] ), .O(n4340) );
  NAND_GATE U5356 ( .I1(n3501), .I2(\registres[8][19] ), .O(n4338) );
  NAND_GATE U5357 ( .I1(n3502), .I2(\registres[2][19] ), .O(n4337) );
  NAND_GATE U5358 ( .I1(n3503), .I2(\registres[16][19] ), .O(n4336) );
  AND_GATE U5359 ( .I1(n4344), .I2(n3432), .O(data_src1[18]) );
  NAND4_GATE U5360 ( .I1(n4345), .I2(n4346), .I3(n4347), .I4(n4348), .O(n4344)
         );
  AND5_GATE U5361 ( .I1(n4349), .I2(n4350), .I3(n4351), .I4(n4352), .I5(n4353), 
        .O(n4348) );
  AND4_GATE U5362 ( .I1(n4354), .I2(n4355), .I3(n4356), .I4(n4357), .O(n4353)
         );
  NAND_GATE U5363 ( .I1(n3447), .I2(\registres[24][18] ), .O(n4357) );
  NAND_GATE U5364 ( .I1(n3448), .I2(\registres[25][18] ), .O(n4356) );
  NAND_GATE U5365 ( .I1(n3449), .I2(\registres[3][18] ), .O(n4355) );
  NAND_GATE U5366 ( .I1(n3450), .I2(\registres[26][18] ), .O(n4354) );
  NAND_GATE U5367 ( .I1(n3451), .I2(\registres[27][18] ), .O(n4352) );
  NAND_GATE U5368 ( .I1(n3452), .I2(\registres[10][18] ), .O(n4351) );
  NAND_GATE U5369 ( .I1(n3453), .I2(\registres[18][18] ), .O(n4350) );
  NAND_GATE U5370 ( .I1(n3454), .I2(\registres[5][18] ), .O(n4349) );
  AND5_GATE U5371 ( .I1(n4358), .I2(n4359), .I3(n4360), .I4(n4361), .I5(n4362), 
        .O(n4347) );
  AND4_GATE U5372 ( .I1(n4363), .I2(n4364), .I3(n4365), .I4(n4366), .O(n4362)
         );
  NAND_GATE U5373 ( .I1(n3464), .I2(\registres[28][18] ), .O(n4366) );
  NAND_GATE U5374 ( .I1(n3465), .I2(\registres[29][18] ), .O(n4365) );
  NAND_GATE U5375 ( .I1(n3466), .I2(\registres[12][18] ), .O(n4364) );
  NAND_GATE U5376 ( .I1(n3467), .I2(\registres[20][18] ), .O(n4363) );
  NAND_GATE U5377 ( .I1(n3468), .I2(\registres[1][18] ), .O(n4361) );
  NAND_GATE U5378 ( .I1(n3469), .I2(\registres[9][18] ), .O(n4360) );
  NAND_GATE U5379 ( .I1(n3470), .I2(\registres[11][18] ), .O(n4359) );
  NAND_GATE U5380 ( .I1(n3471), .I2(\registres[13][18] ), .O(n4358) );
  AND5_GATE U5381 ( .I1(n4367), .I2(n4368), .I3(n4369), .I4(n4370), .I5(n4371), 
        .O(n4346) );
  AND4_GATE U5382 ( .I1(n4372), .I2(n4373), .I3(n4374), .I4(n4375), .O(n4371)
         );
  NAND_GATE U5383 ( .I1(n3481), .I2(\registres[17][18] ), .O(n4375) );
  NAND_GATE U5384 ( .I1(n3482), .I2(\registres[19][18] ), .O(n4374) );
  NAND_GATE U5385 ( .I1(n3483), .I2(\registres[21][18] ), .O(n4373) );
  NAND_GATE U5386 ( .I1(n3484), .I2(\registres[6][18] ), .O(n4372) );
  NAND_GATE U5387 ( .I1(n3485), .I2(\registres[7][18] ), .O(n4370) );
  NAND_GATE U5388 ( .I1(n3486), .I2(\registres[30][18] ), .O(n4369) );
  NAND_GATE U5389 ( .I1(n3487), .I2(\registres[31][18] ), .O(n4368) );
  NAND_GATE U5390 ( .I1(n3488), .I2(\registres[14][18] ), .O(n4367) );
  AND4_GATE U5391 ( .I1(n4376), .I2(n4377), .I3(n4378), .I4(n4379), .O(n4345)
         );
  AND4_GATE U5392 ( .I1(n4380), .I2(n4381), .I3(n4382), .I4(n4383), .O(n4379)
         );
  NAND_GATE U5393 ( .I1(n3497), .I2(\registres[22][18] ), .O(n4383) );
  NAND_GATE U5394 ( .I1(n3498), .I2(\registres[15][18] ), .O(n4382) );
  NAND_GATE U5395 ( .I1(n3499), .I2(\registres[23][18] ), .O(n4381) );
  NAND_GATE U5396 ( .I1(n3500), .I2(\registres[4][18] ), .O(n4380) );
  NAND_GATE U5397 ( .I1(n3501), .I2(\registres[8][18] ), .O(n4378) );
  NAND_GATE U5398 ( .I1(n3502), .I2(\registres[2][18] ), .O(n4377) );
  NAND_GATE U5399 ( .I1(n3503), .I2(\registres[16][18] ), .O(n4376) );
  AND_GATE U5400 ( .I1(n4384), .I2(n3432), .O(data_src1[17]) );
  NAND4_GATE U5401 ( .I1(n4385), .I2(n4386), .I3(n4387), .I4(n4388), .O(n4384)
         );
  AND5_GATE U5402 ( .I1(n4389), .I2(n4390), .I3(n4391), .I4(n4392), .I5(n4393), 
        .O(n4388) );
  AND4_GATE U5403 ( .I1(n4394), .I2(n4395), .I3(n4396), .I4(n4397), .O(n4393)
         );
  NAND_GATE U5404 ( .I1(n3447), .I2(\registres[24][17] ), .O(n4397) );
  NAND_GATE U5405 ( .I1(n3448), .I2(\registres[25][17] ), .O(n4396) );
  NAND_GATE U5406 ( .I1(n3449), .I2(\registres[3][17] ), .O(n4395) );
  NAND_GATE U5407 ( .I1(n3450), .I2(\registres[26][17] ), .O(n4394) );
  NAND_GATE U5408 ( .I1(n3451), .I2(\registres[27][17] ), .O(n4392) );
  NAND_GATE U5409 ( .I1(n3452), .I2(\registres[10][17] ), .O(n4391) );
  NAND_GATE U5410 ( .I1(n3453), .I2(\registres[18][17] ), .O(n4390) );
  NAND_GATE U5411 ( .I1(n3454), .I2(\registres[5][17] ), .O(n4389) );
  AND5_GATE U5412 ( .I1(n4398), .I2(n4399), .I3(n4400), .I4(n4401), .I5(n4402), 
        .O(n4387) );
  AND4_GATE U5413 ( .I1(n4403), .I2(n4404), .I3(n4405), .I4(n4406), .O(n4402)
         );
  NAND_GATE U5414 ( .I1(n3464), .I2(\registres[28][17] ), .O(n4406) );
  NAND_GATE U5415 ( .I1(n3465), .I2(\registres[29][17] ), .O(n4405) );
  NAND_GATE U5416 ( .I1(n3466), .I2(\registres[12][17] ), .O(n4404) );
  NAND_GATE U5417 ( .I1(n3467), .I2(\registres[20][17] ), .O(n4403) );
  NAND_GATE U5418 ( .I1(n3468), .I2(\registres[1][17] ), .O(n4401) );
  NAND_GATE U5419 ( .I1(n3469), .I2(\registres[9][17] ), .O(n4400) );
  NAND_GATE U5420 ( .I1(n3470), .I2(\registres[11][17] ), .O(n4399) );
  NAND_GATE U5421 ( .I1(n3471), .I2(\registres[13][17] ), .O(n4398) );
  AND5_GATE U5422 ( .I1(n4407), .I2(n4408), .I3(n4409), .I4(n4410), .I5(n4411), 
        .O(n4386) );
  AND4_GATE U5423 ( .I1(n4412), .I2(n4413), .I3(n4414), .I4(n4415), .O(n4411)
         );
  NAND_GATE U5424 ( .I1(n3481), .I2(\registres[17][17] ), .O(n4415) );
  NAND_GATE U5425 ( .I1(n3482), .I2(\registres[19][17] ), .O(n4414) );
  NAND_GATE U5426 ( .I1(n3483), .I2(\registres[21][17] ), .O(n4413) );
  NAND_GATE U5427 ( .I1(n3484), .I2(\registres[6][17] ), .O(n4412) );
  NAND_GATE U5428 ( .I1(n3485), .I2(\registres[7][17] ), .O(n4410) );
  NAND_GATE U5429 ( .I1(n3486), .I2(\registres[30][17] ), .O(n4409) );
  NAND_GATE U5430 ( .I1(n3487), .I2(\registres[31][17] ), .O(n4408) );
  NAND_GATE U5431 ( .I1(n3488), .I2(\registres[14][17] ), .O(n4407) );
  AND4_GATE U5432 ( .I1(n4416), .I2(n4417), .I3(n4418), .I4(n4419), .O(n4385)
         );
  AND4_GATE U5433 ( .I1(n4420), .I2(n4421), .I3(n4422), .I4(n4423), .O(n4419)
         );
  NAND_GATE U5434 ( .I1(n3497), .I2(\registres[22][17] ), .O(n4423) );
  NAND_GATE U5435 ( .I1(n3498), .I2(\registres[15][17] ), .O(n4422) );
  NAND_GATE U5436 ( .I1(n3499), .I2(\registres[23][17] ), .O(n4421) );
  NAND_GATE U5437 ( .I1(n3500), .I2(\registres[4][17] ), .O(n4420) );
  NAND_GATE U5438 ( .I1(n3501), .I2(\registres[8][17] ), .O(n4418) );
  NAND_GATE U5439 ( .I1(n3502), .I2(\registres[2][17] ), .O(n4417) );
  NAND_GATE U5440 ( .I1(n3503), .I2(\registres[16][17] ), .O(n4416) );
  AND_GATE U5441 ( .I1(n4424), .I2(n3432), .O(data_src1[16]) );
  NAND4_GATE U5442 ( .I1(n4425), .I2(n4426), .I3(n4427), .I4(n4428), .O(n4424)
         );
  AND5_GATE U5443 ( .I1(n4429), .I2(n4430), .I3(n4431), .I4(n4432), .I5(n4433), 
        .O(n4428) );
  AND4_GATE U5444 ( .I1(n4434), .I2(n4435), .I3(n4436), .I4(n4437), .O(n4433)
         );
  NAND_GATE U5445 ( .I1(n3447), .I2(\registres[24][16] ), .O(n4437) );
  NAND_GATE U5446 ( .I1(n3448), .I2(\registres[25][16] ), .O(n4436) );
  NAND_GATE U5447 ( .I1(n3449), .I2(\registres[3][16] ), .O(n4435) );
  NAND_GATE U5448 ( .I1(n3450), .I2(\registres[26][16] ), .O(n4434) );
  NAND_GATE U5449 ( .I1(n3451), .I2(\registres[27][16] ), .O(n4432) );
  NAND_GATE U5450 ( .I1(n3452), .I2(\registres[10][16] ), .O(n4431) );
  NAND_GATE U5451 ( .I1(n3453), .I2(\registres[18][16] ), .O(n4430) );
  NAND_GATE U5452 ( .I1(n3454), .I2(\registres[5][16] ), .O(n4429) );
  AND5_GATE U5453 ( .I1(n4438), .I2(n4439), .I3(n4440), .I4(n4441), .I5(n4442), 
        .O(n4427) );
  AND4_GATE U5454 ( .I1(n4443), .I2(n4444), .I3(n4445), .I4(n4446), .O(n4442)
         );
  NAND_GATE U5455 ( .I1(n3464), .I2(\registres[28][16] ), .O(n4446) );
  NAND_GATE U5456 ( .I1(n3465), .I2(\registres[29][16] ), .O(n4445) );
  NAND_GATE U5457 ( .I1(n3466), .I2(\registres[12][16] ), .O(n4444) );
  NAND_GATE U5458 ( .I1(n3467), .I2(\registres[20][16] ), .O(n4443) );
  NAND_GATE U5459 ( .I1(n3468), .I2(\registres[1][16] ), .O(n4441) );
  NAND_GATE U5460 ( .I1(n3469), .I2(\registres[9][16] ), .O(n4440) );
  NAND_GATE U5461 ( .I1(n3470), .I2(\registres[11][16] ), .O(n4439) );
  NAND_GATE U5462 ( .I1(n3471), .I2(\registres[13][16] ), .O(n4438) );
  AND5_GATE U5463 ( .I1(n4447), .I2(n4448), .I3(n4449), .I4(n4450), .I5(n4451), 
        .O(n4426) );
  AND4_GATE U5464 ( .I1(n4452), .I2(n4453), .I3(n4454), .I4(n4455), .O(n4451)
         );
  NAND_GATE U5465 ( .I1(n3481), .I2(\registres[17][16] ), .O(n4455) );
  NAND_GATE U5466 ( .I1(n3482), .I2(\registres[19][16] ), .O(n4454) );
  NAND_GATE U5467 ( .I1(n3483), .I2(\registres[21][16] ), .O(n4453) );
  NAND_GATE U5468 ( .I1(n3484), .I2(\registres[6][16] ), .O(n4452) );
  NAND_GATE U5469 ( .I1(n3485), .I2(\registres[7][16] ), .O(n4450) );
  NAND_GATE U5470 ( .I1(n3486), .I2(\registres[30][16] ), .O(n4449) );
  NAND_GATE U5471 ( .I1(n3487), .I2(\registres[31][16] ), .O(n4448) );
  NAND_GATE U5472 ( .I1(n3488), .I2(\registres[14][16] ), .O(n4447) );
  AND4_GATE U5473 ( .I1(n4456), .I2(n4457), .I3(n4458), .I4(n4459), .O(n4425)
         );
  AND4_GATE U5474 ( .I1(n4460), .I2(n4461), .I3(n4462), .I4(n4463), .O(n4459)
         );
  NAND_GATE U5475 ( .I1(n3497), .I2(\registres[22][16] ), .O(n4463) );
  NAND_GATE U5476 ( .I1(n3498), .I2(\registres[15][16] ), .O(n4462) );
  NAND_GATE U5477 ( .I1(n3499), .I2(\registres[23][16] ), .O(n4461) );
  NAND_GATE U5478 ( .I1(n3500), .I2(\registres[4][16] ), .O(n4460) );
  NAND_GATE U5479 ( .I1(n3501), .I2(\registres[8][16] ), .O(n4458) );
  NAND_GATE U5480 ( .I1(n3502), .I2(\registres[2][16] ), .O(n4457) );
  NAND_GATE U5481 ( .I1(n3503), .I2(\registres[16][16] ), .O(n4456) );
  AND_GATE U5482 ( .I1(n4464), .I2(n3432), .O(data_src1[15]) );
  NAND4_GATE U5483 ( .I1(n4465), .I2(n4466), .I3(n4467), .I4(n4468), .O(n4464)
         );
  AND5_GATE U5484 ( .I1(n4469), .I2(n4470), .I3(n4471), .I4(n4472), .I5(n4473), 
        .O(n4468) );
  AND4_GATE U5485 ( .I1(n4474), .I2(n4475), .I3(n4476), .I4(n4477), .O(n4473)
         );
  NAND_GATE U5486 ( .I1(n3447), .I2(\registres[24][15] ), .O(n4477) );
  NAND_GATE U5487 ( .I1(n3448), .I2(\registres[25][15] ), .O(n4476) );
  NAND_GATE U5488 ( .I1(n3449), .I2(\registres[3][15] ), .O(n4475) );
  NAND_GATE U5489 ( .I1(n3450), .I2(\registres[26][15] ), .O(n4474) );
  NAND_GATE U5490 ( .I1(n3451), .I2(\registres[27][15] ), .O(n4472) );
  NAND_GATE U5491 ( .I1(n3452), .I2(\registres[10][15] ), .O(n4471) );
  NAND_GATE U5492 ( .I1(n3453), .I2(\registres[18][15] ), .O(n4470) );
  NAND_GATE U5493 ( .I1(n3454), .I2(\registres[5][15] ), .O(n4469) );
  AND5_GATE U5494 ( .I1(n4478), .I2(n4479), .I3(n4480), .I4(n4481), .I5(n4482), 
        .O(n4467) );
  AND4_GATE U5495 ( .I1(n4483), .I2(n4484), .I3(n4485), .I4(n4486), .O(n4482)
         );
  NAND_GATE U5496 ( .I1(n3464), .I2(\registres[28][15] ), .O(n4486) );
  NAND_GATE U5497 ( .I1(n3465), .I2(\registres[29][15] ), .O(n4485) );
  NAND_GATE U5498 ( .I1(n3466), .I2(\registres[12][15] ), .O(n4484) );
  NAND_GATE U5499 ( .I1(n3467), .I2(\registres[20][15] ), .O(n4483) );
  NAND_GATE U5500 ( .I1(n3468), .I2(\registres[1][15] ), .O(n4481) );
  NAND_GATE U5501 ( .I1(n3469), .I2(\registres[9][15] ), .O(n4480) );
  NAND_GATE U5502 ( .I1(n3470), .I2(\registres[11][15] ), .O(n4479) );
  NAND_GATE U5503 ( .I1(n3471), .I2(\registres[13][15] ), .O(n4478) );
  AND5_GATE U5504 ( .I1(n4487), .I2(n4488), .I3(n4489), .I4(n4490), .I5(n4491), 
        .O(n4466) );
  AND4_GATE U5505 ( .I1(n4492), .I2(n4493), .I3(n4494), .I4(n4495), .O(n4491)
         );
  NAND_GATE U5506 ( .I1(n3481), .I2(\registres[17][15] ), .O(n4495) );
  NAND_GATE U5507 ( .I1(n3482), .I2(\registres[19][15] ), .O(n4494) );
  NAND_GATE U5508 ( .I1(n3483), .I2(\registres[21][15] ), .O(n4493) );
  NAND_GATE U5509 ( .I1(n3484), .I2(\registres[6][15] ), .O(n4492) );
  NAND_GATE U5510 ( .I1(n3485), .I2(\registres[7][15] ), .O(n4490) );
  NAND_GATE U5511 ( .I1(n3486), .I2(\registres[30][15] ), .O(n4489) );
  NAND_GATE U5512 ( .I1(n3487), .I2(\registres[31][15] ), .O(n4488) );
  NAND_GATE U5513 ( .I1(n3488), .I2(\registres[14][15] ), .O(n4487) );
  AND4_GATE U5514 ( .I1(n4496), .I2(n4497), .I3(n4498), .I4(n4499), .O(n4465)
         );
  AND4_GATE U5515 ( .I1(n4500), .I2(n4501), .I3(n4502), .I4(n4503), .O(n4499)
         );
  NAND_GATE U5516 ( .I1(n3497), .I2(\registres[22][15] ), .O(n4503) );
  NAND_GATE U5517 ( .I1(n3498), .I2(\registres[15][15] ), .O(n4502) );
  NAND_GATE U5518 ( .I1(n3499), .I2(\registres[23][15] ), .O(n4501) );
  NAND_GATE U5519 ( .I1(n3500), .I2(\registres[4][15] ), .O(n4500) );
  NAND_GATE U5520 ( .I1(n3501), .I2(\registres[8][15] ), .O(n4498) );
  NAND_GATE U5521 ( .I1(n3502), .I2(\registres[2][15] ), .O(n4497) );
  NAND_GATE U5522 ( .I1(n3503), .I2(\registres[16][15] ), .O(n4496) );
  AND_GATE U5523 ( .I1(n4504), .I2(n3432), .O(data_src1[14]) );
  NAND4_GATE U5524 ( .I1(n4505), .I2(n4506), .I3(n4507), .I4(n4508), .O(n4504)
         );
  AND5_GATE U5525 ( .I1(n4509), .I2(n4510), .I3(n4511), .I4(n4512), .I5(n4513), 
        .O(n4508) );
  AND4_GATE U5526 ( .I1(n4514), .I2(n4515), .I3(n4516), .I4(n4517), .O(n4513)
         );
  NAND_GATE U5527 ( .I1(n3447), .I2(\registres[24][14] ), .O(n4517) );
  NAND_GATE U5528 ( .I1(n3448), .I2(\registres[25][14] ), .O(n4516) );
  NAND_GATE U5529 ( .I1(n3449), .I2(\registres[3][14] ), .O(n4515) );
  NAND_GATE U5530 ( .I1(n3450), .I2(\registres[26][14] ), .O(n4514) );
  NAND_GATE U5531 ( .I1(n3451), .I2(\registres[27][14] ), .O(n4512) );
  NAND_GATE U5532 ( .I1(n3452), .I2(\registres[10][14] ), .O(n4511) );
  NAND_GATE U5533 ( .I1(n3453), .I2(\registres[18][14] ), .O(n4510) );
  NAND_GATE U5534 ( .I1(n3454), .I2(\registres[5][14] ), .O(n4509) );
  AND5_GATE U5535 ( .I1(n4518), .I2(n4519), .I3(n4520), .I4(n4521), .I5(n4522), 
        .O(n4507) );
  AND4_GATE U5536 ( .I1(n4523), .I2(n4524), .I3(n4525), .I4(n4526), .O(n4522)
         );
  NAND_GATE U5537 ( .I1(n3464), .I2(\registres[28][14] ), .O(n4526) );
  NAND_GATE U5538 ( .I1(n3465), .I2(\registres[29][14] ), .O(n4525) );
  NAND_GATE U5539 ( .I1(n3466), .I2(\registres[12][14] ), .O(n4524) );
  NAND_GATE U5540 ( .I1(n3467), .I2(\registres[20][14] ), .O(n4523) );
  NAND_GATE U5541 ( .I1(n3468), .I2(\registres[1][14] ), .O(n4521) );
  NAND_GATE U5542 ( .I1(n3469), .I2(\registres[9][14] ), .O(n4520) );
  NAND_GATE U5543 ( .I1(n3470), .I2(\registres[11][14] ), .O(n4519) );
  NAND_GATE U5544 ( .I1(n3471), .I2(\registres[13][14] ), .O(n4518) );
  AND5_GATE U5545 ( .I1(n4527), .I2(n4528), .I3(n4529), .I4(n4530), .I5(n4531), 
        .O(n4506) );
  AND4_GATE U5546 ( .I1(n4532), .I2(n4533), .I3(n4534), .I4(n4535), .O(n4531)
         );
  NAND_GATE U5547 ( .I1(n3481), .I2(\registres[17][14] ), .O(n4535) );
  NAND_GATE U5548 ( .I1(n3482), .I2(\registres[19][14] ), .O(n4534) );
  NAND_GATE U5549 ( .I1(n3483), .I2(\registres[21][14] ), .O(n4533) );
  NAND_GATE U5550 ( .I1(n3484), .I2(\registres[6][14] ), .O(n4532) );
  NAND_GATE U5551 ( .I1(n3485), .I2(\registres[7][14] ), .O(n4530) );
  NAND_GATE U5552 ( .I1(n3486), .I2(\registres[30][14] ), .O(n4529) );
  NAND_GATE U5553 ( .I1(n3487), .I2(\registres[31][14] ), .O(n4528) );
  NAND_GATE U5554 ( .I1(n3488), .I2(\registres[14][14] ), .O(n4527) );
  AND4_GATE U5555 ( .I1(n4536), .I2(n4537), .I3(n4538), .I4(n4539), .O(n4505)
         );
  AND4_GATE U5556 ( .I1(n4540), .I2(n4541), .I3(n4542), .I4(n4543), .O(n4539)
         );
  NAND_GATE U5557 ( .I1(n3497), .I2(\registres[22][14] ), .O(n4543) );
  NAND_GATE U5558 ( .I1(n3498), .I2(\registres[15][14] ), .O(n4542) );
  NAND_GATE U5559 ( .I1(n3499), .I2(\registres[23][14] ), .O(n4541) );
  NAND_GATE U5560 ( .I1(n3500), .I2(\registres[4][14] ), .O(n4540) );
  NAND_GATE U5561 ( .I1(n3501), .I2(\registres[8][14] ), .O(n4538) );
  NAND_GATE U5562 ( .I1(n3502), .I2(\registres[2][14] ), .O(n4537) );
  NAND_GATE U5563 ( .I1(n3503), .I2(\registres[16][14] ), .O(n4536) );
  AND_GATE U5564 ( .I1(n4544), .I2(n3432), .O(data_src1[13]) );
  NAND4_GATE U5565 ( .I1(n4545), .I2(n4546), .I3(n4547), .I4(n4548), .O(n4544)
         );
  AND5_GATE U5566 ( .I1(n4549), .I2(n4550), .I3(n4551), .I4(n4552), .I5(n4553), 
        .O(n4548) );
  AND4_GATE U5567 ( .I1(n4554), .I2(n4555), .I3(n4556), .I4(n4557), .O(n4553)
         );
  NAND_GATE U5568 ( .I1(n3447), .I2(\registres[24][13] ), .O(n4557) );
  NAND_GATE U5569 ( .I1(n3448), .I2(\registres[25][13] ), .O(n4556) );
  NAND_GATE U5570 ( .I1(n3449), .I2(\registres[3][13] ), .O(n4555) );
  NAND_GATE U5571 ( .I1(n3450), .I2(\registres[26][13] ), .O(n4554) );
  NAND_GATE U5572 ( .I1(n3451), .I2(\registres[27][13] ), .O(n4552) );
  NAND_GATE U5573 ( .I1(n3452), .I2(\registres[10][13] ), .O(n4551) );
  NAND_GATE U5574 ( .I1(n3453), .I2(\registres[18][13] ), .O(n4550) );
  NAND_GATE U5575 ( .I1(n3454), .I2(\registres[5][13] ), .O(n4549) );
  AND5_GATE U5576 ( .I1(n4558), .I2(n4559), .I3(n4560), .I4(n4561), .I5(n4562), 
        .O(n4547) );
  AND4_GATE U5577 ( .I1(n4563), .I2(n4564), .I3(n4565), .I4(n4566), .O(n4562)
         );
  NAND_GATE U5578 ( .I1(n3464), .I2(\registres[28][13] ), .O(n4566) );
  NAND_GATE U5579 ( .I1(n3465), .I2(\registres[29][13] ), .O(n4565) );
  NAND_GATE U5580 ( .I1(n3466), .I2(\registres[12][13] ), .O(n4564) );
  NAND_GATE U5581 ( .I1(n3467), .I2(\registres[20][13] ), .O(n4563) );
  NAND_GATE U5582 ( .I1(n3468), .I2(\registres[1][13] ), .O(n4561) );
  NAND_GATE U5583 ( .I1(n3469), .I2(\registres[9][13] ), .O(n4560) );
  NAND_GATE U5584 ( .I1(n3470), .I2(\registres[11][13] ), .O(n4559) );
  NAND_GATE U5585 ( .I1(n3471), .I2(\registres[13][13] ), .O(n4558) );
  AND5_GATE U5586 ( .I1(n4567), .I2(n4568), .I3(n4569), .I4(n4570), .I5(n4571), 
        .O(n4546) );
  AND4_GATE U5587 ( .I1(n4572), .I2(n4573), .I3(n4574), .I4(n4575), .O(n4571)
         );
  NAND_GATE U5588 ( .I1(n3481), .I2(\registres[17][13] ), .O(n4575) );
  NAND_GATE U5589 ( .I1(n3482), .I2(\registres[19][13] ), .O(n4574) );
  NAND_GATE U5590 ( .I1(n3483), .I2(\registres[21][13] ), .O(n4573) );
  NAND_GATE U5591 ( .I1(n3484), .I2(\registres[6][13] ), .O(n4572) );
  NAND_GATE U5592 ( .I1(n3485), .I2(\registres[7][13] ), .O(n4570) );
  NAND_GATE U5593 ( .I1(n3486), .I2(\registres[30][13] ), .O(n4569) );
  NAND_GATE U5594 ( .I1(n3487), .I2(\registres[31][13] ), .O(n4568) );
  NAND_GATE U5595 ( .I1(n3488), .I2(\registres[14][13] ), .O(n4567) );
  AND4_GATE U5596 ( .I1(n4576), .I2(n4577), .I3(n4578), .I4(n4579), .O(n4545)
         );
  AND4_GATE U5597 ( .I1(n4580), .I2(n4581), .I3(n4582), .I4(n4583), .O(n4579)
         );
  NAND_GATE U5598 ( .I1(n3497), .I2(\registres[22][13] ), .O(n4583) );
  NAND_GATE U5599 ( .I1(n3498), .I2(\registres[15][13] ), .O(n4582) );
  NAND_GATE U5600 ( .I1(n3499), .I2(\registres[23][13] ), .O(n4581) );
  NAND_GATE U5601 ( .I1(n3500), .I2(\registres[4][13] ), .O(n4580) );
  NAND_GATE U5602 ( .I1(n3501), .I2(\registres[8][13] ), .O(n4578) );
  NAND_GATE U5603 ( .I1(n3502), .I2(\registres[2][13] ), .O(n4577) );
  NAND_GATE U5604 ( .I1(n3503), .I2(\registres[16][13] ), .O(n4576) );
  AND_GATE U5605 ( .I1(n4584), .I2(n3432), .O(data_src1[12]) );
  NAND4_GATE U5606 ( .I1(n4585), .I2(n4586), .I3(n4587), .I4(n4588), .O(n4584)
         );
  AND5_GATE U5607 ( .I1(n4589), .I2(n4590), .I3(n4591), .I4(n4592), .I5(n4593), 
        .O(n4588) );
  AND4_GATE U5608 ( .I1(n4594), .I2(n4595), .I3(n4596), .I4(n4597), .O(n4593)
         );
  NAND_GATE U5609 ( .I1(n3447), .I2(\registres[24][12] ), .O(n4597) );
  NAND_GATE U5610 ( .I1(n3448), .I2(\registres[25][12] ), .O(n4596) );
  NAND_GATE U5611 ( .I1(n3449), .I2(\registres[3][12] ), .O(n4595) );
  NAND_GATE U5612 ( .I1(n3450), .I2(\registres[26][12] ), .O(n4594) );
  NAND_GATE U5613 ( .I1(n3451), .I2(\registres[27][12] ), .O(n4592) );
  NAND_GATE U5614 ( .I1(n3452), .I2(\registres[10][12] ), .O(n4591) );
  NAND_GATE U5615 ( .I1(n3453), .I2(\registres[18][12] ), .O(n4590) );
  NAND_GATE U5616 ( .I1(n3454), .I2(\registres[5][12] ), .O(n4589) );
  AND5_GATE U5617 ( .I1(n4598), .I2(n4599), .I3(n4600), .I4(n4601), .I5(n4602), 
        .O(n4587) );
  AND4_GATE U5618 ( .I1(n4603), .I2(n4604), .I3(n4605), .I4(n4606), .O(n4602)
         );
  NAND_GATE U5619 ( .I1(n3464), .I2(\registres[28][12] ), .O(n4606) );
  NAND_GATE U5620 ( .I1(n3465), .I2(\registres[29][12] ), .O(n4605) );
  NAND_GATE U5621 ( .I1(n3466), .I2(\registres[12][12] ), .O(n4604) );
  NAND_GATE U5622 ( .I1(n3467), .I2(\registres[20][12] ), .O(n4603) );
  NAND_GATE U5623 ( .I1(n3468), .I2(\registres[1][12] ), .O(n4601) );
  NAND_GATE U5624 ( .I1(n3469), .I2(\registres[9][12] ), .O(n4600) );
  NAND_GATE U5625 ( .I1(n3470), .I2(\registres[11][12] ), .O(n4599) );
  NAND_GATE U5626 ( .I1(n3471), .I2(\registres[13][12] ), .O(n4598) );
  AND5_GATE U5627 ( .I1(n4607), .I2(n4608), .I3(n4609), .I4(n4610), .I5(n4611), 
        .O(n4586) );
  AND4_GATE U5628 ( .I1(n4612), .I2(n4613), .I3(n4614), .I4(n4615), .O(n4611)
         );
  NAND_GATE U5629 ( .I1(n3481), .I2(\registres[17][12] ), .O(n4615) );
  NAND_GATE U5630 ( .I1(n3482), .I2(\registres[19][12] ), .O(n4614) );
  NAND_GATE U5631 ( .I1(n3483), .I2(\registres[21][12] ), .O(n4613) );
  NAND_GATE U5632 ( .I1(n3484), .I2(\registres[6][12] ), .O(n4612) );
  NAND_GATE U5633 ( .I1(n3485), .I2(\registres[7][12] ), .O(n4610) );
  NAND_GATE U5634 ( .I1(n3486), .I2(\registres[30][12] ), .O(n4609) );
  NAND_GATE U5635 ( .I1(n3487), .I2(\registres[31][12] ), .O(n4608) );
  NAND_GATE U5636 ( .I1(n3488), .I2(\registres[14][12] ), .O(n4607) );
  AND4_GATE U5637 ( .I1(n4616), .I2(n4617), .I3(n4618), .I4(n4619), .O(n4585)
         );
  AND4_GATE U5638 ( .I1(n4620), .I2(n4621), .I3(n4622), .I4(n4623), .O(n4619)
         );
  NAND_GATE U5639 ( .I1(n3497), .I2(\registres[22][12] ), .O(n4623) );
  NAND_GATE U5640 ( .I1(n3498), .I2(\registres[15][12] ), .O(n4622) );
  NAND_GATE U5641 ( .I1(n3499), .I2(\registres[23][12] ), .O(n4621) );
  NAND_GATE U5642 ( .I1(n3500), .I2(\registres[4][12] ), .O(n4620) );
  NAND_GATE U5643 ( .I1(n3501), .I2(\registres[8][12] ), .O(n4618) );
  NAND_GATE U5644 ( .I1(n3502), .I2(\registres[2][12] ), .O(n4617) );
  NAND_GATE U5645 ( .I1(n3503), .I2(\registres[16][12] ), .O(n4616) );
  AND_GATE U5646 ( .I1(n4624), .I2(n3432), .O(data_src1[11]) );
  NAND4_GATE U5647 ( .I1(n4625), .I2(n4626), .I3(n4627), .I4(n4628), .O(n4624)
         );
  AND5_GATE U5648 ( .I1(n4629), .I2(n4630), .I3(n4631), .I4(n4632), .I5(n4633), 
        .O(n4628) );
  AND4_GATE U5649 ( .I1(n4634), .I2(n4635), .I3(n4636), .I4(n4637), .O(n4633)
         );
  NAND_GATE U5650 ( .I1(n3447), .I2(\registres[24][11] ), .O(n4637) );
  NAND_GATE U5651 ( .I1(n3448), .I2(\registres[25][11] ), .O(n4636) );
  NAND_GATE U5652 ( .I1(n3449), .I2(\registres[3][11] ), .O(n4635) );
  NAND_GATE U5653 ( .I1(n3450), .I2(\registres[26][11] ), .O(n4634) );
  NAND_GATE U5654 ( .I1(n3451), .I2(\registres[27][11] ), .O(n4632) );
  NAND_GATE U5655 ( .I1(n3452), .I2(\registres[10][11] ), .O(n4631) );
  NAND_GATE U5656 ( .I1(n3453), .I2(\registres[18][11] ), .O(n4630) );
  NAND_GATE U5657 ( .I1(n3454), .I2(\registres[5][11] ), .O(n4629) );
  AND5_GATE U5658 ( .I1(n4638), .I2(n4639), .I3(n4640), .I4(n4641), .I5(n4642), 
        .O(n4627) );
  AND4_GATE U5659 ( .I1(n4643), .I2(n4644), .I3(n4645), .I4(n4646), .O(n4642)
         );
  NAND_GATE U5660 ( .I1(n3464), .I2(\registres[28][11] ), .O(n4646) );
  NAND_GATE U5661 ( .I1(n3465), .I2(\registres[29][11] ), .O(n4645) );
  NAND_GATE U5662 ( .I1(n3466), .I2(\registres[12][11] ), .O(n4644) );
  NAND_GATE U5663 ( .I1(n3467), .I2(\registres[20][11] ), .O(n4643) );
  NAND_GATE U5664 ( .I1(n3468), .I2(\registres[1][11] ), .O(n4641) );
  NAND_GATE U5665 ( .I1(n3469), .I2(\registres[9][11] ), .O(n4640) );
  NAND_GATE U5666 ( .I1(n3470), .I2(\registres[11][11] ), .O(n4639) );
  NAND_GATE U5667 ( .I1(n3471), .I2(\registres[13][11] ), .O(n4638) );
  AND5_GATE U5668 ( .I1(n4647), .I2(n4648), .I3(n4649), .I4(n4650), .I5(n4651), 
        .O(n4626) );
  AND4_GATE U5669 ( .I1(n4652), .I2(n4653), .I3(n4654), .I4(n4655), .O(n4651)
         );
  NAND_GATE U5670 ( .I1(n3481), .I2(\registres[17][11] ), .O(n4655) );
  NAND_GATE U5671 ( .I1(n3482), .I2(\registres[19][11] ), .O(n4654) );
  NAND_GATE U5672 ( .I1(n3483), .I2(\registres[21][11] ), .O(n4653) );
  NAND_GATE U5673 ( .I1(n3484), .I2(\registres[6][11] ), .O(n4652) );
  NAND_GATE U5674 ( .I1(n3485), .I2(\registres[7][11] ), .O(n4650) );
  NAND_GATE U5675 ( .I1(n3486), .I2(\registres[30][11] ), .O(n4649) );
  NAND_GATE U5676 ( .I1(n3487), .I2(\registres[31][11] ), .O(n4648) );
  NAND_GATE U5677 ( .I1(n3488), .I2(\registres[14][11] ), .O(n4647) );
  AND4_GATE U5678 ( .I1(n4656), .I2(n4657), .I3(n4658), .I4(n4659), .O(n4625)
         );
  AND4_GATE U5679 ( .I1(n4660), .I2(n4661), .I3(n4662), .I4(n4663), .O(n4659)
         );
  NAND_GATE U5680 ( .I1(n3497), .I2(\registres[22][11] ), .O(n4663) );
  NAND_GATE U5681 ( .I1(n3498), .I2(\registres[15][11] ), .O(n4662) );
  NAND_GATE U5682 ( .I1(n3499), .I2(\registres[23][11] ), .O(n4661) );
  NAND_GATE U5683 ( .I1(n3500), .I2(\registres[4][11] ), .O(n4660) );
  NAND_GATE U5684 ( .I1(n3501), .I2(\registres[8][11] ), .O(n4658) );
  NAND_GATE U5685 ( .I1(n3502), .I2(\registres[2][11] ), .O(n4657) );
  NAND_GATE U5686 ( .I1(n3503), .I2(\registres[16][11] ), .O(n4656) );
  AND_GATE U5687 ( .I1(n4664), .I2(n3432), .O(data_src1[10]) );
  NAND4_GATE U5688 ( .I1(n4665), .I2(n4666), .I3(n4667), .I4(n4668), .O(n4664)
         );
  AND5_GATE U5689 ( .I1(n4669), .I2(n4670), .I3(n4671), .I4(n4672), .I5(n4673), 
        .O(n4668) );
  AND4_GATE U5690 ( .I1(n4674), .I2(n4675), .I3(n4676), .I4(n4677), .O(n4673)
         );
  NAND_GATE U5691 ( .I1(n3447), .I2(\registres[24][10] ), .O(n4677) );
  NAND_GATE U5692 ( .I1(n3448), .I2(\registres[25][10] ), .O(n4676) );
  NAND_GATE U5693 ( .I1(n3449), .I2(\registres[3][10] ), .O(n4675) );
  NAND_GATE U5694 ( .I1(n3450), .I2(\registres[26][10] ), .O(n4674) );
  NAND_GATE U5695 ( .I1(n3451), .I2(\registres[27][10] ), .O(n4672) );
  NAND_GATE U5696 ( .I1(n3452), .I2(\registres[10][10] ), .O(n4671) );
  NAND_GATE U5697 ( .I1(n3453), .I2(\registres[18][10] ), .O(n4670) );
  NAND_GATE U5698 ( .I1(n3454), .I2(\registres[5][10] ), .O(n4669) );
  AND5_GATE U5699 ( .I1(n4678), .I2(n4679), .I3(n4680), .I4(n4681), .I5(n4682), 
        .O(n4667) );
  AND4_GATE U5700 ( .I1(n4683), .I2(n4684), .I3(n4685), .I4(n4686), .O(n4682)
         );
  NAND_GATE U5701 ( .I1(n3464), .I2(\registres[28][10] ), .O(n4686) );
  NAND_GATE U5702 ( .I1(n3465), .I2(\registres[29][10] ), .O(n4685) );
  NAND_GATE U5703 ( .I1(n3466), .I2(\registres[12][10] ), .O(n4684) );
  NAND_GATE U5704 ( .I1(n3467), .I2(\registres[20][10] ), .O(n4683) );
  NAND_GATE U5705 ( .I1(n3468), .I2(\registres[1][10] ), .O(n4681) );
  NAND_GATE U5706 ( .I1(n3469), .I2(\registres[9][10] ), .O(n4680) );
  NAND_GATE U5707 ( .I1(n3470), .I2(\registres[11][10] ), .O(n4679) );
  NAND_GATE U5708 ( .I1(n3471), .I2(\registres[13][10] ), .O(n4678) );
  AND5_GATE U5709 ( .I1(n4687), .I2(n4688), .I3(n4689), .I4(n4690), .I5(n4691), 
        .O(n4666) );
  AND4_GATE U5710 ( .I1(n4692), .I2(n4693), .I3(n4694), .I4(n4695), .O(n4691)
         );
  NAND_GATE U5711 ( .I1(n3481), .I2(\registres[17][10] ), .O(n4695) );
  NAND_GATE U5712 ( .I1(n3482), .I2(\registres[19][10] ), .O(n4694) );
  NAND_GATE U5713 ( .I1(n3483), .I2(\registres[21][10] ), .O(n4693) );
  NAND_GATE U5714 ( .I1(n3484), .I2(\registres[6][10] ), .O(n4692) );
  NAND_GATE U5715 ( .I1(n3485), .I2(\registres[7][10] ), .O(n4690) );
  NAND_GATE U5716 ( .I1(n3486), .I2(\registres[30][10] ), .O(n4689) );
  NAND_GATE U5717 ( .I1(n3487), .I2(\registres[31][10] ), .O(n4688) );
  NAND_GATE U5718 ( .I1(n3488), .I2(\registres[14][10] ), .O(n4687) );
  AND4_GATE U5719 ( .I1(n4696), .I2(n4697), .I3(n4698), .I4(n4699), .O(n4665)
         );
  AND4_GATE U5720 ( .I1(n4700), .I2(n4701), .I3(n4702), .I4(n4703), .O(n4699)
         );
  NAND_GATE U5721 ( .I1(n3497), .I2(\registres[22][10] ), .O(n4703) );
  NAND_GATE U5722 ( .I1(n3498), .I2(\registres[15][10] ), .O(n4702) );
  NAND_GATE U5723 ( .I1(n3499), .I2(\registres[23][10] ), .O(n4701) );
  NAND_GATE U5724 ( .I1(n3500), .I2(\registres[4][10] ), .O(n4700) );
  NAND_GATE U5725 ( .I1(n3501), .I2(\registres[8][10] ), .O(n4698) );
  NAND_GATE U5726 ( .I1(n3502), .I2(\registres[2][10] ), .O(n4697) );
  NAND_GATE U5727 ( .I1(n3503), .I2(\registres[16][10] ), .O(n4696) );
  AND_GATE U5728 ( .I1(n4704), .I2(n3432), .O(data_src1[0]) );
  NAND_GATE U5729 ( .I1(n3501), .I2(n8), .O(n3432) );
  NAND4_GATE U5730 ( .I1(n4705), .I2(n4706), .I3(n4707), .I4(n4708), .O(n4704)
         );
  AND5_GATE U5731 ( .I1(n4709), .I2(n4710), .I3(n4711), .I4(n4712), .I5(n4713), 
        .O(n4708) );
  AND4_GATE U5732 ( .I1(n4714), .I2(n4715), .I3(n4716), .I4(n4717), .O(n4713)
         );
  NAND_GATE U5733 ( .I1(n3447), .I2(\registres[24][0] ), .O(n4717) );
  AND_GATE U5734 ( .I1(n4718), .I2(n4719), .O(n3447) );
  NAND_GATE U5735 ( .I1(n3448), .I2(\registres[25][0] ), .O(n4716) );
  AND_GATE U5736 ( .I1(n4720), .I2(n4718), .O(n3448) );
  NAND_GATE U5737 ( .I1(n3449), .I2(\registres[3][0] ), .O(n4715) );
  AND_GATE U5738 ( .I1(n4721), .I2(n4722), .O(n3449) );
  NAND_GATE U5739 ( .I1(n3450), .I2(\registres[26][0] ), .O(n4714) );
  AND_GATE U5740 ( .I1(n4721), .I2(n4719), .O(n3450) );
  NAND_GATE U5741 ( .I1(n3451), .I2(\registres[27][0] ), .O(n4712) );
  AND_GATE U5742 ( .I1(n4721), .I2(n4720), .O(n3451) );
  NAND_GATE U5743 ( .I1(n3452), .I2(\registres[10][0] ), .O(n4711) );
  AND_GATE U5744 ( .I1(n4723), .I2(n4721), .O(n3452) );
  NAND_GATE U5745 ( .I1(n3453), .I2(\registres[18][0] ), .O(n4710) );
  AND_GATE U5746 ( .I1(n4724), .I2(n4721), .O(n3453) );
  NAND_GATE U5747 ( .I1(n3454), .I2(\registres[5][0] ), .O(n4709) );
  AND_GATE U5748 ( .I1(n4725), .I2(n4722), .O(n3454) );
  AND5_GATE U5749 ( .I1(n4726), .I2(n4727), .I3(n4728), .I4(n4729), .I5(n4730), 
        .O(n4707) );
  AND4_GATE U5750 ( .I1(n4731), .I2(n4732), .I3(n4733), .I4(n4734), .O(n4730)
         );
  NAND_GATE U5751 ( .I1(n3464), .I2(\registres[28][0] ), .O(n4734) );
  AND_GATE U5752 ( .I1(n4725), .I2(n4719), .O(n3464) );
  NAND_GATE U5753 ( .I1(n3465), .I2(\registres[29][0] ), .O(n4733) );
  AND_GATE U5754 ( .I1(n4725), .I2(n4720), .O(n3465) );
  NAND_GATE U5755 ( .I1(n3466), .I2(\registres[12][0] ), .O(n4732) );
  AND_GATE U5756 ( .I1(n4725), .I2(n4723), .O(n3466) );
  NAND_GATE U5757 ( .I1(n3467), .I2(\registres[20][0] ), .O(n4731) );
  AND_GATE U5758 ( .I1(n4725), .I2(n4724), .O(n3467) );
  NAND_GATE U5759 ( .I1(n3468), .I2(\registres[1][0] ), .O(n4729) );
  AND_GATE U5760 ( .I1(n4735), .I2(n4718), .O(n3468) );
  NAND_GATE U5761 ( .I1(n3469), .I2(\registres[9][0] ), .O(n4728) );
  AND_GATE U5762 ( .I1(n4736), .I2(n4718), .O(n3469) );
  NAND_GATE U5763 ( .I1(n3470), .I2(\registres[11][0] ), .O(n4727) );
  AND_GATE U5764 ( .I1(n4736), .I2(n4721), .O(n3470) );
  NAND_GATE U5765 ( .I1(n3471), .I2(\registres[13][0] ), .O(n4726) );
  AND_GATE U5766 ( .I1(n4736), .I2(n4725), .O(n3471) );
  AND5_GATE U5767 ( .I1(n4737), .I2(n4738), .I3(n4739), .I4(n4740), .I5(n4741), 
        .O(n4706) );
  AND4_GATE U5768 ( .I1(n4742), .I2(n4743), .I3(n4744), .I4(n4745), .O(n4741)
         );
  NAND_GATE U5769 ( .I1(n3481), .I2(\registres[17][0] ), .O(n4745) );
  AND_GATE U5770 ( .I1(n4746), .I2(n4718), .O(n3481) );
  NAND_GATE U5771 ( .I1(n3482), .I2(\registres[19][0] ), .O(n4744) );
  AND_GATE U5772 ( .I1(n4746), .I2(n4721), .O(n3482) );
  NOR_GATE U5773 ( .I1(n6), .I2(reg_src1[2]), .O(n4721) );
  NAND_GATE U5774 ( .I1(n3483), .I2(\registres[21][0] ), .O(n4743) );
  AND_GATE U5775 ( .I1(n4746), .I2(n4725), .O(n3483) );
  NOR_GATE U5776 ( .I1(n7), .I2(reg_src1[1]), .O(n4725) );
  NAND_GATE U5777 ( .I1(n3484), .I2(\registres[6][0] ), .O(n4742) );
  AND_GATE U5778 ( .I1(n4747), .I2(n4748), .O(n3484) );
  NAND_GATE U5779 ( .I1(n3485), .I2(\registres[7][0] ), .O(n4740) );
  AND_GATE U5780 ( .I1(n4747), .I2(n4722), .O(n3485) );
  AND_GATE U5781 ( .I1(n4735), .I2(reg_src1[0]), .O(n4722) );
  NAND_GATE U5782 ( .I1(n3486), .I2(\registres[30][0] ), .O(n4739) );
  AND_GATE U5783 ( .I1(n4747), .I2(n4719), .O(n3486) );
  AND_GATE U5784 ( .I1(n4749), .I2(n5), .O(n4719) );
  NAND_GATE U5785 ( .I1(n3487), .I2(\registres[31][0] ), .O(n4738) );
  AND_GATE U5786 ( .I1(n4747), .I2(n4720), .O(n3487) );
  AND_GATE U5787 ( .I1(reg_src1[0]), .I2(n4749), .O(n4720) );
  NOR_GATE U5788 ( .I1(n9), .I2(n8), .O(n4749) );
  NAND_GATE U5789 ( .I1(n3488), .I2(\registres[14][0] ), .O(n4737) );
  AND_GATE U5790 ( .I1(n4747), .I2(n4723), .O(n3488) );
  NOR3_GATE U5791 ( .I1(reg_src1[0]), .I2(reg_src1[4]), .I3(n8), .O(n4723) );
  AND4_GATE U5792 ( .I1(n4750), .I2(n4751), .I3(n4752), .I4(n4753), .O(n4705)
         );
  AND4_GATE U5793 ( .I1(n4754), .I2(n4755), .I3(n4756), .I4(n4757), .O(n4753)
         );
  NAND_GATE U5794 ( .I1(n3497), .I2(\registres[22][0] ), .O(n4757) );
  AND_GATE U5795 ( .I1(n4747), .I2(n4724), .O(n3497) );
  NOR3_GATE U5796 ( .I1(reg_src1[0]), .I2(reg_src1[3]), .I3(n9), .O(n4724) );
  NAND_GATE U5797 ( .I1(n3498), .I2(\registres[15][0] ), .O(n4756) );
  AND_GATE U5798 ( .I1(n4747), .I2(n4736), .O(n3498) );
  NOR3_GATE U5799 ( .I1(n8), .I2(reg_src1[4]), .I3(n5), .O(n4736) );
  NAND_GATE U5800 ( .I1(n3499), .I2(\registres[23][0] ), .O(n4755) );
  AND_GATE U5801 ( .I1(n4747), .I2(n4746), .O(n3499) );
  NOR3_GATE U5802 ( .I1(n9), .I2(reg_src1[3]), .I3(n5), .O(n4746) );
  NOR_GATE U5803 ( .I1(n7), .I2(n6), .O(n4747) );
  NAND_GATE U5804 ( .I1(n3500), .I2(\registres[4][0] ), .O(n4754) );
  AND_GATE U5805 ( .I1(n4748), .I2(n6), .O(n3500) );
  NAND_GATE U5806 ( .I1(n3501), .I2(\registres[8][0] ), .O(n4752) );
  AND_GATE U5807 ( .I1(n4758), .I2(n9), .O(n3501) );
  NAND_GATE U5808 ( .I1(n3502), .I2(\registres[2][0] ), .O(n4751) );
  AND_GATE U5809 ( .I1(n4748), .I2(n7), .O(n3502) );
  AND_GATE U5810 ( .I1(n4735), .I2(n5), .O(n4748) );
  NOR_GATE U5811 ( .I1(reg_src1[4]), .I2(reg_src1[3]), .O(n4735) );
  NAND_GATE U5812 ( .I1(n3503), .I2(\registres[16][0] ), .O(n4750) );
  AND_GATE U5813 ( .I1(n4758), .I2(n8), .O(n3503) );
  AND_GATE U5814 ( .I1(n4718), .I2(n5), .O(n4758) );
  NOR_GATE U5815 ( .I1(reg_src1[2]), .I2(reg_src1[1]), .O(n4718) );
  INV_GATE U3 ( .I1(reset), .O(n1) );
  INV_GATE U4 ( .I1(reg_dest[4]), .O(n2) );
  INV_GATE U5 ( .I1(reg_dest[1]), .O(n3) );
  INV_GATE U6 ( .I1(reg_dest[0]), .O(n4) );
  INV_GATE U7 ( .I1(reg_src1[0]), .O(n5) );
  INV_GATE U8 ( .I1(reg_src1[1]), .O(n6) );
  INV_GATE U9 ( .I1(reg_src1[2]), .O(n7) );
  INV_GATE U10 ( .I1(reg_src1[3]), .O(n8) );
  INV_GATE U11 ( .I1(reg_src1[4]), .O(n9) );
  INV_GATE U12 ( .I1(reg_src2[0]), .O(n10) );
  INV_GATE U13 ( .I1(reg_src2[1]), .O(n11) );
  INV_GATE U14 ( .I1(reg_src2[2]), .O(n12) );
  INV_GATE U15 ( .I1(reg_src2[3]), .O(n13) );
  INV_GATE U16 ( .I1(reg_src2[4]), .O(n14) );
endmodule


module renvoi ( adr1, adr2, use1, use2, data1, data2, alea, DI_level, DI_adr, 
        DI_ecr, DI_data, EX_level, EX_adr, EX_ecr, EX_data, MEM_level, MEM_adr, 
        MEM_ecr, MEM_data, interrupt, write_data, write_adr, write_GPR, 
        write_SCP, read_adr1, read_adr2, read_data1_GPR, read_data2_GPR, 
        read_data1_SCP, read_data2_SCP );
  input [5:0] adr1;
  input [5:0] adr2;
  output [31:0] data1;
  output [31:0] data2;
  input [1:0] DI_level;
  input [5:0] DI_adr;
  input [31:0] DI_data;
  input [1:0] EX_level;
  input [5:0] EX_adr;
  input [31:0] EX_data;
  input [1:0] MEM_level;
  input [5:0] MEM_adr;
  input [31:0] MEM_data;
  output [31:0] write_data;
  output [4:0] write_adr;
  output [4:0] read_adr1;
  output [4:0] read_adr2;
  input [31:0] read_data1_GPR;
  input [31:0] read_data2_GPR;
  input [31:0] read_data1_SCP;
  input [31:0] read_data2_SCP;
  input use1, use2, DI_ecr, EX_ecr, MEM_ecr, interrupt;
  output alea, write_GPR, write_SCP;
  wire   N250, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484;
  assign write_data[31] = MEM_data[31];
  assign write_data[30] = MEM_data[30];
  assign write_data[29] = MEM_data[29];
  assign write_data[28] = MEM_data[28];
  assign write_data[27] = MEM_data[27];
  assign write_data[26] = MEM_data[26];
  assign write_data[25] = MEM_data[25];
  assign write_data[24] = MEM_data[24];
  assign write_data[23] = MEM_data[23];
  assign write_data[22] = MEM_data[22];
  assign write_data[21] = MEM_data[21];
  assign write_data[20] = MEM_data[20];
  assign write_data[19] = MEM_data[19];
  assign write_data[18] = MEM_data[18];
  assign write_data[17] = MEM_data[17];
  assign write_data[16] = MEM_data[16];
  assign write_data[15] = MEM_data[15];
  assign write_data[14] = MEM_data[14];
  assign write_data[13] = MEM_data[13];
  assign write_data[12] = MEM_data[12];
  assign write_data[11] = MEM_data[11];
  assign write_data[10] = MEM_data[10];
  assign write_data[9] = MEM_data[9];
  assign write_data[8] = MEM_data[8];
  assign write_data[7] = MEM_data[7];
  assign write_data[6] = MEM_data[6];
  assign write_data[5] = MEM_data[5];
  assign write_data[4] = MEM_data[4];
  assign write_data[3] = MEM_data[3];
  assign write_data[2] = MEM_data[2];
  assign write_data[1] = MEM_data[1];
  assign write_data[0] = MEM_data[0];
  assign write_adr[4] = MEM_adr[4];
  assign write_adr[3] = MEM_adr[3];
  assign write_adr[2] = MEM_adr[2];
  assign write_adr[1] = MEM_adr[1];
  assign write_adr[0] = MEM_adr[0];
  assign read_adr1[4] = adr1[4];
  assign read_adr1[3] = adr1[3];
  assign read_adr1[2] = adr1[2];
  assign read_adr1[1] = adr1[1];
  assign read_adr1[0] = adr1[0];
  assign read_adr2[4] = adr2[4];
  assign read_adr2[3] = adr2[3];
  assign read_adr2[2] = adr2[2];
  assign read_adr2[1] = adr2[1];
  assign read_adr2[0] = adr2[0];
  assign N250 = EX_level[1];

  AND_GATE U3 ( .I1(MEM_ecr), .I2(MEM_adr[5]), .O(write_SCP) );
  NOR3_GATE U4 ( .I1(n1), .I2(interrupt), .I3(MEM_adr[5]), .O(write_GPR) );
  INV_GATE U5 ( .I1(MEM_ecr), .O(n1) );
  NAND5_GATE U6 ( .I1(n2), .I2(n3), .I3(n4), .I4(n5), .I5(n6), .O(data2[9]) );
  NAND_GATE U7 ( .I1(EX_data[9]), .I2(n7), .O(n6) );
  NAND_GATE U8 ( .I1(MEM_data[9]), .I2(n8), .O(n5) );
  NAND_GATE U9 ( .I1(read_data2_SCP[9]), .I2(n9), .O(n4) );
  NAND_GATE U10 ( .I1(DI_data[9]), .I2(n10), .O(n3) );
  NAND_GATE U11 ( .I1(read_data2_GPR[9]), .I2(n11), .O(n2) );
  NAND5_GATE U12 ( .I1(n12), .I2(n13), .I3(n14), .I4(n15), .I5(n16), .O(
        data2[8]) );
  NAND_GATE U13 ( .I1(EX_data[8]), .I2(n7), .O(n16) );
  NAND_GATE U14 ( .I1(MEM_data[8]), .I2(n8), .O(n15) );
  NAND_GATE U15 ( .I1(read_data2_SCP[8]), .I2(n9), .O(n14) );
  NAND_GATE U16 ( .I1(DI_data[8]), .I2(n10), .O(n13) );
  NAND_GATE U17 ( .I1(read_data2_GPR[8]), .I2(n11), .O(n12) );
  NAND5_GATE U18 ( .I1(n17), .I2(n18), .I3(n19), .I4(n20), .I5(n21), .O(
        data2[7]) );
  NAND_GATE U19 ( .I1(EX_data[7]), .I2(n7), .O(n21) );
  NAND_GATE U20 ( .I1(MEM_data[7]), .I2(n8), .O(n20) );
  NAND_GATE U21 ( .I1(read_data2_SCP[7]), .I2(n9), .O(n19) );
  NAND_GATE U22 ( .I1(DI_data[7]), .I2(n10), .O(n18) );
  NAND_GATE U23 ( .I1(read_data2_GPR[7]), .I2(n11), .O(n17) );
  NAND5_GATE U24 ( .I1(n22), .I2(n23), .I3(n24), .I4(n25), .I5(n26), .O(
        data2[6]) );
  NAND_GATE U25 ( .I1(EX_data[6]), .I2(n7), .O(n26) );
  NAND_GATE U26 ( .I1(MEM_data[6]), .I2(n8), .O(n25) );
  NAND_GATE U27 ( .I1(read_data2_SCP[6]), .I2(n9), .O(n24) );
  NAND_GATE U28 ( .I1(DI_data[6]), .I2(n10), .O(n23) );
  NAND_GATE U29 ( .I1(read_data2_GPR[6]), .I2(n11), .O(n22) );
  NAND5_GATE U30 ( .I1(n27), .I2(n28), .I3(n29), .I4(n30), .I5(n31), .O(
        data2[5]) );
  NAND_GATE U31 ( .I1(EX_data[5]), .I2(n7), .O(n31) );
  NAND_GATE U32 ( .I1(MEM_data[5]), .I2(n8), .O(n30) );
  NAND_GATE U33 ( .I1(read_data2_SCP[5]), .I2(n9), .O(n29) );
  NAND_GATE U34 ( .I1(DI_data[5]), .I2(n10), .O(n28) );
  NAND_GATE U35 ( .I1(read_data2_GPR[5]), .I2(n11), .O(n27) );
  NAND5_GATE U36 ( .I1(n32), .I2(n33), .I3(n34), .I4(n35), .I5(n36), .O(
        data2[4]) );
  NAND_GATE U37 ( .I1(EX_data[4]), .I2(n7), .O(n36) );
  NAND_GATE U38 ( .I1(MEM_data[4]), .I2(n8), .O(n35) );
  NAND_GATE U39 ( .I1(read_data2_SCP[4]), .I2(n9), .O(n34) );
  NAND_GATE U40 ( .I1(DI_data[4]), .I2(n10), .O(n33) );
  NAND_GATE U41 ( .I1(read_data2_GPR[4]), .I2(n11), .O(n32) );
  NAND5_GATE U42 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .I5(n41), .O(
        data2[3]) );
  NAND_GATE U43 ( .I1(EX_data[3]), .I2(n7), .O(n41) );
  NAND_GATE U44 ( .I1(MEM_data[3]), .I2(n8), .O(n40) );
  NAND_GATE U45 ( .I1(read_data2_SCP[3]), .I2(n9), .O(n39) );
  NAND_GATE U46 ( .I1(DI_data[3]), .I2(n10), .O(n38) );
  NAND_GATE U47 ( .I1(read_data2_GPR[3]), .I2(n11), .O(n37) );
  NAND5_GATE U48 ( .I1(n42), .I2(n43), .I3(n44), .I4(n45), .I5(n46), .O(
        data2[31]) );
  NAND_GATE U49 ( .I1(EX_data[31]), .I2(n7), .O(n46) );
  NAND_GATE U50 ( .I1(MEM_data[31]), .I2(n8), .O(n45) );
  NAND_GATE U51 ( .I1(read_data2_SCP[31]), .I2(n9), .O(n44) );
  NAND_GATE U52 ( .I1(DI_data[31]), .I2(n10), .O(n43) );
  NAND_GATE U53 ( .I1(read_data2_GPR[31]), .I2(n11), .O(n42) );
  NAND5_GATE U54 ( .I1(n47), .I2(n48), .I3(n49), .I4(n50), .I5(n51), .O(
        data2[30]) );
  NAND_GATE U55 ( .I1(EX_data[30]), .I2(n7), .O(n51) );
  NAND_GATE U56 ( .I1(MEM_data[30]), .I2(n8), .O(n50) );
  NAND_GATE U57 ( .I1(read_data2_SCP[30]), .I2(n9), .O(n49) );
  NAND_GATE U58 ( .I1(DI_data[30]), .I2(n10), .O(n48) );
  NAND_GATE U59 ( .I1(read_data2_GPR[30]), .I2(n11), .O(n47) );
  NAND5_GATE U60 ( .I1(n52), .I2(n53), .I3(n54), .I4(n55), .I5(n56), .O(
        data2[2]) );
  NAND_GATE U61 ( .I1(EX_data[2]), .I2(n7), .O(n56) );
  NAND_GATE U62 ( .I1(MEM_data[2]), .I2(n8), .O(n55) );
  NAND_GATE U63 ( .I1(read_data2_SCP[2]), .I2(n9), .O(n54) );
  NAND_GATE U64 ( .I1(DI_data[2]), .I2(n10), .O(n53) );
  NAND_GATE U65 ( .I1(read_data2_GPR[2]), .I2(n11), .O(n52) );
  NAND5_GATE U66 ( .I1(n57), .I2(n58), .I3(n59), .I4(n60), .I5(n61), .O(
        data2[29]) );
  NAND_GATE U67 ( .I1(EX_data[29]), .I2(n7), .O(n61) );
  NAND_GATE U68 ( .I1(MEM_data[29]), .I2(n8), .O(n60) );
  NAND_GATE U69 ( .I1(read_data2_SCP[29]), .I2(n9), .O(n59) );
  NAND_GATE U70 ( .I1(DI_data[29]), .I2(n10), .O(n58) );
  NAND_GATE U71 ( .I1(read_data2_GPR[29]), .I2(n11), .O(n57) );
  NAND5_GATE U72 ( .I1(n62), .I2(n63), .I3(n64), .I4(n65), .I5(n66), .O(
        data2[28]) );
  NAND_GATE U73 ( .I1(EX_data[28]), .I2(n7), .O(n66) );
  NAND_GATE U74 ( .I1(MEM_data[28]), .I2(n8), .O(n65) );
  NAND_GATE U75 ( .I1(read_data2_SCP[28]), .I2(n9), .O(n64) );
  NAND_GATE U76 ( .I1(DI_data[28]), .I2(n10), .O(n63) );
  NAND_GATE U77 ( .I1(read_data2_GPR[28]), .I2(n11), .O(n62) );
  NAND5_GATE U78 ( .I1(n67), .I2(n68), .I3(n69), .I4(n70), .I5(n71), .O(
        data2[27]) );
  NAND_GATE U79 ( .I1(EX_data[27]), .I2(n7), .O(n71) );
  NAND_GATE U80 ( .I1(MEM_data[27]), .I2(n8), .O(n70) );
  NAND_GATE U81 ( .I1(read_data2_SCP[27]), .I2(n9), .O(n69) );
  NAND_GATE U82 ( .I1(DI_data[27]), .I2(n10), .O(n68) );
  NAND_GATE U83 ( .I1(read_data2_GPR[27]), .I2(n11), .O(n67) );
  NAND5_GATE U84 ( .I1(n72), .I2(n73), .I3(n74), .I4(n75), .I5(n76), .O(
        data2[26]) );
  NAND_GATE U85 ( .I1(EX_data[26]), .I2(n7), .O(n76) );
  NAND_GATE U86 ( .I1(MEM_data[26]), .I2(n8), .O(n75) );
  NAND_GATE U87 ( .I1(read_data2_SCP[26]), .I2(n9), .O(n74) );
  NAND_GATE U88 ( .I1(DI_data[26]), .I2(n10), .O(n73) );
  NAND_GATE U89 ( .I1(read_data2_GPR[26]), .I2(n11), .O(n72) );
  NAND5_GATE U90 ( .I1(n77), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(
        data2[25]) );
  NAND_GATE U91 ( .I1(EX_data[25]), .I2(n7), .O(n81) );
  NAND_GATE U92 ( .I1(MEM_data[25]), .I2(n8), .O(n80) );
  NAND_GATE U93 ( .I1(read_data2_SCP[25]), .I2(n9), .O(n79) );
  NAND_GATE U94 ( .I1(DI_data[25]), .I2(n10), .O(n78) );
  NAND_GATE U95 ( .I1(read_data2_GPR[25]), .I2(n11), .O(n77) );
  NAND5_GATE U96 ( .I1(n82), .I2(n83), .I3(n84), .I4(n85), .I5(n86), .O(
        data2[24]) );
  NAND_GATE U97 ( .I1(EX_data[24]), .I2(n7), .O(n86) );
  NAND_GATE U98 ( .I1(MEM_data[24]), .I2(n8), .O(n85) );
  NAND_GATE U99 ( .I1(read_data2_SCP[24]), .I2(n9), .O(n84) );
  NAND_GATE U100 ( .I1(DI_data[24]), .I2(n10), .O(n83) );
  NAND_GATE U101 ( .I1(read_data2_GPR[24]), .I2(n11), .O(n82) );
  NAND5_GATE U102 ( .I1(n87), .I2(n88), .I3(n89), .I4(n90), .I5(n91), .O(
        data2[23]) );
  NAND_GATE U103 ( .I1(EX_data[23]), .I2(n7), .O(n91) );
  NAND_GATE U104 ( .I1(MEM_data[23]), .I2(n8), .O(n90) );
  NAND_GATE U105 ( .I1(read_data2_SCP[23]), .I2(n9), .O(n89) );
  NAND_GATE U106 ( .I1(DI_data[23]), .I2(n10), .O(n88) );
  NAND_GATE U107 ( .I1(read_data2_GPR[23]), .I2(n11), .O(n87) );
  NAND5_GATE U108 ( .I1(n92), .I2(n93), .I3(n94), .I4(n95), .I5(n96), .O(
        data2[22]) );
  NAND_GATE U109 ( .I1(EX_data[22]), .I2(n7), .O(n96) );
  NAND_GATE U110 ( .I1(MEM_data[22]), .I2(n8), .O(n95) );
  NAND_GATE U111 ( .I1(read_data2_SCP[22]), .I2(n9), .O(n94) );
  NAND_GATE U112 ( .I1(DI_data[22]), .I2(n10), .O(n93) );
  NAND_GATE U113 ( .I1(read_data2_GPR[22]), .I2(n11), .O(n92) );
  NAND5_GATE U114 ( .I1(n97), .I2(n98), .I3(n99), .I4(n100), .I5(n101), .O(
        data2[21]) );
  NAND_GATE U115 ( .I1(EX_data[21]), .I2(n7), .O(n101) );
  NAND_GATE U116 ( .I1(MEM_data[21]), .I2(n8), .O(n100) );
  NAND_GATE U117 ( .I1(read_data2_SCP[21]), .I2(n9), .O(n99) );
  NAND_GATE U118 ( .I1(DI_data[21]), .I2(n10), .O(n98) );
  NAND_GATE U119 ( .I1(read_data2_GPR[21]), .I2(n11), .O(n97) );
  NAND5_GATE U120 ( .I1(n102), .I2(n103), .I3(n104), .I4(n105), .I5(n106), .O(
        data2[20]) );
  NAND_GATE U121 ( .I1(EX_data[20]), .I2(n7), .O(n106) );
  NAND_GATE U122 ( .I1(MEM_data[20]), .I2(n8), .O(n105) );
  NAND_GATE U123 ( .I1(read_data2_SCP[20]), .I2(n9), .O(n104) );
  NAND_GATE U124 ( .I1(DI_data[20]), .I2(n10), .O(n103) );
  NAND_GATE U125 ( .I1(read_data2_GPR[20]), .I2(n11), .O(n102) );
  NAND5_GATE U126 ( .I1(n107), .I2(n108), .I3(n109), .I4(n110), .I5(n111), .O(
        data2[1]) );
  NAND_GATE U127 ( .I1(EX_data[1]), .I2(n7), .O(n111) );
  NAND_GATE U128 ( .I1(MEM_data[1]), .I2(n8), .O(n110) );
  NAND_GATE U129 ( .I1(read_data2_SCP[1]), .I2(n9), .O(n109) );
  NAND_GATE U130 ( .I1(DI_data[1]), .I2(n10), .O(n108) );
  NAND_GATE U131 ( .I1(read_data2_GPR[1]), .I2(n11), .O(n107) );
  NAND5_GATE U132 ( .I1(n112), .I2(n113), .I3(n114), .I4(n115), .I5(n116), .O(
        data2[19]) );
  NAND_GATE U133 ( .I1(EX_data[19]), .I2(n7), .O(n116) );
  NAND_GATE U134 ( .I1(MEM_data[19]), .I2(n8), .O(n115) );
  NAND_GATE U135 ( .I1(read_data2_SCP[19]), .I2(n9), .O(n114) );
  NAND_GATE U136 ( .I1(DI_data[19]), .I2(n10), .O(n113) );
  NAND_GATE U137 ( .I1(read_data2_GPR[19]), .I2(n11), .O(n112) );
  NAND5_GATE U138 ( .I1(n117), .I2(n118), .I3(n119), .I4(n120), .I5(n121), .O(
        data2[18]) );
  NAND_GATE U139 ( .I1(EX_data[18]), .I2(n7), .O(n121) );
  NAND_GATE U140 ( .I1(MEM_data[18]), .I2(n8), .O(n120) );
  NAND_GATE U141 ( .I1(read_data2_SCP[18]), .I2(n9), .O(n119) );
  NAND_GATE U142 ( .I1(DI_data[18]), .I2(n10), .O(n118) );
  NAND_GATE U143 ( .I1(read_data2_GPR[18]), .I2(n11), .O(n117) );
  NAND5_GATE U144 ( .I1(n122), .I2(n123), .I3(n124), .I4(n125), .I5(n126), .O(
        data2[17]) );
  NAND_GATE U145 ( .I1(EX_data[17]), .I2(n7), .O(n126) );
  NAND_GATE U146 ( .I1(MEM_data[17]), .I2(n8), .O(n125) );
  NAND_GATE U147 ( .I1(read_data2_SCP[17]), .I2(n9), .O(n124) );
  NAND_GATE U148 ( .I1(DI_data[17]), .I2(n10), .O(n123) );
  NAND_GATE U149 ( .I1(read_data2_GPR[17]), .I2(n11), .O(n122) );
  NAND5_GATE U150 ( .I1(n127), .I2(n128), .I3(n129), .I4(n130), .I5(n131), .O(
        data2[16]) );
  NAND_GATE U151 ( .I1(EX_data[16]), .I2(n7), .O(n131) );
  NAND_GATE U152 ( .I1(MEM_data[16]), .I2(n8), .O(n130) );
  NAND_GATE U153 ( .I1(read_data2_SCP[16]), .I2(n9), .O(n129) );
  NAND_GATE U154 ( .I1(DI_data[16]), .I2(n10), .O(n128) );
  NAND_GATE U155 ( .I1(read_data2_GPR[16]), .I2(n11), .O(n127) );
  NAND5_GATE U156 ( .I1(n132), .I2(n133), .I3(n134), .I4(n135), .I5(n136), .O(
        data2[15]) );
  NAND_GATE U157 ( .I1(EX_data[15]), .I2(n7), .O(n136) );
  NAND_GATE U158 ( .I1(MEM_data[15]), .I2(n8), .O(n135) );
  NAND_GATE U159 ( .I1(read_data2_SCP[15]), .I2(n9), .O(n134) );
  NAND_GATE U160 ( .I1(DI_data[15]), .I2(n10), .O(n133) );
  NAND_GATE U161 ( .I1(read_data2_GPR[15]), .I2(n11), .O(n132) );
  NAND5_GATE U162 ( .I1(n137), .I2(n138), .I3(n139), .I4(n140), .I5(n141), .O(
        data2[14]) );
  NAND_GATE U163 ( .I1(EX_data[14]), .I2(n7), .O(n141) );
  NAND_GATE U164 ( .I1(MEM_data[14]), .I2(n8), .O(n140) );
  NAND_GATE U165 ( .I1(read_data2_SCP[14]), .I2(n9), .O(n139) );
  NAND_GATE U166 ( .I1(DI_data[14]), .I2(n10), .O(n138) );
  NAND_GATE U167 ( .I1(read_data2_GPR[14]), .I2(n11), .O(n137) );
  NAND5_GATE U168 ( .I1(n142), .I2(n143), .I3(n144), .I4(n145), .I5(n146), .O(
        data2[13]) );
  NAND_GATE U169 ( .I1(EX_data[13]), .I2(n7), .O(n146) );
  NAND_GATE U170 ( .I1(MEM_data[13]), .I2(n8), .O(n145) );
  NAND_GATE U171 ( .I1(read_data2_SCP[13]), .I2(n9), .O(n144) );
  NAND_GATE U172 ( .I1(DI_data[13]), .I2(n10), .O(n143) );
  NAND_GATE U173 ( .I1(read_data2_GPR[13]), .I2(n11), .O(n142) );
  NAND5_GATE U174 ( .I1(n147), .I2(n148), .I3(n149), .I4(n150), .I5(n151), .O(
        data2[12]) );
  NAND_GATE U175 ( .I1(EX_data[12]), .I2(n7), .O(n151) );
  NAND_GATE U176 ( .I1(MEM_data[12]), .I2(n8), .O(n150) );
  NAND_GATE U177 ( .I1(read_data2_SCP[12]), .I2(n9), .O(n149) );
  NAND_GATE U178 ( .I1(DI_data[12]), .I2(n10), .O(n148) );
  NAND_GATE U179 ( .I1(read_data2_GPR[12]), .I2(n11), .O(n147) );
  NAND5_GATE U180 ( .I1(n152), .I2(n153), .I3(n154), .I4(n155), .I5(n156), .O(
        data2[11]) );
  NAND_GATE U181 ( .I1(EX_data[11]), .I2(n7), .O(n156) );
  NAND_GATE U182 ( .I1(MEM_data[11]), .I2(n8), .O(n155) );
  NAND_GATE U183 ( .I1(read_data2_SCP[11]), .I2(n9), .O(n154) );
  NAND_GATE U184 ( .I1(DI_data[11]), .I2(n10), .O(n153) );
  NAND_GATE U185 ( .I1(read_data2_GPR[11]), .I2(n11), .O(n152) );
  NAND5_GATE U186 ( .I1(n157), .I2(n158), .I3(n159), .I4(n160), .I5(n161), .O(
        data2[10]) );
  NAND_GATE U187 ( .I1(EX_data[10]), .I2(n7), .O(n161) );
  NAND_GATE U188 ( .I1(MEM_data[10]), .I2(n8), .O(n160) );
  NAND_GATE U189 ( .I1(read_data2_SCP[10]), .I2(n9), .O(n159) );
  NAND_GATE U190 ( .I1(DI_data[10]), .I2(n10), .O(n158) );
  NAND_GATE U191 ( .I1(read_data2_GPR[10]), .I2(n11), .O(n157) );
  NAND5_GATE U192 ( .I1(n162), .I2(n163), .I3(n164), .I4(n165), .I5(n166), .O(
        data2[0]) );
  NAND_GATE U193 ( .I1(EX_data[0]), .I2(n7), .O(n166) );
  NAND_GATE U194 ( .I1(MEM_data[0]), .I2(n8), .O(n165) );
  NAND_GATE U195 ( .I1(read_data2_SCP[0]), .I2(n9), .O(n164) );
  AND_GATE U196 ( .I1(n167), .I2(adr2[5]), .O(n9) );
  NAND_GATE U197 ( .I1(DI_data[0]), .I2(n10), .O(n163) );
  NOR3_GATE U198 ( .I1(n7), .I2(n8), .I3(n167), .O(n10) );
  NAND_GATE U199 ( .I1(read_data2_GPR[0]), .I2(n11), .O(n162) );
  AND_GATE U200 ( .I1(n167), .I2(n168), .O(n11) );
  NOR_GATE U201 ( .I1(n169), .I2(n170), .O(n167) );
  NAND5_GATE U202 ( .I1(n171), .I2(n172), .I3(n173), .I4(n174), .I5(n175), .O(
        data1[9]) );
  NAND_GATE U203 ( .I1(n176), .I2(EX_data[9]), .O(n175) );
  NAND_GATE U204 ( .I1(n177), .I2(MEM_data[9]), .O(n174) );
  NAND_GATE U205 ( .I1(read_data1_SCP[9]), .I2(n178), .O(n173) );
  NAND_GATE U206 ( .I1(n179), .I2(DI_data[9]), .O(n172) );
  NAND_GATE U207 ( .I1(read_data1_GPR[9]), .I2(n180), .O(n171) );
  NAND5_GATE U208 ( .I1(n181), .I2(n182), .I3(n183), .I4(n184), .I5(n185), .O(
        data1[8]) );
  NAND_GATE U209 ( .I1(n176), .I2(EX_data[8]), .O(n185) );
  NAND_GATE U210 ( .I1(n177), .I2(MEM_data[8]), .O(n184) );
  NAND_GATE U211 ( .I1(read_data1_SCP[8]), .I2(n178), .O(n183) );
  NAND_GATE U212 ( .I1(n179), .I2(DI_data[8]), .O(n182) );
  NAND_GATE U213 ( .I1(read_data1_GPR[8]), .I2(n180), .O(n181) );
  NAND5_GATE U214 ( .I1(n186), .I2(n187), .I3(n188), .I4(n189), .I5(n190), .O(
        data1[7]) );
  NAND_GATE U215 ( .I1(n176), .I2(EX_data[7]), .O(n190) );
  NAND_GATE U216 ( .I1(n177), .I2(MEM_data[7]), .O(n189) );
  NAND_GATE U217 ( .I1(read_data1_SCP[7]), .I2(n178), .O(n188) );
  NAND_GATE U218 ( .I1(n179), .I2(DI_data[7]), .O(n187) );
  NAND_GATE U219 ( .I1(read_data1_GPR[7]), .I2(n180), .O(n186) );
  NAND5_GATE U220 ( .I1(n191), .I2(n192), .I3(n193), .I4(n194), .I5(n195), .O(
        data1[6]) );
  NAND_GATE U221 ( .I1(n176), .I2(EX_data[6]), .O(n195) );
  NAND_GATE U222 ( .I1(n177), .I2(MEM_data[6]), .O(n194) );
  NAND_GATE U223 ( .I1(read_data1_SCP[6]), .I2(n178), .O(n193) );
  NAND_GATE U224 ( .I1(n179), .I2(DI_data[6]), .O(n192) );
  NAND_GATE U225 ( .I1(read_data1_GPR[6]), .I2(n180), .O(n191) );
  NAND5_GATE U226 ( .I1(n196), .I2(n197), .I3(n198), .I4(n199), .I5(n200), .O(
        data1[5]) );
  NAND_GATE U227 ( .I1(n176), .I2(EX_data[5]), .O(n200) );
  NAND_GATE U228 ( .I1(n177), .I2(MEM_data[5]), .O(n199) );
  NAND_GATE U229 ( .I1(read_data1_SCP[5]), .I2(n178), .O(n198) );
  NAND_GATE U230 ( .I1(n179), .I2(DI_data[5]), .O(n197) );
  NAND_GATE U231 ( .I1(read_data1_GPR[5]), .I2(n180), .O(n196) );
  NAND5_GATE U232 ( .I1(n201), .I2(n202), .I3(n203), .I4(n204), .I5(n205), .O(
        data1[4]) );
  NAND_GATE U233 ( .I1(n176), .I2(EX_data[4]), .O(n205) );
  NAND_GATE U234 ( .I1(n177), .I2(MEM_data[4]), .O(n204) );
  NAND_GATE U235 ( .I1(read_data1_SCP[4]), .I2(n178), .O(n203) );
  NAND_GATE U236 ( .I1(n179), .I2(DI_data[4]), .O(n202) );
  NAND_GATE U237 ( .I1(read_data1_GPR[4]), .I2(n180), .O(n201) );
  NAND5_GATE U238 ( .I1(n206), .I2(n207), .I3(n208), .I4(n209), .I5(n210), .O(
        data1[3]) );
  NAND_GATE U239 ( .I1(n176), .I2(EX_data[3]), .O(n210) );
  NAND_GATE U240 ( .I1(n177), .I2(MEM_data[3]), .O(n209) );
  NAND_GATE U241 ( .I1(read_data1_SCP[3]), .I2(n178), .O(n208) );
  NAND_GATE U242 ( .I1(n179), .I2(DI_data[3]), .O(n207) );
  NAND_GATE U243 ( .I1(read_data1_GPR[3]), .I2(n180), .O(n206) );
  NAND5_GATE U244 ( .I1(n211), .I2(n212), .I3(n213), .I4(n214), .I5(n215), .O(
        data1[31]) );
  NAND_GATE U245 ( .I1(n176), .I2(EX_data[31]), .O(n215) );
  NAND_GATE U246 ( .I1(n177), .I2(MEM_data[31]), .O(n214) );
  NAND_GATE U247 ( .I1(read_data1_SCP[31]), .I2(n178), .O(n213) );
  NAND_GATE U248 ( .I1(n179), .I2(DI_data[31]), .O(n212) );
  NAND_GATE U249 ( .I1(read_data1_GPR[31]), .I2(n180), .O(n211) );
  NAND5_GATE U250 ( .I1(n216), .I2(n217), .I3(n218), .I4(n219), .I5(n220), .O(
        data1[30]) );
  NAND_GATE U251 ( .I1(n176), .I2(EX_data[30]), .O(n220) );
  NAND_GATE U252 ( .I1(n177), .I2(MEM_data[30]), .O(n219) );
  NAND_GATE U253 ( .I1(read_data1_SCP[30]), .I2(n178), .O(n218) );
  NAND_GATE U254 ( .I1(n179), .I2(DI_data[30]), .O(n217) );
  NAND_GATE U255 ( .I1(read_data1_GPR[30]), .I2(n180), .O(n216) );
  NAND5_GATE U256 ( .I1(n221), .I2(n222), .I3(n223), .I4(n224), .I5(n225), .O(
        data1[2]) );
  NAND_GATE U257 ( .I1(n176), .I2(EX_data[2]), .O(n225) );
  NAND_GATE U258 ( .I1(n177), .I2(MEM_data[2]), .O(n224) );
  NAND_GATE U259 ( .I1(read_data1_SCP[2]), .I2(n178), .O(n223) );
  NAND_GATE U260 ( .I1(n179), .I2(DI_data[2]), .O(n222) );
  NAND_GATE U261 ( .I1(read_data1_GPR[2]), .I2(n180), .O(n221) );
  NAND5_GATE U262 ( .I1(n226), .I2(n227), .I3(n228), .I4(n229), .I5(n230), .O(
        data1[29]) );
  NAND_GATE U263 ( .I1(n176), .I2(EX_data[29]), .O(n230) );
  NAND_GATE U264 ( .I1(n177), .I2(MEM_data[29]), .O(n229) );
  NAND_GATE U265 ( .I1(read_data1_SCP[29]), .I2(n178), .O(n228) );
  NAND_GATE U266 ( .I1(n179), .I2(DI_data[29]), .O(n227) );
  NAND_GATE U267 ( .I1(read_data1_GPR[29]), .I2(n180), .O(n226) );
  NAND5_GATE U268 ( .I1(n231), .I2(n232), .I3(n233), .I4(n234), .I5(n235), .O(
        data1[28]) );
  NAND_GATE U269 ( .I1(n176), .I2(EX_data[28]), .O(n235) );
  NAND_GATE U270 ( .I1(n177), .I2(MEM_data[28]), .O(n234) );
  NAND_GATE U271 ( .I1(read_data1_SCP[28]), .I2(n178), .O(n233) );
  NAND_GATE U272 ( .I1(n179), .I2(DI_data[28]), .O(n232) );
  NAND_GATE U273 ( .I1(read_data1_GPR[28]), .I2(n180), .O(n231) );
  NAND5_GATE U274 ( .I1(n236), .I2(n237), .I3(n238), .I4(n239), .I5(n240), .O(
        data1[27]) );
  NAND_GATE U275 ( .I1(n176), .I2(EX_data[27]), .O(n240) );
  NAND_GATE U276 ( .I1(n177), .I2(MEM_data[27]), .O(n239) );
  NAND_GATE U277 ( .I1(read_data1_SCP[27]), .I2(n178), .O(n238) );
  NAND_GATE U278 ( .I1(n179), .I2(DI_data[27]), .O(n237) );
  NAND_GATE U279 ( .I1(read_data1_GPR[27]), .I2(n180), .O(n236) );
  NAND5_GATE U280 ( .I1(n241), .I2(n242), .I3(n243), .I4(n244), .I5(n245), .O(
        data1[26]) );
  NAND_GATE U281 ( .I1(n176), .I2(EX_data[26]), .O(n245) );
  NAND_GATE U282 ( .I1(n177), .I2(MEM_data[26]), .O(n244) );
  NAND_GATE U283 ( .I1(read_data1_SCP[26]), .I2(n178), .O(n243) );
  NAND_GATE U284 ( .I1(n179), .I2(DI_data[26]), .O(n242) );
  NAND_GATE U285 ( .I1(read_data1_GPR[26]), .I2(n180), .O(n241) );
  NAND5_GATE U286 ( .I1(n246), .I2(n247), .I3(n248), .I4(n249), .I5(n250), .O(
        data1[25]) );
  NAND_GATE U287 ( .I1(n176), .I2(EX_data[25]), .O(n250) );
  NAND_GATE U288 ( .I1(n177), .I2(MEM_data[25]), .O(n249) );
  NAND_GATE U289 ( .I1(read_data1_SCP[25]), .I2(n178), .O(n248) );
  NAND_GATE U290 ( .I1(n179), .I2(DI_data[25]), .O(n247) );
  NAND_GATE U291 ( .I1(read_data1_GPR[25]), .I2(n180), .O(n246) );
  NAND5_GATE U292 ( .I1(n251), .I2(n252), .I3(n253), .I4(n254), .I5(n255), .O(
        data1[24]) );
  NAND_GATE U293 ( .I1(n176), .I2(EX_data[24]), .O(n255) );
  NAND_GATE U294 ( .I1(n177), .I2(MEM_data[24]), .O(n254) );
  NAND_GATE U295 ( .I1(read_data1_SCP[24]), .I2(n178), .O(n253) );
  NAND_GATE U296 ( .I1(n179), .I2(DI_data[24]), .O(n252) );
  NAND_GATE U297 ( .I1(read_data1_GPR[24]), .I2(n180), .O(n251) );
  NAND5_GATE U298 ( .I1(n256), .I2(n257), .I3(n258), .I4(n259), .I5(n260), .O(
        data1[23]) );
  NAND_GATE U299 ( .I1(n176), .I2(EX_data[23]), .O(n260) );
  NAND_GATE U300 ( .I1(n177), .I2(MEM_data[23]), .O(n259) );
  NAND_GATE U301 ( .I1(read_data1_SCP[23]), .I2(n178), .O(n258) );
  NAND_GATE U302 ( .I1(n179), .I2(DI_data[23]), .O(n257) );
  NAND_GATE U303 ( .I1(read_data1_GPR[23]), .I2(n180), .O(n256) );
  NAND5_GATE U304 ( .I1(n261), .I2(n262), .I3(n263), .I4(n264), .I5(n265), .O(
        data1[22]) );
  NAND_GATE U305 ( .I1(n176), .I2(EX_data[22]), .O(n265) );
  NAND_GATE U306 ( .I1(n177), .I2(MEM_data[22]), .O(n264) );
  NAND_GATE U307 ( .I1(read_data1_SCP[22]), .I2(n178), .O(n263) );
  NAND_GATE U308 ( .I1(n179), .I2(DI_data[22]), .O(n262) );
  NAND_GATE U309 ( .I1(read_data1_GPR[22]), .I2(n180), .O(n261) );
  NAND5_GATE U310 ( .I1(n266), .I2(n267), .I3(n268), .I4(n269), .I5(n270), .O(
        data1[21]) );
  NAND_GATE U311 ( .I1(n176), .I2(EX_data[21]), .O(n270) );
  NAND_GATE U312 ( .I1(n177), .I2(MEM_data[21]), .O(n269) );
  NAND_GATE U313 ( .I1(read_data1_SCP[21]), .I2(n178), .O(n268) );
  NAND_GATE U314 ( .I1(n179), .I2(DI_data[21]), .O(n267) );
  NAND_GATE U315 ( .I1(read_data1_GPR[21]), .I2(n180), .O(n266) );
  NAND5_GATE U316 ( .I1(n271), .I2(n272), .I3(n273), .I4(n274), .I5(n275), .O(
        data1[20]) );
  NAND_GATE U317 ( .I1(n176), .I2(EX_data[20]), .O(n275) );
  NAND_GATE U318 ( .I1(n177), .I2(MEM_data[20]), .O(n274) );
  NAND_GATE U319 ( .I1(read_data1_SCP[20]), .I2(n178), .O(n273) );
  NAND_GATE U320 ( .I1(n179), .I2(DI_data[20]), .O(n272) );
  NAND_GATE U321 ( .I1(read_data1_GPR[20]), .I2(n180), .O(n271) );
  NAND5_GATE U322 ( .I1(n276), .I2(n277), .I3(n278), .I4(n279), .I5(n280), .O(
        data1[1]) );
  NAND_GATE U323 ( .I1(n176), .I2(EX_data[1]), .O(n280) );
  NAND_GATE U324 ( .I1(n177), .I2(MEM_data[1]), .O(n279) );
  NAND_GATE U325 ( .I1(read_data1_SCP[1]), .I2(n178), .O(n278) );
  NAND_GATE U326 ( .I1(n179), .I2(DI_data[1]), .O(n277) );
  NAND_GATE U327 ( .I1(read_data1_GPR[1]), .I2(n180), .O(n276) );
  NAND5_GATE U328 ( .I1(n281), .I2(n282), .I3(n283), .I4(n284), .I5(n285), .O(
        data1[19]) );
  NAND_GATE U329 ( .I1(n176), .I2(EX_data[19]), .O(n285) );
  NAND_GATE U330 ( .I1(n177), .I2(MEM_data[19]), .O(n284) );
  NAND_GATE U331 ( .I1(read_data1_SCP[19]), .I2(n178), .O(n283) );
  NAND_GATE U332 ( .I1(n179), .I2(DI_data[19]), .O(n282) );
  NAND_GATE U333 ( .I1(read_data1_GPR[19]), .I2(n180), .O(n281) );
  NAND5_GATE U334 ( .I1(n286), .I2(n287), .I3(n288), .I4(n289), .I5(n290), .O(
        data1[18]) );
  NAND_GATE U335 ( .I1(n176), .I2(EX_data[18]), .O(n290) );
  NAND_GATE U336 ( .I1(n177), .I2(MEM_data[18]), .O(n289) );
  NAND_GATE U337 ( .I1(read_data1_SCP[18]), .I2(n178), .O(n288) );
  NAND_GATE U338 ( .I1(n179), .I2(DI_data[18]), .O(n287) );
  NAND_GATE U339 ( .I1(read_data1_GPR[18]), .I2(n180), .O(n286) );
  NAND5_GATE U340 ( .I1(n291), .I2(n292), .I3(n293), .I4(n294), .I5(n295), .O(
        data1[17]) );
  NAND_GATE U341 ( .I1(n176), .I2(EX_data[17]), .O(n295) );
  NAND_GATE U342 ( .I1(n177), .I2(MEM_data[17]), .O(n294) );
  NAND_GATE U343 ( .I1(read_data1_SCP[17]), .I2(n178), .O(n293) );
  NAND_GATE U344 ( .I1(n179), .I2(DI_data[17]), .O(n292) );
  NAND_GATE U345 ( .I1(read_data1_GPR[17]), .I2(n180), .O(n291) );
  NAND5_GATE U346 ( .I1(n296), .I2(n297), .I3(n298), .I4(n299), .I5(n300), .O(
        data1[16]) );
  NAND_GATE U347 ( .I1(n176), .I2(EX_data[16]), .O(n300) );
  NAND_GATE U348 ( .I1(n177), .I2(MEM_data[16]), .O(n299) );
  NAND_GATE U349 ( .I1(read_data1_SCP[16]), .I2(n178), .O(n298) );
  NAND_GATE U350 ( .I1(n179), .I2(DI_data[16]), .O(n297) );
  NAND_GATE U351 ( .I1(read_data1_GPR[16]), .I2(n180), .O(n296) );
  NAND5_GATE U352 ( .I1(n301), .I2(n302), .I3(n303), .I4(n304), .I5(n305), .O(
        data1[15]) );
  NAND_GATE U353 ( .I1(n176), .I2(EX_data[15]), .O(n305) );
  NAND_GATE U354 ( .I1(n177), .I2(MEM_data[15]), .O(n304) );
  NAND_GATE U355 ( .I1(read_data1_SCP[15]), .I2(n178), .O(n303) );
  NAND_GATE U356 ( .I1(n179), .I2(DI_data[15]), .O(n302) );
  NAND_GATE U357 ( .I1(read_data1_GPR[15]), .I2(n180), .O(n301) );
  NAND5_GATE U358 ( .I1(n306), .I2(n307), .I3(n308), .I4(n309), .I5(n310), .O(
        data1[14]) );
  NAND_GATE U359 ( .I1(n176), .I2(EX_data[14]), .O(n310) );
  NAND_GATE U360 ( .I1(n177), .I2(MEM_data[14]), .O(n309) );
  NAND_GATE U361 ( .I1(read_data1_SCP[14]), .I2(n178), .O(n308) );
  NAND_GATE U362 ( .I1(n179), .I2(DI_data[14]), .O(n307) );
  NAND_GATE U363 ( .I1(read_data1_GPR[14]), .I2(n180), .O(n306) );
  NAND5_GATE U364 ( .I1(n311), .I2(n312), .I3(n313), .I4(n314), .I5(n315), .O(
        data1[13]) );
  NAND_GATE U365 ( .I1(n176), .I2(EX_data[13]), .O(n315) );
  NAND_GATE U366 ( .I1(n177), .I2(MEM_data[13]), .O(n314) );
  NAND_GATE U367 ( .I1(read_data1_SCP[13]), .I2(n178), .O(n313) );
  NAND_GATE U368 ( .I1(n179), .I2(DI_data[13]), .O(n312) );
  NAND_GATE U369 ( .I1(read_data1_GPR[13]), .I2(n180), .O(n311) );
  NAND5_GATE U370 ( .I1(n316), .I2(n317), .I3(n318), .I4(n319), .I5(n320), .O(
        data1[12]) );
  NAND_GATE U371 ( .I1(n176), .I2(EX_data[12]), .O(n320) );
  NAND_GATE U372 ( .I1(n177), .I2(MEM_data[12]), .O(n319) );
  NAND_GATE U373 ( .I1(read_data1_SCP[12]), .I2(n178), .O(n318) );
  NAND_GATE U374 ( .I1(n179), .I2(DI_data[12]), .O(n317) );
  NAND_GATE U375 ( .I1(read_data1_GPR[12]), .I2(n180), .O(n316) );
  NAND5_GATE U376 ( .I1(n321), .I2(n322), .I3(n323), .I4(n324), .I5(n325), .O(
        data1[11]) );
  NAND_GATE U377 ( .I1(n176), .I2(EX_data[11]), .O(n325) );
  NAND_GATE U378 ( .I1(n177), .I2(MEM_data[11]), .O(n324) );
  NAND_GATE U379 ( .I1(read_data1_SCP[11]), .I2(n178), .O(n323) );
  NAND_GATE U380 ( .I1(n179), .I2(DI_data[11]), .O(n322) );
  NAND_GATE U381 ( .I1(read_data1_GPR[11]), .I2(n180), .O(n321) );
  NAND5_GATE U382 ( .I1(n326), .I2(n327), .I3(n328), .I4(n329), .I5(n330), .O(
        data1[10]) );
  NAND_GATE U383 ( .I1(n176), .I2(EX_data[10]), .O(n330) );
  NAND_GATE U384 ( .I1(n177), .I2(MEM_data[10]), .O(n329) );
  NAND_GATE U385 ( .I1(read_data1_SCP[10]), .I2(n178), .O(n328) );
  NAND_GATE U386 ( .I1(n179), .I2(DI_data[10]), .O(n327) );
  NAND_GATE U387 ( .I1(read_data1_GPR[10]), .I2(n180), .O(n326) );
  NAND5_GATE U388 ( .I1(n331), .I2(n332), .I3(n333), .I4(n334), .I5(n335), .O(
        data1[0]) );
  NAND_GATE U389 ( .I1(n176), .I2(EX_data[0]), .O(n335) );
  NAND_GATE U390 ( .I1(n177), .I2(MEM_data[0]), .O(n334) );
  NAND_GATE U391 ( .I1(read_data1_SCP[0]), .I2(n178), .O(n333) );
  AND_GATE U392 ( .I1(n336), .I2(adr1[5]), .O(n178) );
  NAND_GATE U393 ( .I1(n179), .I2(DI_data[0]), .O(n332) );
  NOR3_GATE U394 ( .I1(n176), .I2(n177), .I3(n336), .O(n179) );
  NAND_GATE U395 ( .I1(read_data1_GPR[0]), .I2(n180), .O(n331) );
  AND_GATE U396 ( .I1(n336), .I2(n337), .O(n180) );
  NOR_GATE U397 ( .I1(n338), .I2(n339), .O(n336) );
  NAND3_GATE U398 ( .I1(n340), .I2(n341), .I3(n342), .O(alea) );
  OR_GATE U399 ( .I1(N250), .I2(n343), .O(n342) );
  NOR_GATE U400 ( .I1(n176), .I2(n7), .O(n343) );
  NOR_GATE U401 ( .I1(n169), .I2(n344), .O(n7) );
  INV_GATE U402 ( .I1(n345), .O(n169) );
  NOR_GATE U403 ( .I1(n338), .I2(n346), .O(n176) );
  INV_GATE U404 ( .I1(n347), .O(n338) );
  NAND_GATE U405 ( .I1(n348), .I2(n349), .O(n341) );
  NAND_GATE U406 ( .I1(n350), .I2(n351), .O(n349) );
  OR_GATE U407 ( .I1(n344), .I2(n345), .O(n351) );
  OR_GATE U408 ( .I1(n346), .I2(n347), .O(n350) );
  NAND_GATE U409 ( .I1(DI_level[1]), .I2(DI_level[0]), .O(n348) );
  OR3_GATE U410 ( .I1(MEM_level[1]), .I2(MEM_level[0]), .I3(n352), .O(n340) );
  NOR_GATE U411 ( .I1(n177), .I2(n8), .O(n352) );
  NOR_GATE U412 ( .I1(n170), .I2(n345), .O(n8) );
  AND_GATE U413 ( .I1(n353), .I2(n354), .O(n345) );
  NAND5_GATE U414 ( .I1(MEM_ecr), .I2(n355), .I3(n356), .I4(n357), .I5(n358), 
        .O(n353) );
  AND5_GATE U415 ( .I1(n359), .I2(n360), .I3(n361), .I4(n362), .I5(n363), .O(
        n358) );
  AND4_GATE U416 ( .I1(n364), .I2(n365), .I3(n366), .I4(n367), .O(n363) );
  OR_GATE U417 ( .I1(n368), .I2(adr2[1]), .O(n367) );
  OR_GATE U418 ( .I1(n369), .I2(MEM_adr[1]), .O(n366) );
  OR_GATE U419 ( .I1(n370), .I2(adr2[2]), .O(n365) );
  OR_GATE U420 ( .I1(n371), .I2(MEM_adr[2]), .O(n364) );
  OR_GATE U421 ( .I1(n372), .I2(adr2[3]), .O(n362) );
  OR_GATE U422 ( .I1(n373), .I2(MEM_adr[3]), .O(n361) );
  OR_GATE U423 ( .I1(n374), .I2(adr2[4]), .O(n360) );
  OR_GATE U424 ( .I1(n375), .I2(MEM_adr[4]), .O(n359) );
  AND4_GATE U425 ( .I1(n376), .I2(n377), .I3(n378), .I4(n379), .O(n357) );
  OR_GATE U426 ( .I1(n168), .I2(MEM_adr[5]), .O(n379) );
  OR_GATE U427 ( .I1(n380), .I2(adr2[5]), .O(n378) );
  OR_GATE U428 ( .I1(n381), .I2(adr2[0]), .O(n377) );
  OR_GATE U429 ( .I1(n382), .I2(MEM_adr[0]), .O(n376) );
  INV_GATE U430 ( .I1(n344), .O(n170) );
  AND_GATE U431 ( .I1(n354), .I2(n383), .O(n344) );
  OR_GATE U432 ( .I1(n355), .I2(n384), .O(n383) );
  NAND5_GATE U433 ( .I1(n385), .I2(n386), .I3(n387), .I4(n388), .I5(n389), .O(
        n355) );
  AND3_GATE U434 ( .I1(n390), .I2(n391), .I3(EX_ecr), .O(n389) );
  OR_GATE U435 ( .I1(n382), .I2(EX_adr[0]), .O(n391) );
  OR_GATE U436 ( .I1(n392), .I2(adr2[0]), .O(n390) );
  AND4_GATE U437 ( .I1(n393), .I2(n394), .I3(n395), .I4(n396), .O(n388) );
  OR_GATE U438 ( .I1(n369), .I2(EX_adr[1]), .O(n396) );
  OR_GATE U439 ( .I1(n397), .I2(adr2[1]), .O(n395) );
  OR_GATE U440 ( .I1(n371), .I2(EX_adr[2]), .O(n394) );
  OR_GATE U441 ( .I1(n398), .I2(adr2[2]), .O(n393) );
  AND4_GATE U442 ( .I1(n399), .I2(n400), .I3(n401), .I4(n402), .O(n387) );
  OR_GATE U443 ( .I1(n168), .I2(EX_adr[5]), .O(n402) );
  OR_GATE U444 ( .I1(n403), .I2(adr2[5]), .O(n401) );
  OR_GATE U445 ( .I1(n373), .I2(EX_adr[3]), .O(n400) );
  OR_GATE U446 ( .I1(n404), .I2(adr2[3]), .O(n399) );
  OR_GATE U447 ( .I1(n375), .I2(EX_adr[4]), .O(n386) );
  OR_GATE U448 ( .I1(n405), .I2(adr2[4]), .O(n385) );
  NAND5_GATE U449 ( .I1(DI_ecr), .I2(n356), .I3(n406), .I4(n407), .I5(n408), 
        .O(n354) );
  AND4_GATE U450 ( .I1(n409), .I2(n410), .I3(n411), .I4(n412), .O(n408) );
  OR_GATE U451 ( .I1(n371), .I2(DI_adr[2]), .O(n412) );
  OR_GATE U452 ( .I1(n413), .I2(adr2[2]), .O(n411) );
  OR_GATE U453 ( .I1(n373), .I2(DI_adr[3]), .O(n410) );
  OR_GATE U454 ( .I1(n414), .I2(adr2[3]), .O(n409) );
  AND4_GATE U455 ( .I1(n415), .I2(n416), .I3(n417), .I4(n418), .O(n407) );
  OR_GATE U456 ( .I1(n375), .I2(DI_adr[4]), .O(n418) );
  OR_GATE U457 ( .I1(n419), .I2(adr2[4]), .O(n417) );
  OR_GATE U458 ( .I1(n168), .I2(DI_adr[5]), .O(n416) );
  INV_GATE U459 ( .I1(adr2[5]), .O(n168) );
  OR_GATE U460 ( .I1(n420), .I2(adr2[5]), .O(n415) );
  AND4_GATE U461 ( .I1(n421), .I2(n422), .I3(n423), .I4(n424), .O(n406) );
  OR_GATE U462 ( .I1(n382), .I2(DI_adr[0]), .O(n424) );
  OR_GATE U463 ( .I1(n425), .I2(adr2[0]), .O(n423) );
  OR_GATE U464 ( .I1(n369), .I2(DI_adr[1]), .O(n422) );
  OR_GATE U465 ( .I1(n426), .I2(adr2[1]), .O(n421) );
  INV_GATE U466 ( .I1(n384), .O(n356) );
  NAND_GATE U467 ( .I1(use2), .I2(n427), .O(n384) );
  NAND5_GATE U468 ( .I1(n375), .I2(n373), .I3(n371), .I4(n369), .I5(n382), .O(
        n427) );
  INV_GATE U469 ( .I1(adr2[0]), .O(n382) );
  INV_GATE U470 ( .I1(adr2[1]), .O(n369) );
  INV_GATE U471 ( .I1(adr2[2]), .O(n371) );
  INV_GATE U472 ( .I1(adr2[3]), .O(n373) );
  INV_GATE U473 ( .I1(adr2[4]), .O(n375) );
  NOR_GATE U474 ( .I1(n339), .I2(n347), .O(n177) );
  AND_GATE U475 ( .I1(n428), .I2(n429), .O(n347) );
  NAND5_GATE U476 ( .I1(MEM_ecr), .I2(n430), .I3(n431), .I4(n432), .I5(n433), 
        .O(n428) );
  AND5_GATE U477 ( .I1(n434), .I2(n435), .I3(n436), .I4(n437), .I5(n438), .O(
        n433) );
  AND4_GATE U478 ( .I1(n439), .I2(n440), .I3(n441), .I4(n442), .O(n438) );
  OR_GATE U479 ( .I1(n368), .I2(adr1[1]), .O(n442) );
  INV_GATE U480 ( .I1(MEM_adr[1]), .O(n368) );
  OR_GATE U481 ( .I1(n443), .I2(MEM_adr[1]), .O(n441) );
  OR_GATE U482 ( .I1(n370), .I2(adr1[2]), .O(n440) );
  INV_GATE U483 ( .I1(MEM_adr[2]), .O(n370) );
  OR_GATE U484 ( .I1(n444), .I2(MEM_adr[2]), .O(n439) );
  OR_GATE U485 ( .I1(n372), .I2(adr1[3]), .O(n437) );
  INV_GATE U486 ( .I1(MEM_adr[3]), .O(n372) );
  OR_GATE U487 ( .I1(n445), .I2(MEM_adr[3]), .O(n436) );
  OR_GATE U488 ( .I1(n374), .I2(adr1[4]), .O(n435) );
  INV_GATE U489 ( .I1(MEM_adr[4]), .O(n374) );
  OR_GATE U490 ( .I1(n446), .I2(MEM_adr[4]), .O(n434) );
  AND4_GATE U491 ( .I1(n447), .I2(n448), .I3(n449), .I4(n450), .O(n432) );
  OR_GATE U492 ( .I1(n337), .I2(MEM_adr[5]), .O(n450) );
  OR_GATE U493 ( .I1(n380), .I2(adr1[5]), .O(n449) );
  INV_GATE U494 ( .I1(MEM_adr[5]), .O(n380) );
  OR_GATE U495 ( .I1(n381), .I2(adr1[0]), .O(n448) );
  INV_GATE U496 ( .I1(MEM_adr[0]), .O(n381) );
  OR_GATE U497 ( .I1(n451), .I2(MEM_adr[0]), .O(n447) );
  INV_GATE U498 ( .I1(n346), .O(n339) );
  AND_GATE U499 ( .I1(n429), .I2(n452), .O(n346) );
  OR_GATE U500 ( .I1(n430), .I2(n453), .O(n452) );
  NAND5_GATE U501 ( .I1(n454), .I2(n455), .I3(n456), .I4(n457), .I5(n458), .O(
        n430) );
  AND3_GATE U502 ( .I1(n459), .I2(n460), .I3(EX_ecr), .O(n458) );
  OR_GATE U503 ( .I1(n451), .I2(EX_adr[0]), .O(n460) );
  OR_GATE U504 ( .I1(n392), .I2(adr1[0]), .O(n459) );
  INV_GATE U505 ( .I1(EX_adr[0]), .O(n392) );
  AND4_GATE U506 ( .I1(n461), .I2(n462), .I3(n463), .I4(n464), .O(n457) );
  OR_GATE U507 ( .I1(n443), .I2(EX_adr[1]), .O(n464) );
  OR_GATE U508 ( .I1(n397), .I2(adr1[1]), .O(n463) );
  INV_GATE U509 ( .I1(EX_adr[1]), .O(n397) );
  OR_GATE U510 ( .I1(n444), .I2(EX_adr[2]), .O(n462) );
  OR_GATE U511 ( .I1(n398), .I2(adr1[2]), .O(n461) );
  INV_GATE U512 ( .I1(EX_adr[2]), .O(n398) );
  AND4_GATE U513 ( .I1(n465), .I2(n466), .I3(n467), .I4(n468), .O(n456) );
  OR_GATE U514 ( .I1(n337), .I2(EX_adr[5]), .O(n468) );
  OR_GATE U515 ( .I1(n403), .I2(adr1[5]), .O(n467) );
  INV_GATE U516 ( .I1(EX_adr[5]), .O(n403) );
  OR_GATE U517 ( .I1(n445), .I2(EX_adr[3]), .O(n466) );
  OR_GATE U518 ( .I1(n404), .I2(adr1[3]), .O(n465) );
  INV_GATE U519 ( .I1(EX_adr[3]), .O(n404) );
  OR_GATE U520 ( .I1(n446), .I2(EX_adr[4]), .O(n455) );
  OR_GATE U521 ( .I1(n405), .I2(adr1[4]), .O(n454) );
  INV_GATE U522 ( .I1(EX_adr[4]), .O(n405) );
  NAND5_GATE U523 ( .I1(n431), .I2(DI_ecr), .I3(n469), .I4(n470), .I5(n471), 
        .O(n429) );
  AND4_GATE U524 ( .I1(n472), .I2(n473), .I3(n474), .I4(n475), .O(n471) );
  OR_GATE U525 ( .I1(n444), .I2(DI_adr[2]), .O(n475) );
  OR_GATE U526 ( .I1(n413), .I2(adr1[2]), .O(n474) );
  INV_GATE U527 ( .I1(DI_adr[2]), .O(n413) );
  OR_GATE U528 ( .I1(n445), .I2(DI_adr[3]), .O(n473) );
  OR_GATE U529 ( .I1(n414), .I2(adr1[3]), .O(n472) );
  INV_GATE U530 ( .I1(DI_adr[3]), .O(n414) );
  AND4_GATE U531 ( .I1(n476), .I2(n477), .I3(n478), .I4(n479), .O(n470) );
  OR_GATE U532 ( .I1(n446), .I2(DI_adr[4]), .O(n479) );
  OR_GATE U533 ( .I1(n419), .I2(adr1[4]), .O(n478) );
  INV_GATE U534 ( .I1(DI_adr[4]), .O(n419) );
  OR_GATE U535 ( .I1(n337), .I2(DI_adr[5]), .O(n477) );
  INV_GATE U536 ( .I1(adr1[5]), .O(n337) );
  OR_GATE U537 ( .I1(n420), .I2(adr1[5]), .O(n476) );
  INV_GATE U538 ( .I1(DI_adr[5]), .O(n420) );
  AND4_GATE U539 ( .I1(n480), .I2(n481), .I3(n482), .I4(n483), .O(n469) );
  OR_GATE U540 ( .I1(n451), .I2(DI_adr[0]), .O(n483) );
  OR_GATE U541 ( .I1(n425), .I2(adr1[0]), .O(n482) );
  INV_GATE U542 ( .I1(DI_adr[0]), .O(n425) );
  OR_GATE U543 ( .I1(n443), .I2(DI_adr[1]), .O(n481) );
  OR_GATE U544 ( .I1(n426), .I2(adr1[1]), .O(n480) );
  INV_GATE U545 ( .I1(DI_adr[1]), .O(n426) );
  INV_GATE U546 ( .I1(n453), .O(n431) );
  NAND_GATE U547 ( .I1(use1), .I2(n484), .O(n453) );
  NAND5_GATE U548 ( .I1(n446), .I2(n445), .I3(n444), .I4(n443), .I5(n451), .O(
        n484) );
  INV_GATE U549 ( .I1(adr1[0]), .O(n451) );
  INV_GATE U550 ( .I1(adr1[1]), .O(n443) );
  INV_GATE U551 ( .I1(adr1[2]), .O(n444) );
  INV_GATE U552 ( .I1(adr1[3]), .O(n445) );
  INV_GATE U553 ( .I1(adr1[4]), .O(n446) );
endmodule


module pps_mem ( clock, reset, stop_all, clear, MTC_data, MTC_adr, MTC_r_w, 
        MTC_req, CTM_data, EX_adr, EX_data_ual, EX_adresse, EX_adr_reg_dest, 
        EX_ecr_reg, EX_op_mem, EX_r_w, EX_exc_cause, EX_level, EX_it_ok, 
        MEM_adr, MEM_adr_reg_dest, MEM_ecr_reg, MEM_data_ecr, MEM_exc_cause, 
        MEM_level, MEM_it_ok );
  output [31:0] MTC_data;
  output [31:0] MTC_adr;
  input [31:0] CTM_data;
  input [31:0] EX_adr;
  input [31:0] EX_data_ual;
  input [31:0] EX_adresse;
  input [5:0] EX_adr_reg_dest;
  input [31:0] EX_exc_cause;
  input [1:0] EX_level;
  output [31:0] MEM_adr;
  output [5:0] MEM_adr_reg_dest;
  output [31:0] MEM_data_ecr;
  output [31:0] MEM_exc_cause;
  output [1:0] MEM_level;
  input clock, reset, stop_all, clear, EX_ecr_reg, EX_op_mem, EX_r_w, EX_it_ok;
  output MTC_r_w, MTC_req, MEM_ecr_reg, MEM_it_ok;
  wire   EX_r_w, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n1, n2, n3;
  assign MTC_data[31] = EX_data_ual[31];
  assign MTC_data[30] = EX_data_ual[30];
  assign MTC_data[29] = EX_data_ual[29];
  assign MTC_data[28] = EX_data_ual[28];
  assign MTC_data[27] = EX_data_ual[27];
  assign MTC_data[26] = EX_data_ual[26];
  assign MTC_data[25] = EX_data_ual[25];
  assign MTC_data[24] = EX_data_ual[24];
  assign MTC_data[23] = EX_data_ual[23];
  assign MTC_data[22] = EX_data_ual[22];
  assign MTC_data[21] = EX_data_ual[21];
  assign MTC_data[20] = EX_data_ual[20];
  assign MTC_data[19] = EX_data_ual[19];
  assign MTC_data[18] = EX_data_ual[18];
  assign MTC_data[17] = EX_data_ual[17];
  assign MTC_data[16] = EX_data_ual[16];
  assign MTC_data[15] = EX_data_ual[15];
  assign MTC_data[14] = EX_data_ual[14];
  assign MTC_data[13] = EX_data_ual[13];
  assign MTC_data[12] = EX_data_ual[12];
  assign MTC_data[11] = EX_data_ual[11];
  assign MTC_data[10] = EX_data_ual[10];
  assign MTC_data[9] = EX_data_ual[9];
  assign MTC_data[8] = EX_data_ual[8];
  assign MTC_data[7] = EX_data_ual[7];
  assign MTC_data[6] = EX_data_ual[6];
  assign MTC_data[5] = EX_data_ual[5];
  assign MTC_data[4] = EX_data_ual[4];
  assign MTC_data[3] = EX_data_ual[3];
  assign MTC_data[2] = EX_data_ual[2];
  assign MTC_data[1] = EX_data_ual[1];
  assign MTC_data[0] = EX_data_ual[0];
  assign MTC_adr[31] = EX_adresse[31];
  assign MTC_adr[30] = EX_adresse[30];
  assign MTC_adr[29] = EX_adresse[29];
  assign MTC_adr[28] = EX_adresse[28];
  assign MTC_adr[27] = EX_adresse[27];
  assign MTC_adr[26] = EX_adresse[26];
  assign MTC_adr[25] = EX_adresse[25];
  assign MTC_adr[24] = EX_adresse[24];
  assign MTC_adr[23] = EX_adresse[23];
  assign MTC_adr[22] = EX_adresse[22];
  assign MTC_adr[21] = EX_adresse[21];
  assign MTC_adr[20] = EX_adresse[20];
  assign MTC_adr[19] = EX_adresse[19];
  assign MTC_adr[18] = EX_adresse[18];
  assign MTC_adr[17] = EX_adresse[17];
  assign MTC_adr[16] = EX_adresse[16];
  assign MTC_adr[15] = EX_adresse[15];
  assign MTC_adr[14] = EX_adresse[14];
  assign MTC_adr[13] = EX_adresse[13];
  assign MTC_adr[12] = EX_adresse[12];
  assign MTC_adr[11] = EX_adresse[11];
  assign MTC_adr[10] = EX_adresse[10];
  assign MTC_adr[9] = EX_adresse[9];
  assign MTC_adr[8] = EX_adresse[8];
  assign MTC_adr[7] = EX_adresse[7];
  assign MTC_adr[6] = EX_adresse[6];
  assign MTC_adr[5] = EX_adresse[5];
  assign MTC_adr[4] = EX_adresse[4];
  assign MTC_adr[3] = EX_adresse[3];
  assign MTC_adr[2] = EX_adresse[2];
  assign MTC_adr[1] = EX_adresse[1];
  assign MTC_adr[0] = EX_adresse[0];
  assign MTC_r_w = EX_r_w;

  FLIP_FLOP_D MEM_it_ok_reg ( .D(n362), .CK(clock), .Q(MEM_it_ok) );
  FLIP_FLOP_D \MEM_adr_reg[31]  ( .D(n361), .CK(clock), .Q(MEM_adr[31]) );
  FLIP_FLOP_D \MEM_adr_reg[30]  ( .D(n360), .CK(clock), .Q(MEM_adr[30]) );
  FLIP_FLOP_D \MEM_adr_reg[29]  ( .D(n359), .CK(clock), .Q(MEM_adr[29]) );
  FLIP_FLOP_D \MEM_adr_reg[28]  ( .D(n358), .CK(clock), .Q(MEM_adr[28]) );
  FLIP_FLOP_D \MEM_adr_reg[27]  ( .D(n357), .CK(clock), .Q(MEM_adr[27]) );
  FLIP_FLOP_D \MEM_adr_reg[26]  ( .D(n356), .CK(clock), .Q(MEM_adr[26]) );
  FLIP_FLOP_D \MEM_adr_reg[25]  ( .D(n355), .CK(clock), .Q(MEM_adr[25]) );
  FLIP_FLOP_D \MEM_adr_reg[24]  ( .D(n354), .CK(clock), .Q(MEM_adr[24]) );
  FLIP_FLOP_D \MEM_adr_reg[23]  ( .D(n353), .CK(clock), .Q(MEM_adr[23]) );
  FLIP_FLOP_D \MEM_adr_reg[22]  ( .D(n352), .CK(clock), .Q(MEM_adr[22]) );
  FLIP_FLOP_D \MEM_adr_reg[21]  ( .D(n351), .CK(clock), .Q(MEM_adr[21]) );
  FLIP_FLOP_D \MEM_adr_reg[20]  ( .D(n350), .CK(clock), .Q(MEM_adr[20]) );
  FLIP_FLOP_D \MEM_adr_reg[19]  ( .D(n349), .CK(clock), .Q(MEM_adr[19]) );
  FLIP_FLOP_D \MEM_adr_reg[18]  ( .D(n348), .CK(clock), .Q(MEM_adr[18]) );
  FLIP_FLOP_D \MEM_adr_reg[17]  ( .D(n347), .CK(clock), .Q(MEM_adr[17]) );
  FLIP_FLOP_D \MEM_adr_reg[16]  ( .D(n346), .CK(clock), .Q(MEM_adr[16]) );
  FLIP_FLOP_D \MEM_adr_reg[15]  ( .D(n345), .CK(clock), .Q(MEM_adr[15]) );
  FLIP_FLOP_D \MEM_adr_reg[14]  ( .D(n344), .CK(clock), .Q(MEM_adr[14]) );
  FLIP_FLOP_D \MEM_adr_reg[13]  ( .D(n343), .CK(clock), .Q(MEM_adr[13]) );
  FLIP_FLOP_D \MEM_adr_reg[12]  ( .D(n342), .CK(clock), .Q(MEM_adr[12]) );
  FLIP_FLOP_D \MEM_adr_reg[11]  ( .D(n341), .CK(clock), .Q(MEM_adr[11]) );
  FLIP_FLOP_D \MEM_adr_reg[10]  ( .D(n340), .CK(clock), .Q(MEM_adr[10]) );
  FLIP_FLOP_D \MEM_adr_reg[9]  ( .D(n339), .CK(clock), .Q(MEM_adr[9]) );
  FLIP_FLOP_D \MEM_adr_reg[8]  ( .D(n338), .CK(clock), .Q(MEM_adr[8]) );
  FLIP_FLOP_D \MEM_adr_reg[7]  ( .D(n337), .CK(clock), .Q(MEM_adr[7]) );
  FLIP_FLOP_D \MEM_adr_reg[6]  ( .D(n336), .CK(clock), .Q(MEM_adr[6]) );
  FLIP_FLOP_D \MEM_adr_reg[5]  ( .D(n335), .CK(clock), .Q(MEM_adr[5]) );
  FLIP_FLOP_D \MEM_adr_reg[4]  ( .D(n334), .CK(clock), .Q(MEM_adr[4]) );
  FLIP_FLOP_D \MEM_adr_reg[3]  ( .D(n333), .CK(clock), .Q(MEM_adr[3]) );
  FLIP_FLOP_D \MEM_adr_reg[2]  ( .D(n332), .CK(clock), .Q(MEM_adr[2]) );
  FLIP_FLOP_D \MEM_adr_reg[1]  ( .D(n331), .CK(clock), .Q(MEM_adr[1]) );
  FLIP_FLOP_D \MEM_adr_reg[0]  ( .D(n330), .CK(clock), .Q(MEM_adr[0]) );
  FLIP_FLOP_D \MEM_adr_reg_dest_reg[5]  ( .D(n329), .CK(clock), .Q(
        MEM_adr_reg_dest[5]) );
  FLIP_FLOP_D \MEM_adr_reg_dest_reg[4]  ( .D(n328), .CK(clock), .Q(
        MEM_adr_reg_dest[4]) );
  FLIP_FLOP_D \MEM_adr_reg_dest_reg[3]  ( .D(n327), .CK(clock), .Q(
        MEM_adr_reg_dest[3]) );
  FLIP_FLOP_D \MEM_adr_reg_dest_reg[2]  ( .D(n326), .CK(clock), .Q(
        MEM_adr_reg_dest[2]) );
  FLIP_FLOP_D \MEM_adr_reg_dest_reg[1]  ( .D(n325), .CK(clock), .Q(
        MEM_adr_reg_dest[1]) );
  FLIP_FLOP_D \MEM_adr_reg_dest_reg[0]  ( .D(n324), .CK(clock), .Q(
        MEM_adr_reg_dest[0]) );
  FLIP_FLOP_D MEM_ecr_reg_reg ( .D(n323), .CK(clock), .Q(MEM_ecr_reg) );
  FLIP_FLOP_D \MEM_data_ecr_reg[31]  ( .D(n322), .CK(clock), .Q(
        MEM_data_ecr[31]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[30]  ( .D(n321), .CK(clock), .Q(
        MEM_data_ecr[30]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[29]  ( .D(n320), .CK(clock), .Q(
        MEM_data_ecr[29]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[28]  ( .D(n319), .CK(clock), .Q(
        MEM_data_ecr[28]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[27]  ( .D(n318), .CK(clock), .Q(
        MEM_data_ecr[27]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[26]  ( .D(n317), .CK(clock), .Q(
        MEM_data_ecr[26]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[25]  ( .D(n316), .CK(clock), .Q(
        MEM_data_ecr[25]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[24]  ( .D(n315), .CK(clock), .Q(
        MEM_data_ecr[24]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[23]  ( .D(n314), .CK(clock), .Q(
        MEM_data_ecr[23]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[22]  ( .D(n313), .CK(clock), .Q(
        MEM_data_ecr[22]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[21]  ( .D(n312), .CK(clock), .Q(
        MEM_data_ecr[21]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[20]  ( .D(n311), .CK(clock), .Q(
        MEM_data_ecr[20]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[19]  ( .D(n310), .CK(clock), .Q(
        MEM_data_ecr[19]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[18]  ( .D(n309), .CK(clock), .Q(
        MEM_data_ecr[18]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[17]  ( .D(n308), .CK(clock), .Q(
        MEM_data_ecr[17]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[16]  ( .D(n307), .CK(clock), .Q(
        MEM_data_ecr[16]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[15]  ( .D(n306), .CK(clock), .Q(
        MEM_data_ecr[15]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[14]  ( .D(n305), .CK(clock), .Q(
        MEM_data_ecr[14]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[13]  ( .D(n304), .CK(clock), .Q(
        MEM_data_ecr[13]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[12]  ( .D(n303), .CK(clock), .Q(
        MEM_data_ecr[12]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[11]  ( .D(n302), .CK(clock), .Q(
        MEM_data_ecr[11]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[10]  ( .D(n301), .CK(clock), .Q(
        MEM_data_ecr[10]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[9]  ( .D(n300), .CK(clock), .Q(MEM_data_ecr[9]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[8]  ( .D(n299), .CK(clock), .Q(MEM_data_ecr[8]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[7]  ( .D(n298), .CK(clock), .Q(MEM_data_ecr[7]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[6]  ( .D(n297), .CK(clock), .Q(MEM_data_ecr[6]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[5]  ( .D(n296), .CK(clock), .Q(MEM_data_ecr[5]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[4]  ( .D(n295), .CK(clock), .Q(MEM_data_ecr[4]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[3]  ( .D(n294), .CK(clock), .Q(MEM_data_ecr[3]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[2]  ( .D(n293), .CK(clock), .Q(MEM_data_ecr[2]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[1]  ( .D(n292), .CK(clock), .Q(MEM_data_ecr[1]) );
  FLIP_FLOP_D \MEM_data_ecr_reg[0]  ( .D(n291), .CK(clock), .Q(MEM_data_ecr[0]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[31]  ( .D(n290), .CK(clock), .Q(
        MEM_exc_cause[31]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[30]  ( .D(n289), .CK(clock), .Q(
        MEM_exc_cause[30]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[29]  ( .D(n288), .CK(clock), .Q(
        MEM_exc_cause[29]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[28]  ( .D(n287), .CK(clock), .Q(
        MEM_exc_cause[28]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[27]  ( .D(n286), .CK(clock), .Q(
        MEM_exc_cause[27]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[26]  ( .D(n285), .CK(clock), .Q(
        MEM_exc_cause[26]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[25]  ( .D(n284), .CK(clock), .Q(
        MEM_exc_cause[25]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[24]  ( .D(n283), .CK(clock), .Q(
        MEM_exc_cause[24]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[23]  ( .D(n282), .CK(clock), .Q(
        MEM_exc_cause[23]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[22]  ( .D(n281), .CK(clock), .Q(
        MEM_exc_cause[22]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[21]  ( .D(n280), .CK(clock), .Q(
        MEM_exc_cause[21]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[20]  ( .D(n279), .CK(clock), .Q(
        MEM_exc_cause[20]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[19]  ( .D(n278), .CK(clock), .Q(
        MEM_exc_cause[19]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[18]  ( .D(n277), .CK(clock), .Q(
        MEM_exc_cause[18]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[17]  ( .D(n276), .CK(clock), .Q(
        MEM_exc_cause[17]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[16]  ( .D(n275), .CK(clock), .Q(
        MEM_exc_cause[16]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[15]  ( .D(n274), .CK(clock), .Q(
        MEM_exc_cause[15]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[14]  ( .D(n273), .CK(clock), .Q(
        MEM_exc_cause[14]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[13]  ( .D(n272), .CK(clock), .Q(
        MEM_exc_cause[13]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[12]  ( .D(n271), .CK(clock), .Q(
        MEM_exc_cause[12]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[11]  ( .D(n270), .CK(clock), .Q(
        MEM_exc_cause[11]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[10]  ( .D(n269), .CK(clock), .Q(
        MEM_exc_cause[10]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[9]  ( .D(n268), .CK(clock), .Q(
        MEM_exc_cause[9]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[8]  ( .D(n267), .CK(clock), .Q(
        MEM_exc_cause[8]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[7]  ( .D(n266), .CK(clock), .Q(
        MEM_exc_cause[7]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[6]  ( .D(n265), .CK(clock), .Q(
        MEM_exc_cause[6]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[5]  ( .D(n264), .CK(clock), .Q(
        MEM_exc_cause[5]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[4]  ( .D(n263), .CK(clock), .Q(
        MEM_exc_cause[4]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[3]  ( .D(n262), .CK(clock), .Q(
        MEM_exc_cause[3]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[2]  ( .D(n261), .CK(clock), .Q(
        MEM_exc_cause[2]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[1]  ( .D(n260), .CK(clock), .Q(
        MEM_exc_cause[1]) );
  FLIP_FLOP_D \MEM_exc_cause_reg[0]  ( .D(n259), .CK(clock), .Q(
        MEM_exc_cause[0]) );
  FLIP_FLOP_D \MEM_level_reg[1]  ( .D(n258), .CK(clock), .Q(MEM_level[1]) );
  FLIP_FLOP_D \MEM_level_reg[0]  ( .D(n257), .CK(clock), .Q(MEM_level[0]) );
  NAND_GATE U6 ( .I1(n5), .I2(n6), .O(n257) );
  NAND_GATE U7 ( .I1(n7), .I2(n8), .O(n6) );
  OR_GATE U8 ( .I1(EX_level[0]), .I2(n9), .O(n7) );
  NAND_GATE U9 ( .I1(MEM_level[0]), .I2(n2), .O(n5) );
  NAND_GATE U10 ( .I1(n10), .I2(n11), .O(n258) );
  NAND_GATE U11 ( .I1(n12), .I2(n8), .O(n11) );
  OR_GATE U12 ( .I1(EX_level[1]), .I2(n9), .O(n12) );
  NAND_GATE U13 ( .I1(MEM_level[1]), .I2(n2), .O(n10) );
  NAND_GATE U14 ( .I1(n13), .I2(n14), .O(n259) );
  NAND_GATE U15 ( .I1(EX_exc_cause[0]), .I2(n15), .O(n14) );
  NAND_GATE U16 ( .I1(MEM_exc_cause[0]), .I2(n2), .O(n13) );
  NAND_GATE U17 ( .I1(n16), .I2(n17), .O(n260) );
  NAND_GATE U18 ( .I1(EX_exc_cause[1]), .I2(n15), .O(n17) );
  NAND_GATE U19 ( .I1(MEM_exc_cause[1]), .I2(n2), .O(n16) );
  NAND_GATE U20 ( .I1(n18), .I2(n19), .O(n261) );
  NAND_GATE U21 ( .I1(EX_exc_cause[2]), .I2(n15), .O(n19) );
  NAND_GATE U22 ( .I1(MEM_exc_cause[2]), .I2(n2), .O(n18) );
  NAND_GATE U23 ( .I1(n20), .I2(n21), .O(n262) );
  NAND_GATE U24 ( .I1(EX_exc_cause[3]), .I2(n15), .O(n21) );
  NAND_GATE U25 ( .I1(MEM_exc_cause[3]), .I2(n2), .O(n20) );
  NAND_GATE U26 ( .I1(n22), .I2(n23), .O(n263) );
  NAND_GATE U27 ( .I1(EX_exc_cause[4]), .I2(n15), .O(n23) );
  NAND_GATE U28 ( .I1(MEM_exc_cause[4]), .I2(n2), .O(n22) );
  NAND_GATE U29 ( .I1(n24), .I2(n25), .O(n264) );
  NAND_GATE U30 ( .I1(EX_exc_cause[5]), .I2(n15), .O(n25) );
  NAND_GATE U31 ( .I1(MEM_exc_cause[5]), .I2(n2), .O(n24) );
  NAND_GATE U32 ( .I1(n26), .I2(n27), .O(n265) );
  NAND_GATE U33 ( .I1(EX_exc_cause[6]), .I2(n15), .O(n27) );
  NAND_GATE U34 ( .I1(MEM_exc_cause[6]), .I2(n2), .O(n26) );
  NAND_GATE U35 ( .I1(n28), .I2(n29), .O(n266) );
  NAND_GATE U36 ( .I1(EX_exc_cause[7]), .I2(n15), .O(n29) );
  NAND_GATE U37 ( .I1(MEM_exc_cause[7]), .I2(n2), .O(n28) );
  NAND_GATE U38 ( .I1(n30), .I2(n31), .O(n267) );
  NAND_GATE U39 ( .I1(EX_exc_cause[8]), .I2(n15), .O(n31) );
  NAND_GATE U40 ( .I1(MEM_exc_cause[8]), .I2(n2), .O(n30) );
  NAND_GATE U41 ( .I1(n32), .I2(n33), .O(n268) );
  NAND_GATE U42 ( .I1(EX_exc_cause[9]), .I2(n15), .O(n33) );
  NAND_GATE U43 ( .I1(MEM_exc_cause[9]), .I2(n2), .O(n32) );
  NAND_GATE U44 ( .I1(n34), .I2(n35), .O(n269) );
  NAND_GATE U45 ( .I1(EX_exc_cause[10]), .I2(n15), .O(n35) );
  NAND_GATE U46 ( .I1(MEM_exc_cause[10]), .I2(n2), .O(n34) );
  NAND_GATE U47 ( .I1(n36), .I2(n37), .O(n270) );
  NAND_GATE U48 ( .I1(EX_exc_cause[11]), .I2(n15), .O(n37) );
  NAND_GATE U49 ( .I1(MEM_exc_cause[11]), .I2(n2), .O(n36) );
  NAND_GATE U50 ( .I1(n38), .I2(n39), .O(n271) );
  NAND_GATE U51 ( .I1(EX_exc_cause[12]), .I2(n15), .O(n39) );
  NAND_GATE U52 ( .I1(MEM_exc_cause[12]), .I2(n2), .O(n38) );
  NAND_GATE U53 ( .I1(n40), .I2(n41), .O(n272) );
  NAND_GATE U54 ( .I1(EX_exc_cause[13]), .I2(n15), .O(n41) );
  NAND_GATE U55 ( .I1(MEM_exc_cause[13]), .I2(n2), .O(n40) );
  NAND_GATE U56 ( .I1(n42), .I2(n43), .O(n273) );
  NAND_GATE U57 ( .I1(EX_exc_cause[14]), .I2(n15), .O(n43) );
  NAND_GATE U58 ( .I1(MEM_exc_cause[14]), .I2(n2), .O(n42) );
  NAND_GATE U59 ( .I1(n44), .I2(n45), .O(n274) );
  NAND_GATE U60 ( .I1(EX_exc_cause[15]), .I2(n15), .O(n45) );
  NAND_GATE U61 ( .I1(MEM_exc_cause[15]), .I2(n2), .O(n44) );
  NAND_GATE U62 ( .I1(n46), .I2(n47), .O(n275) );
  NAND_GATE U63 ( .I1(EX_exc_cause[16]), .I2(n15), .O(n47) );
  NAND_GATE U64 ( .I1(MEM_exc_cause[16]), .I2(n2), .O(n46) );
  NAND_GATE U65 ( .I1(n48), .I2(n49), .O(n276) );
  NAND_GATE U66 ( .I1(EX_exc_cause[17]), .I2(n15), .O(n49) );
  NAND_GATE U67 ( .I1(MEM_exc_cause[17]), .I2(n2), .O(n48) );
  NAND_GATE U68 ( .I1(n50), .I2(n51), .O(n277) );
  NAND_GATE U69 ( .I1(EX_exc_cause[18]), .I2(n15), .O(n51) );
  NAND_GATE U70 ( .I1(MEM_exc_cause[18]), .I2(n2), .O(n50) );
  NAND_GATE U71 ( .I1(n52), .I2(n53), .O(n278) );
  NAND_GATE U72 ( .I1(EX_exc_cause[19]), .I2(n15), .O(n53) );
  NAND_GATE U73 ( .I1(MEM_exc_cause[19]), .I2(n2), .O(n52) );
  NAND_GATE U74 ( .I1(n54), .I2(n55), .O(n279) );
  NAND_GATE U75 ( .I1(EX_exc_cause[20]), .I2(n15), .O(n55) );
  NAND_GATE U76 ( .I1(MEM_exc_cause[20]), .I2(n2), .O(n54) );
  NAND_GATE U77 ( .I1(n56), .I2(n57), .O(n280) );
  NAND_GATE U78 ( .I1(EX_exc_cause[21]), .I2(n15), .O(n57) );
  NAND_GATE U79 ( .I1(MEM_exc_cause[21]), .I2(n2), .O(n56) );
  NAND_GATE U80 ( .I1(n58), .I2(n59), .O(n281) );
  NAND_GATE U81 ( .I1(EX_exc_cause[22]), .I2(n15), .O(n59) );
  NAND_GATE U82 ( .I1(MEM_exc_cause[22]), .I2(n2), .O(n58) );
  NAND_GATE U83 ( .I1(n60), .I2(n61), .O(n282) );
  NAND_GATE U84 ( .I1(EX_exc_cause[23]), .I2(n15), .O(n61) );
  NAND_GATE U85 ( .I1(MEM_exc_cause[23]), .I2(n2), .O(n60) );
  NAND_GATE U86 ( .I1(n62), .I2(n63), .O(n283) );
  NAND_GATE U87 ( .I1(EX_exc_cause[24]), .I2(n15), .O(n63) );
  NAND_GATE U88 ( .I1(MEM_exc_cause[24]), .I2(n2), .O(n62) );
  NAND_GATE U89 ( .I1(n64), .I2(n65), .O(n284) );
  NAND_GATE U90 ( .I1(EX_exc_cause[25]), .I2(n15), .O(n65) );
  NAND_GATE U91 ( .I1(MEM_exc_cause[25]), .I2(n2), .O(n64) );
  NAND_GATE U92 ( .I1(n66), .I2(n67), .O(n285) );
  NAND_GATE U93 ( .I1(EX_exc_cause[26]), .I2(n15), .O(n67) );
  NAND_GATE U94 ( .I1(MEM_exc_cause[26]), .I2(n2), .O(n66) );
  NAND_GATE U95 ( .I1(n68), .I2(n69), .O(n286) );
  NAND_GATE U96 ( .I1(EX_exc_cause[27]), .I2(n15), .O(n69) );
  NAND_GATE U97 ( .I1(MEM_exc_cause[27]), .I2(n2), .O(n68) );
  NAND_GATE U98 ( .I1(n70), .I2(n71), .O(n287) );
  NAND_GATE U99 ( .I1(EX_exc_cause[28]), .I2(n15), .O(n71) );
  NAND_GATE U100 ( .I1(MEM_exc_cause[28]), .I2(n2), .O(n70) );
  NAND_GATE U101 ( .I1(n72), .I2(n73), .O(n288) );
  NAND_GATE U102 ( .I1(EX_exc_cause[29]), .I2(n15), .O(n73) );
  NAND_GATE U103 ( .I1(MEM_exc_cause[29]), .I2(n2), .O(n72) );
  NAND_GATE U104 ( .I1(n74), .I2(n75), .O(n289) );
  NAND_GATE U105 ( .I1(EX_exc_cause[30]), .I2(n15), .O(n75) );
  NAND_GATE U106 ( .I1(MEM_exc_cause[30]), .I2(n2), .O(n74) );
  NAND_GATE U107 ( .I1(n76), .I2(n77), .O(n290) );
  NAND_GATE U108 ( .I1(EX_exc_cause[31]), .I2(n15), .O(n77) );
  NAND_GATE U109 ( .I1(MEM_exc_cause[31]), .I2(n2), .O(n76) );
  NAND3_GATE U110 ( .I1(n78), .I2(n79), .I3(n80), .O(n291) );
  NAND_GATE U111 ( .I1(MEM_data_ecr[0]), .I2(n2), .O(n80) );
  NAND_GATE U112 ( .I1(CTM_data[0]), .I2(n81), .O(n79) );
  NAND_GATE U113 ( .I1(EX_data_ual[0]), .I2(n82), .O(n78) );
  NAND3_GATE U114 ( .I1(n83), .I2(n84), .I3(n85), .O(n292) );
  NAND_GATE U115 ( .I1(MEM_data_ecr[1]), .I2(n2), .O(n85) );
  NAND_GATE U116 ( .I1(CTM_data[1]), .I2(n81), .O(n84) );
  NAND_GATE U117 ( .I1(EX_data_ual[1]), .I2(n82), .O(n83) );
  NAND3_GATE U118 ( .I1(n86), .I2(n87), .I3(n88), .O(n293) );
  NAND_GATE U119 ( .I1(MEM_data_ecr[2]), .I2(n2), .O(n88) );
  NAND_GATE U120 ( .I1(CTM_data[2]), .I2(n81), .O(n87) );
  NAND_GATE U121 ( .I1(EX_data_ual[2]), .I2(n82), .O(n86) );
  NAND3_GATE U122 ( .I1(n89), .I2(n90), .I3(n91), .O(n294) );
  NAND_GATE U123 ( .I1(MEM_data_ecr[3]), .I2(n2), .O(n91) );
  NAND_GATE U124 ( .I1(CTM_data[3]), .I2(n81), .O(n90) );
  NAND_GATE U125 ( .I1(EX_data_ual[3]), .I2(n82), .O(n89) );
  NAND3_GATE U126 ( .I1(n92), .I2(n93), .I3(n94), .O(n295) );
  NAND_GATE U127 ( .I1(MEM_data_ecr[4]), .I2(n2), .O(n94) );
  NAND_GATE U128 ( .I1(CTM_data[4]), .I2(n81), .O(n93) );
  NAND_GATE U129 ( .I1(EX_data_ual[4]), .I2(n82), .O(n92) );
  NAND3_GATE U130 ( .I1(n95), .I2(n96), .I3(n97), .O(n296) );
  NAND_GATE U131 ( .I1(MEM_data_ecr[5]), .I2(n2), .O(n97) );
  NAND_GATE U132 ( .I1(CTM_data[5]), .I2(n81), .O(n96) );
  NAND_GATE U133 ( .I1(EX_data_ual[5]), .I2(n82), .O(n95) );
  NAND3_GATE U134 ( .I1(n98), .I2(n99), .I3(n100), .O(n297) );
  NAND_GATE U135 ( .I1(MEM_data_ecr[6]), .I2(n2), .O(n100) );
  NAND_GATE U136 ( .I1(CTM_data[6]), .I2(n81), .O(n99) );
  NAND_GATE U137 ( .I1(EX_data_ual[6]), .I2(n82), .O(n98) );
  NAND3_GATE U138 ( .I1(n101), .I2(n102), .I3(n103), .O(n298) );
  NAND_GATE U139 ( .I1(MEM_data_ecr[7]), .I2(n2), .O(n103) );
  NAND_GATE U140 ( .I1(CTM_data[7]), .I2(n81), .O(n102) );
  NAND_GATE U141 ( .I1(EX_data_ual[7]), .I2(n82), .O(n101) );
  NAND3_GATE U142 ( .I1(n104), .I2(n105), .I3(n106), .O(n299) );
  NAND_GATE U143 ( .I1(MEM_data_ecr[8]), .I2(n2), .O(n106) );
  NAND_GATE U144 ( .I1(CTM_data[8]), .I2(n81), .O(n105) );
  NAND_GATE U145 ( .I1(EX_data_ual[8]), .I2(n82), .O(n104) );
  NAND3_GATE U146 ( .I1(n107), .I2(n108), .I3(n109), .O(n300) );
  NAND_GATE U147 ( .I1(MEM_data_ecr[9]), .I2(n2), .O(n109) );
  NAND_GATE U148 ( .I1(CTM_data[9]), .I2(n81), .O(n108) );
  NAND_GATE U149 ( .I1(EX_data_ual[9]), .I2(n82), .O(n107) );
  NAND3_GATE U150 ( .I1(n110), .I2(n111), .I3(n112), .O(n301) );
  NAND_GATE U151 ( .I1(MEM_data_ecr[10]), .I2(n2), .O(n112) );
  NAND_GATE U152 ( .I1(CTM_data[10]), .I2(n81), .O(n111) );
  NAND_GATE U153 ( .I1(EX_data_ual[10]), .I2(n82), .O(n110) );
  NAND3_GATE U154 ( .I1(n113), .I2(n114), .I3(n115), .O(n302) );
  NAND_GATE U155 ( .I1(MEM_data_ecr[11]), .I2(n2), .O(n115) );
  NAND_GATE U156 ( .I1(CTM_data[11]), .I2(n81), .O(n114) );
  NAND_GATE U157 ( .I1(EX_data_ual[11]), .I2(n82), .O(n113) );
  NAND3_GATE U158 ( .I1(n116), .I2(n117), .I3(n118), .O(n303) );
  NAND_GATE U159 ( .I1(MEM_data_ecr[12]), .I2(n2), .O(n118) );
  NAND_GATE U160 ( .I1(CTM_data[12]), .I2(n81), .O(n117) );
  NAND_GATE U161 ( .I1(EX_data_ual[12]), .I2(n82), .O(n116) );
  NAND3_GATE U162 ( .I1(n119), .I2(n120), .I3(n121), .O(n304) );
  NAND_GATE U163 ( .I1(MEM_data_ecr[13]), .I2(n2), .O(n121) );
  NAND_GATE U164 ( .I1(CTM_data[13]), .I2(n81), .O(n120) );
  NAND_GATE U165 ( .I1(EX_data_ual[13]), .I2(n82), .O(n119) );
  NAND3_GATE U166 ( .I1(n122), .I2(n123), .I3(n124), .O(n305) );
  NAND_GATE U167 ( .I1(MEM_data_ecr[14]), .I2(n2), .O(n124) );
  NAND_GATE U168 ( .I1(CTM_data[14]), .I2(n81), .O(n123) );
  NAND_GATE U169 ( .I1(EX_data_ual[14]), .I2(n82), .O(n122) );
  NAND3_GATE U170 ( .I1(n125), .I2(n126), .I3(n127), .O(n306) );
  NAND_GATE U171 ( .I1(MEM_data_ecr[15]), .I2(n2), .O(n127) );
  NAND_GATE U172 ( .I1(CTM_data[15]), .I2(n81), .O(n126) );
  NAND_GATE U173 ( .I1(EX_data_ual[15]), .I2(n82), .O(n125) );
  NAND3_GATE U174 ( .I1(n128), .I2(n129), .I3(n130), .O(n307) );
  NAND_GATE U175 ( .I1(MEM_data_ecr[16]), .I2(n2), .O(n130) );
  NAND_GATE U176 ( .I1(CTM_data[16]), .I2(n81), .O(n129) );
  NAND_GATE U177 ( .I1(EX_data_ual[16]), .I2(n82), .O(n128) );
  NAND3_GATE U178 ( .I1(n131), .I2(n132), .I3(n133), .O(n308) );
  NAND_GATE U179 ( .I1(MEM_data_ecr[17]), .I2(n2), .O(n133) );
  NAND_GATE U180 ( .I1(CTM_data[17]), .I2(n81), .O(n132) );
  NAND_GATE U181 ( .I1(EX_data_ual[17]), .I2(n82), .O(n131) );
  NAND3_GATE U182 ( .I1(n134), .I2(n135), .I3(n136), .O(n309) );
  NAND_GATE U183 ( .I1(MEM_data_ecr[18]), .I2(n2), .O(n136) );
  NAND_GATE U184 ( .I1(CTM_data[18]), .I2(n81), .O(n135) );
  NAND_GATE U185 ( .I1(EX_data_ual[18]), .I2(n82), .O(n134) );
  NAND3_GATE U186 ( .I1(n137), .I2(n138), .I3(n139), .O(n310) );
  NAND_GATE U187 ( .I1(MEM_data_ecr[19]), .I2(n2), .O(n139) );
  NAND_GATE U188 ( .I1(CTM_data[19]), .I2(n81), .O(n138) );
  NAND_GATE U189 ( .I1(EX_data_ual[19]), .I2(n82), .O(n137) );
  NAND3_GATE U190 ( .I1(n140), .I2(n141), .I3(n142), .O(n311) );
  NAND_GATE U191 ( .I1(MEM_data_ecr[20]), .I2(n2), .O(n142) );
  NAND_GATE U192 ( .I1(CTM_data[20]), .I2(n81), .O(n141) );
  NAND_GATE U193 ( .I1(EX_data_ual[20]), .I2(n82), .O(n140) );
  NAND3_GATE U194 ( .I1(n143), .I2(n144), .I3(n145), .O(n312) );
  NAND_GATE U195 ( .I1(MEM_data_ecr[21]), .I2(n2), .O(n145) );
  NAND_GATE U196 ( .I1(CTM_data[21]), .I2(n81), .O(n144) );
  NAND_GATE U197 ( .I1(EX_data_ual[21]), .I2(n82), .O(n143) );
  NAND3_GATE U198 ( .I1(n146), .I2(n147), .I3(n148), .O(n313) );
  NAND_GATE U199 ( .I1(MEM_data_ecr[22]), .I2(n2), .O(n148) );
  NAND_GATE U200 ( .I1(CTM_data[22]), .I2(n81), .O(n147) );
  NAND_GATE U201 ( .I1(EX_data_ual[22]), .I2(n82), .O(n146) );
  NAND3_GATE U202 ( .I1(n149), .I2(n150), .I3(n151), .O(n314) );
  NAND_GATE U203 ( .I1(MEM_data_ecr[23]), .I2(n2), .O(n151) );
  NAND_GATE U204 ( .I1(CTM_data[23]), .I2(n81), .O(n150) );
  NAND_GATE U205 ( .I1(EX_data_ual[23]), .I2(n82), .O(n149) );
  NAND3_GATE U206 ( .I1(n152), .I2(n153), .I3(n154), .O(n315) );
  NAND_GATE U207 ( .I1(MEM_data_ecr[24]), .I2(n2), .O(n154) );
  NAND_GATE U208 ( .I1(CTM_data[24]), .I2(n81), .O(n153) );
  NAND_GATE U209 ( .I1(EX_data_ual[24]), .I2(n82), .O(n152) );
  NAND3_GATE U210 ( .I1(n155), .I2(n156), .I3(n157), .O(n316) );
  NAND_GATE U211 ( .I1(MEM_data_ecr[25]), .I2(n2), .O(n157) );
  NAND_GATE U212 ( .I1(CTM_data[25]), .I2(n81), .O(n156) );
  NAND_GATE U213 ( .I1(EX_data_ual[25]), .I2(n82), .O(n155) );
  NAND3_GATE U214 ( .I1(n158), .I2(n159), .I3(n160), .O(n317) );
  NAND_GATE U215 ( .I1(MEM_data_ecr[26]), .I2(n2), .O(n160) );
  NAND_GATE U216 ( .I1(CTM_data[26]), .I2(n81), .O(n159) );
  NAND_GATE U217 ( .I1(EX_data_ual[26]), .I2(n82), .O(n158) );
  NAND3_GATE U218 ( .I1(n161), .I2(n162), .I3(n163), .O(n318) );
  NAND_GATE U219 ( .I1(MEM_data_ecr[27]), .I2(n2), .O(n163) );
  NAND_GATE U220 ( .I1(CTM_data[27]), .I2(n81), .O(n162) );
  NAND_GATE U221 ( .I1(EX_data_ual[27]), .I2(n82), .O(n161) );
  NAND3_GATE U222 ( .I1(n164), .I2(n165), .I3(n166), .O(n319) );
  NAND_GATE U223 ( .I1(MEM_data_ecr[28]), .I2(n2), .O(n166) );
  NAND_GATE U224 ( .I1(CTM_data[28]), .I2(n81), .O(n165) );
  NAND_GATE U225 ( .I1(EX_data_ual[28]), .I2(n82), .O(n164) );
  NAND3_GATE U226 ( .I1(n167), .I2(n168), .I3(n169), .O(n320) );
  NAND_GATE U227 ( .I1(MEM_data_ecr[29]), .I2(n2), .O(n169) );
  NAND_GATE U228 ( .I1(CTM_data[29]), .I2(n81), .O(n168) );
  NAND_GATE U229 ( .I1(EX_data_ual[29]), .I2(n82), .O(n167) );
  NAND3_GATE U230 ( .I1(n170), .I2(n171), .I3(n172), .O(n321) );
  NAND_GATE U231 ( .I1(MEM_data_ecr[30]), .I2(n2), .O(n172) );
  NAND_GATE U232 ( .I1(CTM_data[30]), .I2(n81), .O(n171) );
  NAND_GATE U233 ( .I1(EX_data_ual[30]), .I2(n82), .O(n170) );
  NAND3_GATE U234 ( .I1(n173), .I2(n174), .I3(n175), .O(n322) );
  NAND_GATE U235 ( .I1(MEM_data_ecr[31]), .I2(n2), .O(n175) );
  NAND_GATE U236 ( .I1(CTM_data[31]), .I2(n81), .O(n174) );
  AND3_GATE U237 ( .I1(n8), .I2(n1), .I3(MTC_req), .O(n81) );
  NAND_GATE U238 ( .I1(EX_data_ual[31]), .I2(n82), .O(n173) );
  NOR3_GATE U239 ( .I1(n2), .I2(EX_op_mem), .I3(n9), .O(n82) );
  NAND_GATE U240 ( .I1(n3), .I2(n1), .O(n9) );
  NAND_GATE U241 ( .I1(n176), .I2(n177), .O(n323) );
  NAND_GATE U242 ( .I1(EX_ecr_reg), .I2(n15), .O(n177) );
  NAND_GATE U243 ( .I1(MEM_ecr_reg), .I2(n2), .O(n176) );
  NAND_GATE U244 ( .I1(n178), .I2(n179), .O(n324) );
  NAND_GATE U245 ( .I1(EX_adr_reg_dest[0]), .I2(n15), .O(n179) );
  NAND_GATE U246 ( .I1(MEM_adr_reg_dest[0]), .I2(n2), .O(n178) );
  NAND_GATE U247 ( .I1(n180), .I2(n181), .O(n325) );
  NAND_GATE U248 ( .I1(EX_adr_reg_dest[1]), .I2(n15), .O(n181) );
  NAND_GATE U249 ( .I1(MEM_adr_reg_dest[1]), .I2(n2), .O(n180) );
  NAND_GATE U250 ( .I1(n182), .I2(n183), .O(n326) );
  NAND_GATE U251 ( .I1(EX_adr_reg_dest[2]), .I2(n15), .O(n183) );
  NAND_GATE U252 ( .I1(MEM_adr_reg_dest[2]), .I2(n2), .O(n182) );
  NAND_GATE U253 ( .I1(n184), .I2(n185), .O(n327) );
  NAND_GATE U254 ( .I1(EX_adr_reg_dest[3]), .I2(n15), .O(n185) );
  NAND_GATE U255 ( .I1(MEM_adr_reg_dest[3]), .I2(n2), .O(n184) );
  NAND_GATE U256 ( .I1(n186), .I2(n187), .O(n328) );
  NAND_GATE U257 ( .I1(EX_adr_reg_dest[4]), .I2(n15), .O(n187) );
  NAND_GATE U258 ( .I1(MEM_adr_reg_dest[4]), .I2(n2), .O(n186) );
  NAND_GATE U259 ( .I1(n188), .I2(n189), .O(n329) );
  NAND_GATE U260 ( .I1(EX_adr_reg_dest[5]), .I2(n15), .O(n189) );
  NAND_GATE U261 ( .I1(MEM_adr_reg_dest[5]), .I2(n2), .O(n188) );
  NAND_GATE U262 ( .I1(n190), .I2(n191), .O(n330) );
  NAND_GATE U263 ( .I1(EX_adr[0]), .I2(n192), .O(n191) );
  NAND_GATE U264 ( .I1(MEM_adr[0]), .I2(n2), .O(n190) );
  NAND_GATE U265 ( .I1(n193), .I2(n194), .O(n331) );
  NAND_GATE U266 ( .I1(EX_adr[1]), .I2(n192), .O(n194) );
  NAND_GATE U267 ( .I1(MEM_adr[1]), .I2(n2), .O(n193) );
  NAND_GATE U268 ( .I1(n195), .I2(n196), .O(n332) );
  NAND_GATE U269 ( .I1(EX_adr[2]), .I2(n192), .O(n196) );
  NAND_GATE U270 ( .I1(MEM_adr[2]), .I2(n2), .O(n195) );
  NAND_GATE U271 ( .I1(n197), .I2(n198), .O(n333) );
  NAND_GATE U272 ( .I1(EX_adr[3]), .I2(n192), .O(n198) );
  NAND_GATE U273 ( .I1(MEM_adr[3]), .I2(n2), .O(n197) );
  NAND_GATE U274 ( .I1(n199), .I2(n200), .O(n334) );
  NAND_GATE U275 ( .I1(EX_adr[4]), .I2(n192), .O(n200) );
  NAND_GATE U276 ( .I1(MEM_adr[4]), .I2(n2), .O(n199) );
  NAND_GATE U277 ( .I1(n201), .I2(n202), .O(n335) );
  NAND_GATE U278 ( .I1(EX_adr[5]), .I2(n192), .O(n202) );
  NAND_GATE U279 ( .I1(MEM_adr[5]), .I2(n2), .O(n201) );
  NAND_GATE U280 ( .I1(n203), .I2(n204), .O(n336) );
  NAND_GATE U281 ( .I1(EX_adr[6]), .I2(n192), .O(n204) );
  NAND_GATE U282 ( .I1(MEM_adr[6]), .I2(n2), .O(n203) );
  NAND_GATE U283 ( .I1(n205), .I2(n206), .O(n337) );
  NAND_GATE U284 ( .I1(EX_adr[7]), .I2(n192), .O(n206) );
  NAND_GATE U285 ( .I1(MEM_adr[7]), .I2(n2), .O(n205) );
  NAND_GATE U286 ( .I1(n207), .I2(n208), .O(n338) );
  NAND_GATE U287 ( .I1(EX_adr[8]), .I2(n192), .O(n208) );
  NAND_GATE U288 ( .I1(MEM_adr[8]), .I2(n2), .O(n207) );
  NAND_GATE U289 ( .I1(n209), .I2(n210), .O(n339) );
  NAND_GATE U290 ( .I1(EX_adr[9]), .I2(n192), .O(n210) );
  NAND_GATE U291 ( .I1(MEM_adr[9]), .I2(n2), .O(n209) );
  NAND_GATE U292 ( .I1(n211), .I2(n212), .O(n340) );
  NAND_GATE U293 ( .I1(EX_adr[10]), .I2(n192), .O(n212) );
  NAND_GATE U294 ( .I1(MEM_adr[10]), .I2(n2), .O(n211) );
  NAND_GATE U295 ( .I1(n213), .I2(n214), .O(n341) );
  NAND_GATE U296 ( .I1(EX_adr[11]), .I2(n192), .O(n214) );
  NAND_GATE U297 ( .I1(MEM_adr[11]), .I2(n2), .O(n213) );
  NAND_GATE U298 ( .I1(n215), .I2(n216), .O(n342) );
  NAND_GATE U299 ( .I1(EX_adr[12]), .I2(n192), .O(n216) );
  NAND_GATE U300 ( .I1(MEM_adr[12]), .I2(n2), .O(n215) );
  NAND_GATE U301 ( .I1(n217), .I2(n218), .O(n343) );
  NAND_GATE U302 ( .I1(EX_adr[13]), .I2(n192), .O(n218) );
  NAND_GATE U303 ( .I1(MEM_adr[13]), .I2(n2), .O(n217) );
  NAND_GATE U304 ( .I1(n219), .I2(n220), .O(n344) );
  NAND_GATE U305 ( .I1(EX_adr[14]), .I2(n192), .O(n220) );
  NAND_GATE U306 ( .I1(MEM_adr[14]), .I2(n2), .O(n219) );
  NAND_GATE U307 ( .I1(n221), .I2(n222), .O(n345) );
  NAND_GATE U308 ( .I1(EX_adr[15]), .I2(n192), .O(n222) );
  NAND_GATE U309 ( .I1(MEM_adr[15]), .I2(n2), .O(n221) );
  NAND_GATE U310 ( .I1(n223), .I2(n224), .O(n346) );
  NAND_GATE U311 ( .I1(EX_adr[16]), .I2(n192), .O(n224) );
  NAND_GATE U312 ( .I1(MEM_adr[16]), .I2(n2), .O(n223) );
  NAND_GATE U313 ( .I1(n225), .I2(n226), .O(n347) );
  NAND_GATE U314 ( .I1(EX_adr[17]), .I2(n192), .O(n226) );
  NAND_GATE U315 ( .I1(MEM_adr[17]), .I2(n2), .O(n225) );
  NAND_GATE U316 ( .I1(n227), .I2(n228), .O(n348) );
  NAND_GATE U317 ( .I1(EX_adr[18]), .I2(n192), .O(n228) );
  NAND_GATE U318 ( .I1(MEM_adr[18]), .I2(n2), .O(n227) );
  NAND_GATE U319 ( .I1(n229), .I2(n230), .O(n349) );
  NAND_GATE U320 ( .I1(EX_adr[19]), .I2(n192), .O(n230) );
  NAND_GATE U321 ( .I1(MEM_adr[19]), .I2(n2), .O(n229) );
  NAND_GATE U322 ( .I1(n231), .I2(n232), .O(n350) );
  NAND_GATE U323 ( .I1(EX_adr[20]), .I2(n192), .O(n232) );
  NAND_GATE U324 ( .I1(MEM_adr[20]), .I2(n2), .O(n231) );
  NAND_GATE U325 ( .I1(n233), .I2(n234), .O(n351) );
  NAND_GATE U326 ( .I1(EX_adr[21]), .I2(n192), .O(n234) );
  NAND_GATE U327 ( .I1(MEM_adr[21]), .I2(n2), .O(n233) );
  NAND_GATE U328 ( .I1(n235), .I2(n236), .O(n352) );
  NAND_GATE U329 ( .I1(EX_adr[22]), .I2(n192), .O(n236) );
  NAND_GATE U330 ( .I1(MEM_adr[22]), .I2(n2), .O(n235) );
  NAND_GATE U331 ( .I1(n237), .I2(n238), .O(n353) );
  NAND_GATE U332 ( .I1(EX_adr[23]), .I2(n192), .O(n238) );
  NAND_GATE U333 ( .I1(MEM_adr[23]), .I2(n2), .O(n237) );
  NAND_GATE U334 ( .I1(n239), .I2(n240), .O(n354) );
  NAND_GATE U335 ( .I1(EX_adr[24]), .I2(n192), .O(n240) );
  NAND_GATE U336 ( .I1(MEM_adr[24]), .I2(n2), .O(n239) );
  NAND_GATE U337 ( .I1(n241), .I2(n242), .O(n355) );
  NAND_GATE U338 ( .I1(EX_adr[25]), .I2(n192), .O(n242) );
  NAND_GATE U339 ( .I1(MEM_adr[25]), .I2(n2), .O(n241) );
  NAND_GATE U340 ( .I1(n243), .I2(n244), .O(n356) );
  NAND_GATE U341 ( .I1(EX_adr[26]), .I2(n192), .O(n244) );
  NAND_GATE U342 ( .I1(MEM_adr[26]), .I2(n2), .O(n243) );
  NAND_GATE U343 ( .I1(n245), .I2(n246), .O(n357) );
  NAND_GATE U344 ( .I1(EX_adr[27]), .I2(n192), .O(n246) );
  NAND_GATE U345 ( .I1(MEM_adr[27]), .I2(n2), .O(n245) );
  NAND_GATE U346 ( .I1(n247), .I2(n248), .O(n358) );
  NAND_GATE U347 ( .I1(EX_adr[28]), .I2(n192), .O(n248) );
  NAND_GATE U348 ( .I1(MEM_adr[28]), .I2(n2), .O(n247) );
  NAND_GATE U349 ( .I1(n249), .I2(n250), .O(n359) );
  NAND_GATE U350 ( .I1(EX_adr[29]), .I2(n192), .O(n250) );
  NAND_GATE U351 ( .I1(MEM_adr[29]), .I2(n2), .O(n249) );
  NAND_GATE U352 ( .I1(n251), .I2(n252), .O(n360) );
  NAND_GATE U353 ( .I1(EX_adr[30]), .I2(n192), .O(n252) );
  NAND_GATE U354 ( .I1(MEM_adr[30]), .I2(n2), .O(n251) );
  NAND_GATE U355 ( .I1(n253), .I2(n254), .O(n361) );
  NAND_GATE U356 ( .I1(EX_adr[31]), .I2(n192), .O(n254) );
  NAND_GATE U357 ( .I1(MEM_adr[31]), .I2(n2), .O(n253) );
  NAND_GATE U358 ( .I1(n255), .I2(n256), .O(n362) );
  NAND_GATE U359 ( .I1(EX_it_ok), .I2(n15), .O(n256) );
  AND_GATE U360 ( .I1(n192), .I2(n3), .O(n15) );
  NOR_GATE U361 ( .I1(stop_all), .I2(reset), .O(n192) );
  NAND_GATE U362 ( .I1(MEM_it_ok), .I2(n2), .O(n255) );
  NAND_GATE U363 ( .I1(stop_all), .I2(n1), .O(n8) );
  AND_GATE U364 ( .I1(EX_op_mem), .I2(n3), .O(MTC_req) );
  INV_GATE U3 ( .I1(reset), .O(n1) );
  INV_GATE U4 ( .I1(n8), .O(n2) );
  INV_GATE U5 ( .I1(clear), .O(n3) );
endmodule


module pps_ex ( clock, reset, stop_all, clear, DI_bra, DI_link, DI_op1, DI_op2, 
        DI_code_ual, DI_offset, DI_adr_reg_dest, DI_ecr_reg, DI_mode, 
        DI_op_mem, DI_r_w, DI_adr, DI_exc_cause, DI_level, DI_it_ok, EX_adr, 
        EX_bra_confirm, EX_data_ual, EX_adresse, EX_adr_reg_dest, EX_ecr_reg, 
        EX_op_mem, EX_r_w, EX_exc_cause, EX_level, EX_it_ok );
  input [31:0] DI_op1;
  input [31:0] DI_op2;
  input [27:0] DI_code_ual;
  input [31:0] DI_offset;
  input [5:0] DI_adr_reg_dest;
  input [31:0] DI_adr;
  input [31:0] DI_exc_cause;
  input [1:0] DI_level;
  output [31:0] EX_adr;
  output [31:0] EX_data_ual;
  output [31:0] EX_adresse;
  output [5:0] EX_adr_reg_dest;
  output [31:0] EX_exc_cause;
  output [1:0] EX_level;
  input clock, reset, stop_all, clear, DI_bra, DI_link, DI_ecr_reg, DI_mode,
         DI_op_mem, DI_r_w, DI_it_ok;
  output EX_bra_confirm, EX_ecr_reg, EX_op_mem, EX_r_w, EX_it_ok;
  wire   overflow_ual, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, n14, n15, n16, n17, n19, n20, n21, n22, n23, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n381, n382, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n18,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n101,
         n102, n103, n104, n105, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n380, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n588, n589, n590, n591, n592, n593, n594;
  wire   [31:0] res_ual;
  wire   [31:0] base_adr;

  FLIP_FLOP_D EX_it_ok_reg ( .D(n587), .CK(clock), .Q(EX_it_ok) );
  FLIP_FLOP_D \EX_adr_reg[31]  ( .D(n586), .CK(clock), .Q(EX_adr[31]) );
  FLIP_FLOP_D \EX_adr_reg[30]  ( .D(n585), .CK(clock), .Q(EX_adr[30]) );
  FLIP_FLOP_D \EX_adr_reg[29]  ( .D(n584), .CK(clock), .Q(EX_adr[29]) );
  FLIP_FLOP_D \EX_adr_reg[28]  ( .D(n583), .CK(clock), .Q(EX_adr[28]) );
  FLIP_FLOP_D \EX_adr_reg[27]  ( .D(n582), .CK(clock), .Q(EX_adr[27]) );
  FLIP_FLOP_D \EX_adr_reg[26]  ( .D(n581), .CK(clock), .Q(EX_adr[26]) );
  FLIP_FLOP_D \EX_adr_reg[25]  ( .D(n580), .CK(clock), .Q(EX_adr[25]) );
  FLIP_FLOP_D \EX_adr_reg[24]  ( .D(n579), .CK(clock), .Q(EX_adr[24]) );
  FLIP_FLOP_D \EX_adr_reg[23]  ( .D(n578), .CK(clock), .Q(EX_adr[23]) );
  FLIP_FLOP_D \EX_adr_reg[22]  ( .D(n577), .CK(clock), .Q(EX_adr[22]) );
  FLIP_FLOP_D \EX_adr_reg[21]  ( .D(n576), .CK(clock), .Q(EX_adr[21]) );
  FLIP_FLOP_D \EX_adr_reg[20]  ( .D(n575), .CK(clock), .Q(EX_adr[20]) );
  FLIP_FLOP_D \EX_adr_reg[19]  ( .D(n574), .CK(clock), .Q(EX_adr[19]) );
  FLIP_FLOP_D \EX_adr_reg[18]  ( .D(n573), .CK(clock), .Q(EX_adr[18]) );
  FLIP_FLOP_D \EX_adr_reg[17]  ( .D(n572), .CK(clock), .Q(EX_adr[17]) );
  FLIP_FLOP_D \EX_adr_reg[16]  ( .D(n571), .CK(clock), .Q(EX_adr[16]) );
  FLIP_FLOP_D \EX_adr_reg[15]  ( .D(n570), .CK(clock), .Q(EX_adr[15]) );
  FLIP_FLOP_D \EX_adr_reg[14]  ( .D(n569), .CK(clock), .Q(EX_adr[14]) );
  FLIP_FLOP_D \EX_adr_reg[13]  ( .D(n568), .CK(clock), .Q(EX_adr[13]) );
  FLIP_FLOP_D \EX_adr_reg[12]  ( .D(n567), .CK(clock), .Q(EX_adr[12]) );
  FLIP_FLOP_D \EX_adr_reg[11]  ( .D(n566), .CK(clock), .Q(EX_adr[11]) );
  FLIP_FLOP_D \EX_adr_reg[10]  ( .D(n565), .CK(clock), .Q(EX_adr[10]) );
  FLIP_FLOP_D \EX_adr_reg[9]  ( .D(n564), .CK(clock), .Q(EX_adr[9]) );
  FLIP_FLOP_D \EX_adr_reg[8]  ( .D(n563), .CK(clock), .Q(EX_adr[8]) );
  FLIP_FLOP_D \EX_adr_reg[7]  ( .D(n562), .CK(clock), .Q(EX_adr[7]) );
  FLIP_FLOP_D \EX_adr_reg[6]  ( .D(n561), .CK(clock), .Q(EX_adr[6]) );
  FLIP_FLOP_D \EX_adr_reg[5]  ( .D(n560), .CK(clock), .Q(EX_adr[5]) );
  FLIP_FLOP_D \EX_adr_reg[4]  ( .D(n559), .CK(clock), .Q(EX_adr[4]) );
  FLIP_FLOP_D \EX_adr_reg[3]  ( .D(n558), .CK(clock), .Q(EX_adr[3]) );
  FLIP_FLOP_D \EX_adr_reg[2]  ( .D(n557), .CK(clock), .Q(EX_adr[2]) );
  FLIP_FLOP_D \EX_adr_reg[1]  ( .D(n556), .CK(clock), .Q(EX_adr[1]) );
  FLIP_FLOP_D \EX_adr_reg[0]  ( .D(n555), .CK(clock), .Q(EX_adr[0]) );
  FLIP_FLOP_D EX_bra_confirm_reg ( .D(n554), .CK(clock), .Q(EX_bra_confirm) );
  FLIP_FLOP_D \EX_data_ual_reg[31]  ( .D(n553), .CK(clock), .Q(EX_data_ual[31]) );
  FLIP_FLOP_D \EX_data_ual_reg[30]  ( .D(n552), .CK(clock), .Q(EX_data_ual[30]) );
  FLIP_FLOP_D \EX_data_ual_reg[29]  ( .D(n551), .CK(clock), .Q(EX_data_ual[29]) );
  FLIP_FLOP_D \EX_data_ual_reg[28]  ( .D(n550), .CK(clock), .Q(EX_data_ual[28]) );
  FLIP_FLOP_D \EX_data_ual_reg[27]  ( .D(n549), .CK(clock), .Q(EX_data_ual[27]) );
  FLIP_FLOP_D \EX_data_ual_reg[26]  ( .D(n548), .CK(clock), .Q(EX_data_ual[26]) );
  FLIP_FLOP_D \EX_data_ual_reg[25]  ( .D(n547), .CK(clock), .Q(EX_data_ual[25]) );
  FLIP_FLOP_D \EX_data_ual_reg[24]  ( .D(n546), .CK(clock), .Q(EX_data_ual[24]) );
  FLIP_FLOP_D \EX_data_ual_reg[23]  ( .D(n545), .CK(clock), .Q(EX_data_ual[23]) );
  FLIP_FLOP_D \EX_data_ual_reg[22]  ( .D(n544), .CK(clock), .Q(EX_data_ual[22]) );
  FLIP_FLOP_D \EX_data_ual_reg[21]  ( .D(n543), .CK(clock), .Q(EX_data_ual[21]) );
  FLIP_FLOP_D \EX_data_ual_reg[20]  ( .D(n542), .CK(clock), .Q(EX_data_ual[20]) );
  FLIP_FLOP_D \EX_data_ual_reg[19]  ( .D(n541), .CK(clock), .Q(EX_data_ual[19]) );
  FLIP_FLOP_D \EX_data_ual_reg[18]  ( .D(n540), .CK(clock), .Q(EX_data_ual[18]) );
  FLIP_FLOP_D \EX_data_ual_reg[17]  ( .D(n539), .CK(clock), .Q(EX_data_ual[17]) );
  FLIP_FLOP_D \EX_data_ual_reg[16]  ( .D(n538), .CK(clock), .Q(EX_data_ual[16]) );
  FLIP_FLOP_D \EX_data_ual_reg[15]  ( .D(n537), .CK(clock), .Q(EX_data_ual[15]) );
  FLIP_FLOP_D \EX_data_ual_reg[14]  ( .D(n536), .CK(clock), .Q(EX_data_ual[14]) );
  FLIP_FLOP_D \EX_data_ual_reg[13]  ( .D(n535), .CK(clock), .Q(EX_data_ual[13]) );
  FLIP_FLOP_D \EX_data_ual_reg[12]  ( .D(n534), .CK(clock), .Q(EX_data_ual[12]) );
  FLIP_FLOP_D \EX_data_ual_reg[11]  ( .D(n533), .CK(clock), .Q(EX_data_ual[11]) );
  FLIP_FLOP_D \EX_data_ual_reg[10]  ( .D(n532), .CK(clock), .Q(EX_data_ual[10]) );
  FLIP_FLOP_D \EX_data_ual_reg[9]  ( .D(n531), .CK(clock), .Q(EX_data_ual[9])
         );
  FLIP_FLOP_D \EX_data_ual_reg[8]  ( .D(n530), .CK(clock), .Q(EX_data_ual[8])
         );
  FLIP_FLOP_D \EX_data_ual_reg[7]  ( .D(n529), .CK(clock), .Q(EX_data_ual[7])
         );
  FLIP_FLOP_D \EX_data_ual_reg[6]  ( .D(n528), .CK(clock), .Q(EX_data_ual[6])
         );
  FLIP_FLOP_D \EX_data_ual_reg[5]  ( .D(n527), .CK(clock), .Q(EX_data_ual[5])
         );
  FLIP_FLOP_D \EX_data_ual_reg[4]  ( .D(n526), .CK(clock), .Q(EX_data_ual[4])
         );
  FLIP_FLOP_D \EX_data_ual_reg[3]  ( .D(n525), .CK(clock), .Q(EX_data_ual[3])
         );
  FLIP_FLOP_D \EX_data_ual_reg[2]  ( .D(n524), .CK(clock), .Q(EX_data_ual[2])
         );
  FLIP_FLOP_D \EX_data_ual_reg[1]  ( .D(n523), .CK(clock), .Q(EX_data_ual[1])
         );
  FLIP_FLOP_D \EX_data_ual_reg[0]  ( .D(n522), .CK(clock), .Q(EX_data_ual[0])
         );
  FLIP_FLOP_D \EX_adresse_reg[31]  ( .D(n521), .CK(clock), .Q(EX_adresse[31])
         );
  FLIP_FLOP_D \EX_adresse_reg[30]  ( .D(n520), .CK(clock), .Q(EX_adresse[30])
         );
  FLIP_FLOP_D \EX_adresse_reg[29]  ( .D(n519), .CK(clock), .Q(EX_adresse[29])
         );
  FLIP_FLOP_D \EX_adresse_reg[28]  ( .D(n518), .CK(clock), .Q(EX_adresse[28])
         );
  FLIP_FLOP_D \EX_adresse_reg[27]  ( .D(n517), .CK(clock), .Q(EX_adresse[27])
         );
  FLIP_FLOP_D \EX_adresse_reg[26]  ( .D(n516), .CK(clock), .Q(EX_adresse[26])
         );
  FLIP_FLOP_D \EX_adresse_reg[25]  ( .D(n515), .CK(clock), .Q(EX_adresse[25])
         );
  FLIP_FLOP_D \EX_adresse_reg[24]  ( .D(n514), .CK(clock), .Q(EX_adresse[24])
         );
  FLIP_FLOP_D \EX_adresse_reg[23]  ( .D(n513), .CK(clock), .Q(EX_adresse[23])
         );
  FLIP_FLOP_D \EX_adresse_reg[22]  ( .D(n512), .CK(clock), .Q(EX_adresse[22])
         );
  FLIP_FLOP_D \EX_adresse_reg[21]  ( .D(n511), .CK(clock), .Q(EX_adresse[21])
         );
  FLIP_FLOP_D \EX_adresse_reg[20]  ( .D(n510), .CK(clock), .Q(EX_adresse[20])
         );
  FLIP_FLOP_D \EX_adresse_reg[19]  ( .D(n509), .CK(clock), .Q(EX_adresse[19])
         );
  FLIP_FLOP_D \EX_adresse_reg[18]  ( .D(n508), .CK(clock), .Q(EX_adresse[18])
         );
  FLIP_FLOP_D \EX_adresse_reg[17]  ( .D(n507), .CK(clock), .Q(EX_adresse[17])
         );
  FLIP_FLOP_D \EX_adresse_reg[16]  ( .D(n506), .CK(clock), .Q(EX_adresse[16])
         );
  FLIP_FLOP_D \EX_adresse_reg[15]  ( .D(n505), .CK(clock), .Q(EX_adresse[15])
         );
  FLIP_FLOP_D \EX_adresse_reg[14]  ( .D(n504), .CK(clock), .Q(EX_adresse[14])
         );
  FLIP_FLOP_D \EX_adresse_reg[13]  ( .D(n503), .CK(clock), .Q(EX_adresse[13])
         );
  FLIP_FLOP_D \EX_adresse_reg[12]  ( .D(n502), .CK(clock), .Q(EX_adresse[12])
         );
  FLIP_FLOP_D \EX_adresse_reg[11]  ( .D(n501), .CK(clock), .Q(EX_adresse[11])
         );
  FLIP_FLOP_D \EX_adresse_reg[10]  ( .D(n500), .CK(clock), .Q(EX_adresse[10])
         );
  FLIP_FLOP_D \EX_adresse_reg[9]  ( .D(n499), .CK(clock), .Q(EX_adresse[9]) );
  FLIP_FLOP_D \EX_adresse_reg[8]  ( .D(n498), .CK(clock), .Q(EX_adresse[8]) );
  FLIP_FLOP_D \EX_adresse_reg[7]  ( .D(n497), .CK(clock), .Q(EX_adresse[7]) );
  FLIP_FLOP_D \EX_adresse_reg[6]  ( .D(n496), .CK(clock), .Q(EX_adresse[6]) );
  FLIP_FLOP_D \EX_adresse_reg[5]  ( .D(n495), .CK(clock), .Q(EX_adresse[5]) );
  FLIP_FLOP_D \EX_adresse_reg[4]  ( .D(n494), .CK(clock), .Q(EX_adresse[4]) );
  FLIP_FLOP_D \EX_adresse_reg[3]  ( .D(n493), .CK(clock), .Q(EX_adresse[3]) );
  FLIP_FLOP_D \EX_adresse_reg[2]  ( .D(n492), .CK(clock), .Q(EX_adresse[2]) );
  FLIP_FLOP_D \EX_adresse_reg[1]  ( .D(n491), .CK(clock), .Q(EX_adresse[1]) );
  FLIP_FLOP_D \EX_adresse_reg[0]  ( .D(n490), .CK(clock), .Q(EX_adresse[0]) );
  FLIP_FLOP_D \EX_adr_reg_dest_reg[5]  ( .D(n489), .CK(clock), .Q(
        EX_adr_reg_dest[5]) );
  FLIP_FLOP_D \EX_adr_reg_dest_reg[4]  ( .D(n488), .CK(clock), .Q(
        EX_adr_reg_dest[4]) );
  FLIP_FLOP_D \EX_adr_reg_dest_reg[3]  ( .D(n487), .CK(clock), .Q(
        EX_adr_reg_dest[3]) );
  FLIP_FLOP_D \EX_adr_reg_dest_reg[2]  ( .D(n486), .CK(clock), .Q(
        EX_adr_reg_dest[2]) );
  FLIP_FLOP_D \EX_adr_reg_dest_reg[1]  ( .D(n485), .CK(clock), .Q(
        EX_adr_reg_dest[1]) );
  FLIP_FLOP_D \EX_adr_reg_dest_reg[0]  ( .D(n484), .CK(clock), .Q(
        EX_adr_reg_dest[0]) );
  FLIP_FLOP_D EX_ecr_reg_reg ( .D(n483), .CK(clock), .Q(EX_ecr_reg) );
  FLIP_FLOP_D EX_op_mem_reg ( .D(n482), .CK(clock), .Q(EX_op_mem) );
  FLIP_FLOP_D EX_r_w_reg ( .D(n481), .CK(clock), .Q(EX_r_w) );
  FLIP_FLOP_D \EX_exc_cause_reg[31]  ( .D(n480), .CK(clock), .Q(
        EX_exc_cause[31]) );
  FLIP_FLOP_D \EX_exc_cause_reg[30]  ( .D(n479), .CK(clock), .Q(
        EX_exc_cause[30]) );
  FLIP_FLOP_D \EX_exc_cause_reg[29]  ( .D(n478), .CK(clock), .Q(
        EX_exc_cause[29]) );
  FLIP_FLOP_D \EX_exc_cause_reg[28]  ( .D(n477), .CK(clock), .Q(
        EX_exc_cause[28]) );
  FLIP_FLOP_D \EX_exc_cause_reg[27]  ( .D(n476), .CK(clock), .Q(
        EX_exc_cause[27]) );
  FLIP_FLOP_D \EX_exc_cause_reg[26]  ( .D(n475), .CK(clock), .Q(
        EX_exc_cause[26]) );
  FLIP_FLOP_D \EX_exc_cause_reg[25]  ( .D(n474), .CK(clock), .Q(
        EX_exc_cause[25]) );
  FLIP_FLOP_D \EX_exc_cause_reg[24]  ( .D(n473), .CK(clock), .Q(
        EX_exc_cause[24]) );
  FLIP_FLOP_D \EX_exc_cause_reg[23]  ( .D(n472), .CK(clock), .Q(
        EX_exc_cause[23]) );
  FLIP_FLOP_D \EX_exc_cause_reg[22]  ( .D(n471), .CK(clock), .Q(
        EX_exc_cause[22]) );
  FLIP_FLOP_D \EX_exc_cause_reg[21]  ( .D(n470), .CK(clock), .Q(
        EX_exc_cause[21]) );
  FLIP_FLOP_D \EX_exc_cause_reg[20]  ( .D(n469), .CK(clock), .Q(
        EX_exc_cause[20]) );
  FLIP_FLOP_D \EX_exc_cause_reg[19]  ( .D(n468), .CK(clock), .Q(
        EX_exc_cause[19]) );
  FLIP_FLOP_D \EX_exc_cause_reg[18]  ( .D(n467), .CK(clock), .Q(
        EX_exc_cause[18]) );
  FLIP_FLOP_D \EX_exc_cause_reg[17]  ( .D(n466), .CK(clock), .Q(
        EX_exc_cause[17]) );
  FLIP_FLOP_D \EX_exc_cause_reg[16]  ( .D(n465), .CK(clock), .Q(
        EX_exc_cause[16]) );
  FLIP_FLOP_D \EX_exc_cause_reg[15]  ( .D(n464), .CK(clock), .Q(
        EX_exc_cause[15]) );
  FLIP_FLOP_D \EX_exc_cause_reg[14]  ( .D(n463), .CK(clock), .Q(
        EX_exc_cause[14]) );
  FLIP_FLOP_D \EX_exc_cause_reg[13]  ( .D(n462), .CK(clock), .Q(
        EX_exc_cause[13]) );
  FLIP_FLOP_D \EX_exc_cause_reg[12]  ( .D(n461), .CK(clock), .Q(
        EX_exc_cause[12]) );
  FLIP_FLOP_D \EX_exc_cause_reg[11]  ( .D(n460), .CK(clock), .Q(
        EX_exc_cause[11]) );
  FLIP_FLOP_D \EX_exc_cause_reg[10]  ( .D(n459), .CK(clock), .Q(
        EX_exc_cause[10]) );
  FLIP_FLOP_D \EX_exc_cause_reg[9]  ( .D(n458), .CK(clock), .Q(EX_exc_cause[9]) );
  FLIP_FLOP_D \EX_exc_cause_reg[8]  ( .D(n457), .CK(clock), .Q(EX_exc_cause[8]) );
  FLIP_FLOP_D \EX_exc_cause_reg[7]  ( .D(n456), .CK(clock), .Q(EX_exc_cause[7]) );
  FLIP_FLOP_D \EX_exc_cause_reg[6]  ( .D(n455), .CK(clock), .Q(EX_exc_cause[6]) );
  FLIP_FLOP_D \EX_exc_cause_reg[5]  ( .D(n454), .CK(clock), .Q(EX_exc_cause[5]) );
  FLIP_FLOP_D \EX_exc_cause_reg[4]  ( .D(n453), .CK(clock), .Q(EX_exc_cause[4]) );
  FLIP_FLOP_D \EX_exc_cause_reg[3]  ( .D(n452), .CK(clock), .Q(EX_exc_cause[3]) );
  FLIP_FLOP_D \EX_exc_cause_reg[2]  ( .D(n451), .CK(clock), .Q(EX_exc_cause[2]) );
  FLIP_FLOP_D \EX_exc_cause_reg[1]  ( .D(n450), .CK(clock), .Q(EX_exc_cause[1]) );
  FLIP_FLOP_D \EX_exc_cause_reg[0]  ( .D(n449), .CK(clock), .Q(EX_exc_cause[0]) );
  FLIP_FLOP_D \EX_level_reg[1]  ( .D(n448), .CK(clock), .Q(EX_level[1]) );
  FLIP_FLOP_D \EX_level_reg[0]  ( .D(n447), .CK(clock), .Q(EX_level[0]) );
  NAND_GATE U12 ( .I1(n14), .I2(n15), .O(n447) );
  NAND_GATE U13 ( .I1(n16), .I2(n28), .O(n15) );
  OR_GATE U14 ( .I1(DI_level[0]), .I2(n17), .O(n16) );
  NAND_GATE U15 ( .I1(EX_level[0]), .I2(n25), .O(n14) );
  NAND_GATE U16 ( .I1(n19), .I2(n20), .O(n448) );
  NAND_GATE U17 ( .I1(n21), .I2(n28), .O(n20) );
  OR_GATE U18 ( .I1(DI_level[1]), .I2(n17), .O(n21) );
  NAND_GATE U19 ( .I1(EX_level[1]), .I2(n24), .O(n19) );
  NAND_GATE U20 ( .I1(n22), .I2(n23), .O(n449) );
  NAND_GATE U21 ( .I1(DI_exc_cause[0]), .I2(n4), .O(n23) );
  NAND_GATE U22 ( .I1(EX_exc_cause[0]), .I2(n25), .O(n22) );
  NAND_GATE U36 ( .I1(n37), .I2(n38), .O(n451) );
  NAND_GATE U37 ( .I1(DI_exc_cause[2]), .I2(n4), .O(n38) );
  NAND_GATE U38 ( .I1(EX_exc_cause[2]), .I2(n12), .O(n37) );
  NAND_GATE U39 ( .I1(n39), .I2(n40), .O(n452) );
  NAND_GATE U40 ( .I1(DI_exc_cause[3]), .I2(n4), .O(n40) );
  NAND_GATE U41 ( .I1(EX_exc_cause[3]), .I2(n12), .O(n39) );
  NAND_GATE U42 ( .I1(n41), .I2(n42), .O(n453) );
  NAND_GATE U43 ( .I1(DI_exc_cause[4]), .I2(n4), .O(n42) );
  NAND_GATE U44 ( .I1(EX_exc_cause[4]), .I2(n12), .O(n41) );
  NAND_GATE U45 ( .I1(n43), .I2(n44), .O(n454) );
  NAND_GATE U46 ( .I1(DI_exc_cause[5]), .I2(n4), .O(n44) );
  NAND_GATE U47 ( .I1(EX_exc_cause[5]), .I2(n12), .O(n43) );
  NAND_GATE U48 ( .I1(n45), .I2(n46), .O(n455) );
  NAND_GATE U49 ( .I1(DI_exc_cause[6]), .I2(n4), .O(n46) );
  NAND_GATE U50 ( .I1(EX_exc_cause[6]), .I2(n12), .O(n45) );
  NAND_GATE U51 ( .I1(n47), .I2(n48), .O(n456) );
  NAND_GATE U52 ( .I1(DI_exc_cause[7]), .I2(n4), .O(n48) );
  NAND_GATE U53 ( .I1(EX_exc_cause[7]), .I2(n12), .O(n47) );
  NAND_GATE U54 ( .I1(n49), .I2(n50), .O(n457) );
  NAND_GATE U55 ( .I1(DI_exc_cause[8]), .I2(n4), .O(n50) );
  NAND_GATE U56 ( .I1(EX_exc_cause[8]), .I2(n12), .O(n49) );
  NAND_GATE U57 ( .I1(n51), .I2(n52), .O(n458) );
  NAND_GATE U58 ( .I1(DI_exc_cause[9]), .I2(n4), .O(n52) );
  NAND_GATE U59 ( .I1(EX_exc_cause[9]), .I2(n12), .O(n51) );
  NAND_GATE U60 ( .I1(n53), .I2(n54), .O(n459) );
  NAND_GATE U61 ( .I1(DI_exc_cause[10]), .I2(n4), .O(n54) );
  NAND_GATE U62 ( .I1(EX_exc_cause[10]), .I2(n12), .O(n53) );
  NAND_GATE U63 ( .I1(n55), .I2(n56), .O(n460) );
  NAND_GATE U64 ( .I1(DI_exc_cause[11]), .I2(n4), .O(n56) );
  NAND_GATE U65 ( .I1(EX_exc_cause[11]), .I2(n13), .O(n55) );
  NAND_GATE U66 ( .I1(n57), .I2(n58), .O(n461) );
  NAND_GATE U67 ( .I1(DI_exc_cause[12]), .I2(n4), .O(n58) );
  NAND_GATE U68 ( .I1(EX_exc_cause[12]), .I2(n13), .O(n57) );
  NAND_GATE U69 ( .I1(n59), .I2(n60), .O(n462) );
  NAND_GATE U70 ( .I1(DI_exc_cause[13]), .I2(n4), .O(n60) );
  NAND_GATE U71 ( .I1(EX_exc_cause[13]), .I2(n13), .O(n59) );
  NAND_GATE U72 ( .I1(n61), .I2(n62), .O(n463) );
  NAND_GATE U73 ( .I1(DI_exc_cause[14]), .I2(n4), .O(n62) );
  NAND_GATE U74 ( .I1(EX_exc_cause[14]), .I2(n13), .O(n61) );
  NAND_GATE U75 ( .I1(n63), .I2(n64), .O(n464) );
  NAND_GATE U76 ( .I1(DI_exc_cause[15]), .I2(n4), .O(n64) );
  NAND_GATE U77 ( .I1(EX_exc_cause[15]), .I2(n13), .O(n63) );
  NAND_GATE U78 ( .I1(n65), .I2(n66), .O(n465) );
  NAND_GATE U79 ( .I1(DI_exc_cause[16]), .I2(n4), .O(n66) );
  NAND_GATE U80 ( .I1(EX_exc_cause[16]), .I2(n13), .O(n65) );
  NAND_GATE U81 ( .I1(n67), .I2(n68), .O(n466) );
  NAND_GATE U82 ( .I1(DI_exc_cause[17]), .I2(n4), .O(n68) );
  NAND_GATE U83 ( .I1(EX_exc_cause[17]), .I2(n13), .O(n67) );
  NAND_GATE U84 ( .I1(n69), .I2(n70), .O(n467) );
  NAND_GATE U85 ( .I1(DI_exc_cause[18]), .I2(n4), .O(n70) );
  NAND_GATE U86 ( .I1(EX_exc_cause[18]), .I2(n13), .O(n69) );
  NAND_GATE U87 ( .I1(n71), .I2(n72), .O(n468) );
  NAND_GATE U88 ( .I1(DI_exc_cause[19]), .I2(n4), .O(n72) );
  NAND_GATE U89 ( .I1(EX_exc_cause[19]), .I2(n13), .O(n71) );
  NAND_GATE U90 ( .I1(n73), .I2(n74), .O(n469) );
  NAND_GATE U91 ( .I1(DI_exc_cause[20]), .I2(n4), .O(n74) );
  NAND_GATE U92 ( .I1(EX_exc_cause[20]), .I2(n18), .O(n73) );
  NAND_GATE U93 ( .I1(n75), .I2(n76), .O(n470) );
  NAND_GATE U94 ( .I1(DI_exc_cause[21]), .I2(n4), .O(n76) );
  NAND_GATE U95 ( .I1(EX_exc_cause[21]), .I2(n18), .O(n75) );
  NAND_GATE U96 ( .I1(n77), .I2(n78), .O(n471) );
  NAND_GATE U97 ( .I1(DI_exc_cause[22]), .I2(n4), .O(n78) );
  NAND_GATE U98 ( .I1(EX_exc_cause[22]), .I2(n18), .O(n77) );
  NAND_GATE U99 ( .I1(n79), .I2(n80), .O(n472) );
  NAND_GATE U100 ( .I1(DI_exc_cause[23]), .I2(n4), .O(n80) );
  NAND_GATE U101 ( .I1(EX_exc_cause[23]), .I2(n18), .O(n79) );
  NAND_GATE U102 ( .I1(n81), .I2(n82), .O(n473) );
  NAND_GATE U103 ( .I1(DI_exc_cause[24]), .I2(n4), .O(n82) );
  NAND_GATE U104 ( .I1(EX_exc_cause[24]), .I2(n18), .O(n81) );
  NAND_GATE U105 ( .I1(n83), .I2(n84), .O(n474) );
  NAND_GATE U106 ( .I1(DI_exc_cause[25]), .I2(n4), .O(n84) );
  NAND_GATE U107 ( .I1(EX_exc_cause[25]), .I2(n18), .O(n83) );
  NAND_GATE U108 ( .I1(n85), .I2(n86), .O(n475) );
  NAND_GATE U109 ( .I1(DI_exc_cause[26]), .I2(n4), .O(n86) );
  NAND_GATE U110 ( .I1(EX_exc_cause[26]), .I2(n18), .O(n85) );
  NAND_GATE U111 ( .I1(n87), .I2(n88), .O(n476) );
  NAND_GATE U112 ( .I1(DI_exc_cause[27]), .I2(n4), .O(n88) );
  NAND_GATE U113 ( .I1(EX_exc_cause[27]), .I2(n18), .O(n87) );
  NAND_GATE U114 ( .I1(n89), .I2(n90), .O(n477) );
  NAND_GATE U115 ( .I1(DI_exc_cause[28]), .I2(n4), .O(n90) );
  NAND_GATE U116 ( .I1(EX_exc_cause[28]), .I2(n18), .O(n89) );
  NAND_GATE U117 ( .I1(n91), .I2(n92), .O(n478) );
  NAND_GATE U118 ( .I1(DI_exc_cause[29]), .I2(n4), .O(n92) );
  NAND_GATE U119 ( .I1(EX_exc_cause[29]), .I2(n18), .O(n91) );
  NAND_GATE U120 ( .I1(n93), .I2(n94), .O(n479) );
  NAND_GATE U121 ( .I1(DI_exc_cause[30]), .I2(n4), .O(n94) );
  NAND_GATE U122 ( .I1(EX_exc_cause[30]), .I2(n13), .O(n93) );
  NAND_GATE U123 ( .I1(n95), .I2(n96), .O(n480) );
  NAND_GATE U124 ( .I1(DI_exc_cause[31]), .I2(n4), .O(n96) );
  NAND_GATE U125 ( .I1(EX_exc_cause[31]), .I2(n12), .O(n95) );
  NAND_GATE U126 ( .I1(n97), .I2(n98), .O(n481) );
  NAND_GATE U127 ( .I1(DI_r_w), .I2(n4), .O(n98) );
  NAND_GATE U128 ( .I1(EX_r_w), .I2(n25), .O(n97) );
  NAND_GATE U129 ( .I1(n99), .I2(n100), .O(n482) );
  NAND_GATE U130 ( .I1(DI_op_mem), .I2(n4), .O(n100) );
  NAND_GATE U131 ( .I1(EX_op_mem), .I2(n24), .O(n99) );
  NAND_GATE U136 ( .I1(n106), .I2(n107), .O(n484) );
  NAND_GATE U137 ( .I1(DI_adr_reg_dest[0]), .I2(n4), .O(n107) );
  NAND_GATE U138 ( .I1(EX_adr_reg_dest[0]), .I2(n18), .O(n106) );
  NAND_GATE U139 ( .I1(n108), .I2(n109), .O(n485) );
  NAND_GATE U140 ( .I1(DI_adr_reg_dest[1]), .I2(n4), .O(n109) );
  NAND_GATE U141 ( .I1(EX_adr_reg_dest[1]), .I2(n13), .O(n108) );
  NAND_GATE U142 ( .I1(n110), .I2(n111), .O(n486) );
  NAND_GATE U143 ( .I1(DI_adr_reg_dest[2]), .I2(n4), .O(n111) );
  NAND_GATE U144 ( .I1(EX_adr_reg_dest[2]), .I2(n12), .O(n110) );
  NAND_GATE U145 ( .I1(n112), .I2(n113), .O(n487) );
  NAND_GATE U146 ( .I1(DI_adr_reg_dest[3]), .I2(n4), .O(n113) );
  NAND_GATE U147 ( .I1(EX_adr_reg_dest[3]), .I2(n25), .O(n112) );
  NAND_GATE U148 ( .I1(n114), .I2(n115), .O(n488) );
  NAND_GATE U149 ( .I1(DI_adr_reg_dest[4]), .I2(n4), .O(n115) );
  NAND_GATE U150 ( .I1(EX_adr_reg_dest[4]), .I2(n18), .O(n114) );
  NAND_GATE U151 ( .I1(n116), .I2(n117), .O(n489) );
  NAND_GATE U152 ( .I1(DI_adr_reg_dest[5]), .I2(n4), .O(n117) );
  NAND_GATE U153 ( .I1(EX_adr_reg_dest[5]), .I2(n13), .O(n116) );
  NAND3_GATE U289 ( .I1(n221), .I2(n222), .I3(n223), .O(n523) );
  NAND_GATE U290 ( .I1(EX_data_ual[1]), .I2(n10), .O(n223) );
  NAND_GATE U291 ( .I1(res_ual[1]), .I2(n2), .O(n222) );
  NAND_GATE U292 ( .I1(N11), .I2(n1), .O(n221) );
  NAND3_GATE U293 ( .I1(n224), .I2(n225), .I3(n226), .O(n524) );
  NAND_GATE U294 ( .I1(EX_data_ual[2]), .I2(n9), .O(n226) );
  NAND_GATE U295 ( .I1(res_ual[2]), .I2(n2), .O(n225) );
  NAND_GATE U296 ( .I1(N12), .I2(n1), .O(n224) );
  NAND3_GATE U297 ( .I1(n227), .I2(n228), .I3(n229), .O(n525) );
  NAND_GATE U298 ( .I1(EX_data_ual[3]), .I2(n8), .O(n229) );
  NAND_GATE U299 ( .I1(res_ual[3]), .I2(n2), .O(n228) );
  NAND_GATE U300 ( .I1(N13), .I2(n1), .O(n227) );
  NAND3_GATE U301 ( .I1(n230), .I2(n231), .I3(n232), .O(n526) );
  NAND_GATE U302 ( .I1(EX_data_ual[4]), .I2(n594), .O(n232) );
  NAND_GATE U303 ( .I1(res_ual[4]), .I2(n2), .O(n231) );
  NAND_GATE U304 ( .I1(N14), .I2(n1), .O(n230) );
  NAND3_GATE U305 ( .I1(n233), .I2(n234), .I3(n235), .O(n527) );
  NAND_GATE U306 ( .I1(EX_data_ual[5]), .I2(n594), .O(n235) );
  NAND_GATE U307 ( .I1(res_ual[5]), .I2(n2), .O(n234) );
  NAND_GATE U308 ( .I1(N15), .I2(n1), .O(n233) );
  NAND3_GATE U309 ( .I1(n236), .I2(n237), .I3(n238), .O(n528) );
  NAND_GATE U310 ( .I1(EX_data_ual[6]), .I2(n594), .O(n238) );
  NAND_GATE U311 ( .I1(res_ual[6]), .I2(n2), .O(n237) );
  NAND_GATE U312 ( .I1(N16), .I2(n1), .O(n236) );
  NAND3_GATE U313 ( .I1(n239), .I2(n240), .I3(n241), .O(n529) );
  NAND_GATE U314 ( .I1(EX_data_ual[7]), .I2(n594), .O(n241) );
  NAND_GATE U315 ( .I1(res_ual[7]), .I2(n2), .O(n240) );
  NAND_GATE U316 ( .I1(N17), .I2(n1), .O(n239) );
  NAND_GATE U420 ( .I1(n316), .I2(n317), .O(n555) );
  NAND_GATE U421 ( .I1(DI_adr[0]), .I2(n5), .O(n317) );
  NAND_GATE U422 ( .I1(EX_adr[0]), .I2(n24), .O(n316) );
  NAND_GATE U423 ( .I1(n318), .I2(n319), .O(n556) );
  NAND_GATE U424 ( .I1(DI_adr[1]), .I2(n5), .O(n319) );
  NAND_GATE U425 ( .I1(EX_adr[1]), .I2(n24), .O(n318) );
  NAND_GATE U426 ( .I1(n320), .I2(n321), .O(n557) );
  NAND_GATE U427 ( .I1(DI_adr[2]), .I2(n5), .O(n321) );
  NAND_GATE U428 ( .I1(EX_adr[2]), .I2(n24), .O(n320) );
  NAND_GATE U429 ( .I1(n322), .I2(n323), .O(n558) );
  NAND_GATE U430 ( .I1(DI_adr[3]), .I2(n5), .O(n323) );
  NAND_GATE U431 ( .I1(EX_adr[3]), .I2(n24), .O(n322) );
  NAND_GATE U432 ( .I1(n324), .I2(n325), .O(n559) );
  NAND_GATE U433 ( .I1(DI_adr[4]), .I2(n5), .O(n325) );
  NAND_GATE U434 ( .I1(EX_adr[4]), .I2(n24), .O(n324) );
  NAND_GATE U435 ( .I1(n326), .I2(n327), .O(n560) );
  NAND_GATE U436 ( .I1(DI_adr[5]), .I2(n5), .O(n327) );
  NAND_GATE U437 ( .I1(EX_adr[5]), .I2(n24), .O(n326) );
  NAND_GATE U438 ( .I1(n328), .I2(n329), .O(n561) );
  NAND_GATE U439 ( .I1(DI_adr[6]), .I2(n5), .O(n329) );
  NAND_GATE U440 ( .I1(EX_adr[6]), .I2(n24), .O(n328) );
  NAND_GATE U441 ( .I1(n330), .I2(n331), .O(n562) );
  NAND_GATE U442 ( .I1(DI_adr[7]), .I2(n5), .O(n331) );
  NAND_GATE U443 ( .I1(EX_adr[7]), .I2(n24), .O(n330) );
  NAND_GATE U444 ( .I1(n332), .I2(n333), .O(n563) );
  NAND_GATE U445 ( .I1(DI_adr[8]), .I2(n5), .O(n333) );
  NAND_GATE U446 ( .I1(EX_adr[8]), .I2(n24), .O(n332) );
  NAND_GATE U447 ( .I1(n334), .I2(n335), .O(n564) );
  NAND_GATE U448 ( .I1(DI_adr[9]), .I2(n5), .O(n335) );
  NAND_GATE U449 ( .I1(EX_adr[9]), .I2(n18), .O(n334) );
  NAND_GATE U450 ( .I1(n336), .I2(n337), .O(n565) );
  NAND_GATE U451 ( .I1(DI_adr[10]), .I2(n5), .O(n337) );
  NAND_GATE U452 ( .I1(EX_adr[10]), .I2(n13), .O(n336) );
  NAND_GATE U453 ( .I1(n338), .I2(n339), .O(n566) );
  NAND_GATE U454 ( .I1(DI_adr[11]), .I2(n5), .O(n339) );
  NAND_GATE U455 ( .I1(EX_adr[11]), .I2(n12), .O(n338) );
  NAND_GATE U456 ( .I1(n340), .I2(n341), .O(n567) );
  NAND_GATE U457 ( .I1(DI_adr[12]), .I2(n5), .O(n341) );
  NAND_GATE U458 ( .I1(EX_adr[12]), .I2(n25), .O(n340) );
  NAND_GATE U459 ( .I1(n342), .I2(n343), .O(n568) );
  NAND_GATE U460 ( .I1(DI_adr[13]), .I2(n5), .O(n343) );
  NAND_GATE U461 ( .I1(EX_adr[13]), .I2(n24), .O(n342) );
  NAND_GATE U462 ( .I1(n344), .I2(n345), .O(n569) );
  NAND_GATE U463 ( .I1(DI_adr[14]), .I2(n5), .O(n345) );
  NAND_GATE U464 ( .I1(EX_adr[14]), .I2(n18), .O(n344) );
  NAND_GATE U465 ( .I1(n346), .I2(n347), .O(n570) );
  NAND_GATE U466 ( .I1(DI_adr[15]), .I2(n5), .O(n347) );
  NAND_GATE U467 ( .I1(EX_adr[15]), .I2(n13), .O(n346) );
  NAND_GATE U468 ( .I1(n348), .I2(n349), .O(n571) );
  NAND_GATE U469 ( .I1(DI_adr[16]), .I2(n5), .O(n349) );
  NAND_GATE U470 ( .I1(EX_adr[16]), .I2(n12), .O(n348) );
  NAND_GATE U471 ( .I1(n350), .I2(n351), .O(n572) );
  NAND_GATE U472 ( .I1(DI_adr[17]), .I2(n5), .O(n351) );
  NAND_GATE U473 ( .I1(EX_adr[17]), .I2(n25), .O(n350) );
  NAND_GATE U474 ( .I1(n352), .I2(n353), .O(n573) );
  NAND_GATE U475 ( .I1(DI_adr[18]), .I2(n5), .O(n353) );
  NAND_GATE U476 ( .I1(EX_adr[18]), .I2(n25), .O(n352) );
  NAND_GATE U477 ( .I1(n354), .I2(n355), .O(n574) );
  NAND_GATE U478 ( .I1(DI_adr[19]), .I2(n5), .O(n355) );
  NAND_GATE U479 ( .I1(EX_adr[19]), .I2(n25), .O(n354) );
  NAND_GATE U480 ( .I1(n356), .I2(n357), .O(n575) );
  NAND_GATE U481 ( .I1(DI_adr[20]), .I2(n5), .O(n357) );
  NAND_GATE U482 ( .I1(EX_adr[20]), .I2(n25), .O(n356) );
  NAND_GATE U483 ( .I1(n358), .I2(n359), .O(n576) );
  NAND_GATE U484 ( .I1(DI_adr[21]), .I2(n5), .O(n359) );
  NAND_GATE U485 ( .I1(EX_adr[21]), .I2(n25), .O(n358) );
  NAND_GATE U486 ( .I1(n360), .I2(n361), .O(n577) );
  NAND_GATE U487 ( .I1(DI_adr[22]), .I2(n5), .O(n361) );
  NAND_GATE U488 ( .I1(EX_adr[22]), .I2(n25), .O(n360) );
  NAND_GATE U489 ( .I1(n362), .I2(n363), .O(n578) );
  NAND_GATE U490 ( .I1(DI_adr[23]), .I2(n5), .O(n363) );
  NAND_GATE U491 ( .I1(EX_adr[23]), .I2(n25), .O(n362) );
  NAND_GATE U492 ( .I1(n364), .I2(n365), .O(n579) );
  NAND_GATE U493 ( .I1(DI_adr[24]), .I2(n5), .O(n365) );
  NAND_GATE U494 ( .I1(EX_adr[24]), .I2(n25), .O(n364) );
  NAND_GATE U495 ( .I1(n366), .I2(n367), .O(n580) );
  NAND_GATE U496 ( .I1(DI_adr[25]), .I2(n5), .O(n367) );
  NAND_GATE U497 ( .I1(EX_adr[25]), .I2(n25), .O(n366) );
  NAND_GATE U498 ( .I1(n368), .I2(n369), .O(n581) );
  NAND_GATE U499 ( .I1(DI_adr[26]), .I2(n5), .O(n369) );
  NAND_GATE U500 ( .I1(EX_adr[26]), .I2(n25), .O(n368) );
  NAND_GATE U501 ( .I1(n370), .I2(n371), .O(n582) );
  NAND_GATE U502 ( .I1(DI_adr[27]), .I2(n5), .O(n371) );
  NAND_GATE U503 ( .I1(EX_adr[27]), .I2(n24), .O(n370) );
  NAND_GATE U504 ( .I1(n372), .I2(n373), .O(n583) );
  NAND_GATE U505 ( .I1(DI_adr[28]), .I2(n5), .O(n373) );
  NAND_GATE U506 ( .I1(EX_adr[28]), .I2(n24), .O(n372) );
  NAND_GATE U507 ( .I1(n374), .I2(n375), .O(n584) );
  NAND_GATE U508 ( .I1(DI_adr[29]), .I2(n5), .O(n375) );
  NAND_GATE U509 ( .I1(EX_adr[29]), .I2(n24), .O(n374) );
  NAND_GATE U510 ( .I1(n376), .I2(n377), .O(n585) );
  NAND_GATE U511 ( .I1(DI_adr[30]), .I2(n5), .O(n377) );
  NAND_GATE U512 ( .I1(EX_adr[30]), .I2(n18), .O(n376) );
  NAND_GATE U513 ( .I1(n378), .I2(n379), .O(n586) );
  NAND_GATE U514 ( .I1(DI_adr[31]), .I2(n5), .O(n379) );
  NAND_GATE U515 ( .I1(EX_adr[31]), .I2(n13), .O(n378) );
  NAND_GATE U516 ( .I1(n381), .I2(n382), .O(n587) );
  NAND_GATE U517 ( .I1(DI_it_ok), .I2(n4), .O(n382) );
  NAND_GATE U520 ( .I1(EX_it_ok), .I2(n12), .O(n381) );
  alu U1_alu ( .clock(clock), .reset(reset), .op1(DI_op1), .op2(DI_op2), 
        .ctrl(DI_code_ual), .res(res_ual), .overflow(overflow_ual) );
  pps_ex_DW01_add_0 add_183 ( .A(DI_offset), .B(base_adr), .CI(1'b0), .SUM({
        N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, 
        N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82}) );
  pps_ex_DW01_add_1 r87 ( .A(DI_adr), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N41, N40, N39, N38, N37, N36, N35, N34, 
        N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, 
        N19, N18, N17, N16, N15, N14, N13, N12, N11, N10}) );
  AND_GATE U3 ( .I1(DI_link), .I2(n3), .O(n1) );
  AND_GATE U4 ( .I1(n30), .I2(n3), .O(n2) );
  AND_GATE U5 ( .I1(n29), .I2(n28), .O(n3) );
  AND_GATE U6 ( .I1(n27), .I2(n29), .O(n4) );
  NOR_GATE U7 ( .I1(reset), .I2(stop_all), .O(n5) );
  OR_GATE U8 ( .I1(res_ual[0]), .I2(n6), .O(n189) );
  INV_GATE U9 ( .I1(DI_bra), .O(n6) );
  AND_GATE U10 ( .I1(DI_bra), .I2(res_ual[0]), .O(n7) );
  INV_GATE U11 ( .I1(n28), .O(n8) );
  INV_GATE U23 ( .I1(n28), .O(n9) );
  INV_GATE U24 ( .I1(n28), .O(n10) );
  INV_GATE U25 ( .I1(n28), .O(n11) );
  INV_GATE U26 ( .I1(n28), .O(n12) );
  INV_GATE U27 ( .I1(n28), .O(n13) );
  INV_GATE U28 ( .I1(n28), .O(n18) );
  INV_GATE U29 ( .I1(n28), .O(n24) );
  INV_GATE U30 ( .I1(n28), .O(n25) );
  INV_GATE U31 ( .I1(DI_mode), .O(n26) );
  INV_GATE U32 ( .I1(stop_all), .O(n27) );
  OR_GATE U33 ( .I1(reset), .I2(n27), .O(n28) );
  INV_GATE U34 ( .I1(n28), .O(n594) );
  OR_GATE U35 ( .I1(reset), .I2(clear), .O(n17) );
  INV_GATE U132 ( .I1(n17), .O(n29) );
  INV_GATE U133 ( .I1(DI_link), .O(n30) );
  NAND_GATE U134 ( .I1(EX_exc_cause[1]), .I2(n8), .O(n121) );
  NOR_GATE U135 ( .I1(DI_exc_cause[2]), .I2(DI_exc_cause[3]), .O(n31) );
  AND_GATE U154 ( .I1(overflow_ual), .I2(n31), .O(n105) );
  OR4_GATE U155 ( .I1(DI_exc_cause[4]), .I2(DI_exc_cause[5]), .I3(
        DI_exc_cause[6]), .I4(DI_exc_cause[7]), .O(n34) );
  OR4_GATE U156 ( .I1(DI_exc_cause[12]), .I2(DI_exc_cause[13]), .I3(
        DI_exc_cause[14]), .I4(DI_exc_cause[15]), .O(n33) );
  OR4_GATE U157 ( .I1(DI_exc_cause[8]), .I2(DI_exc_cause[9]), .I3(
        DI_exc_cause[10]), .I4(DI_exc_cause[11]), .O(n32) );
  NOR4_GATE U158 ( .I1(n34), .I2(DI_exc_cause[0]), .I3(n33), .I4(n32), .O(n104) );
  NOR4_GATE U159 ( .I1(DI_exc_cause[18]), .I2(DI_exc_cause[19]), .I3(
        DI_exc_cause[16]), .I4(DI_exc_cause[17]), .O(n102) );
  NOR4_GATE U160 ( .I1(DI_exc_cause[22]), .I2(DI_exc_cause[23]), .I3(
        DI_exc_cause[20]), .I4(DI_exc_cause[21]), .O(n101) );
  NOR4_GATE U161 ( .I1(DI_exc_cause[26]), .I2(DI_exc_cause[27]), .I3(
        DI_exc_cause[24]), .I4(DI_exc_cause[25]), .O(n36) );
  NOR4_GATE U162 ( .I1(DI_exc_cause[30]), .I2(DI_exc_cause[31]), .I3(
        DI_exc_cause[28]), .I4(DI_exc_cause[29]), .O(n35) );
  AND4_GATE U163 ( .I1(n102), .I2(n101), .I3(n36), .I4(n35), .O(n103) );
  AND3_GATE U164 ( .I1(n105), .I2(n104), .I3(n103), .O(n118) );
  OR_GATE U165 ( .I1(DI_exc_cause[1]), .I2(n118), .O(n119) );
  NAND_GATE U166 ( .I1(n3), .I2(n119), .O(n120) );
  NAND_GATE U167 ( .I1(n121), .I2(n120), .O(n450) );
  NAND_GATE U168 ( .I1(n1), .I2(n7), .O(n124) );
  NAND_GATE U169 ( .I1(DI_ecr_reg), .I2(n2), .O(n123) );
  NAND_GATE U170 ( .I1(EX_ecr_reg), .I2(n8), .O(n122) );
  NAND3_GATE U171 ( .I1(n124), .I2(n123), .I3(n122), .O(n483) );
  NAND_GATE U172 ( .I1(DI_mode), .I2(DI_adr[31]), .O(n126) );
  NAND_GATE U173 ( .I1(DI_op1[31]), .I2(n26), .O(n125) );
  NAND_GATE U174 ( .I1(n126), .I2(n125), .O(base_adr[31]) );
  NAND_GATE U175 ( .I1(DI_adr[30]), .I2(DI_mode), .O(n128) );
  NAND_GATE U176 ( .I1(DI_op1[30]), .I2(n26), .O(n127) );
  NAND_GATE U177 ( .I1(n128), .I2(n127), .O(base_adr[30]) );
  NAND_GATE U178 ( .I1(DI_adr[29]), .I2(DI_mode), .O(n130) );
  NAND_GATE U179 ( .I1(DI_op1[29]), .I2(n26), .O(n129) );
  NAND_GATE U180 ( .I1(n130), .I2(n129), .O(base_adr[29]) );
  NAND_GATE U181 ( .I1(DI_adr[28]), .I2(DI_mode), .O(n132) );
  NAND_GATE U182 ( .I1(DI_op1[28]), .I2(n26), .O(n131) );
  NAND_GATE U183 ( .I1(n132), .I2(n131), .O(base_adr[28]) );
  NAND_GATE U184 ( .I1(DI_adr[27]), .I2(DI_mode), .O(n134) );
  NAND_GATE U185 ( .I1(DI_op1[27]), .I2(n26), .O(n133) );
  NAND_GATE U186 ( .I1(n134), .I2(n133), .O(base_adr[27]) );
  NAND_GATE U187 ( .I1(DI_adr[26]), .I2(DI_mode), .O(n136) );
  NAND_GATE U188 ( .I1(DI_op1[26]), .I2(n26), .O(n135) );
  NAND_GATE U189 ( .I1(n136), .I2(n135), .O(base_adr[26]) );
  NAND_GATE U190 ( .I1(DI_adr[25]), .I2(DI_mode), .O(n138) );
  NAND_GATE U191 ( .I1(DI_op1[25]), .I2(n26), .O(n137) );
  NAND_GATE U192 ( .I1(n138), .I2(n137), .O(base_adr[25]) );
  NAND_GATE U193 ( .I1(DI_adr[24]), .I2(DI_mode), .O(n140) );
  NAND_GATE U194 ( .I1(DI_op1[24]), .I2(n26), .O(n139) );
  NAND_GATE U195 ( .I1(n140), .I2(n139), .O(base_adr[24]) );
  NAND_GATE U196 ( .I1(DI_adr[23]), .I2(DI_mode), .O(n142) );
  NAND_GATE U197 ( .I1(DI_op1[23]), .I2(n26), .O(n141) );
  NAND_GATE U198 ( .I1(n142), .I2(n141), .O(base_adr[23]) );
  NAND_GATE U199 ( .I1(DI_adr[22]), .I2(DI_mode), .O(n144) );
  NAND_GATE U200 ( .I1(DI_op1[22]), .I2(n26), .O(n143) );
  NAND_GATE U201 ( .I1(n144), .I2(n143), .O(base_adr[22]) );
  NAND_GATE U202 ( .I1(DI_adr[21]), .I2(DI_mode), .O(n146) );
  NAND_GATE U203 ( .I1(DI_op1[21]), .I2(n26), .O(n145) );
  NAND_GATE U204 ( .I1(n146), .I2(n145), .O(base_adr[21]) );
  NAND_GATE U205 ( .I1(DI_adr[20]), .I2(DI_mode), .O(n148) );
  NAND_GATE U206 ( .I1(DI_op1[20]), .I2(n26), .O(n147) );
  NAND_GATE U207 ( .I1(n148), .I2(n147), .O(base_adr[20]) );
  NAND_GATE U208 ( .I1(DI_adr[19]), .I2(DI_mode), .O(n150) );
  NAND_GATE U209 ( .I1(DI_op1[19]), .I2(n26), .O(n149) );
  NAND_GATE U210 ( .I1(n150), .I2(n149), .O(base_adr[19]) );
  NAND_GATE U211 ( .I1(DI_adr[18]), .I2(DI_mode), .O(n152) );
  NAND_GATE U212 ( .I1(DI_op1[18]), .I2(n26), .O(n151) );
  NAND_GATE U213 ( .I1(n152), .I2(n151), .O(base_adr[18]) );
  NAND_GATE U214 ( .I1(DI_adr[17]), .I2(DI_mode), .O(n154) );
  NAND_GATE U215 ( .I1(DI_op1[17]), .I2(n26), .O(n153) );
  NAND_GATE U216 ( .I1(n154), .I2(n153), .O(base_adr[17]) );
  NAND_GATE U217 ( .I1(DI_adr[16]), .I2(DI_mode), .O(n156) );
  NAND_GATE U218 ( .I1(DI_op1[16]), .I2(n26), .O(n155) );
  NAND_GATE U219 ( .I1(n156), .I2(n155), .O(base_adr[16]) );
  NAND_GATE U220 ( .I1(DI_adr[15]), .I2(DI_mode), .O(n158) );
  NAND_GATE U221 ( .I1(DI_op1[15]), .I2(n26), .O(n157) );
  NAND_GATE U222 ( .I1(n158), .I2(n157), .O(base_adr[15]) );
  NAND_GATE U223 ( .I1(DI_adr[14]), .I2(DI_mode), .O(n160) );
  NAND_GATE U224 ( .I1(DI_op1[14]), .I2(n26), .O(n159) );
  NAND_GATE U225 ( .I1(n160), .I2(n159), .O(base_adr[14]) );
  NAND_GATE U226 ( .I1(DI_adr[13]), .I2(DI_mode), .O(n162) );
  NAND_GATE U227 ( .I1(DI_op1[13]), .I2(n26), .O(n161) );
  NAND_GATE U228 ( .I1(n162), .I2(n161), .O(base_adr[13]) );
  NAND_GATE U229 ( .I1(DI_adr[12]), .I2(DI_mode), .O(n164) );
  NAND_GATE U230 ( .I1(DI_op1[12]), .I2(n26), .O(n163) );
  NAND_GATE U231 ( .I1(n164), .I2(n163), .O(base_adr[12]) );
  NAND_GATE U232 ( .I1(DI_adr[11]), .I2(DI_mode), .O(n166) );
  NAND_GATE U233 ( .I1(DI_op1[11]), .I2(n26), .O(n165) );
  NAND_GATE U234 ( .I1(n166), .I2(n165), .O(base_adr[11]) );
  NAND_GATE U235 ( .I1(DI_adr[10]), .I2(DI_mode), .O(n168) );
  NAND_GATE U236 ( .I1(DI_op1[10]), .I2(n26), .O(n167) );
  NAND_GATE U237 ( .I1(n168), .I2(n167), .O(base_adr[10]) );
  NAND_GATE U238 ( .I1(DI_adr[9]), .I2(DI_mode), .O(n170) );
  NAND_GATE U239 ( .I1(DI_op1[9]), .I2(n26), .O(n169) );
  NAND_GATE U240 ( .I1(n170), .I2(n169), .O(base_adr[9]) );
  NAND_GATE U241 ( .I1(DI_adr[8]), .I2(DI_mode), .O(n172) );
  NAND_GATE U242 ( .I1(DI_op1[8]), .I2(n26), .O(n171) );
  NAND_GATE U243 ( .I1(n172), .I2(n171), .O(base_adr[8]) );
  NAND_GATE U244 ( .I1(DI_adr[7]), .I2(DI_mode), .O(n174) );
  NAND_GATE U245 ( .I1(DI_op1[7]), .I2(n26), .O(n173) );
  NAND_GATE U246 ( .I1(n174), .I2(n173), .O(base_adr[7]) );
  NAND_GATE U247 ( .I1(DI_adr[6]), .I2(DI_mode), .O(n176) );
  NAND_GATE U248 ( .I1(DI_op1[6]), .I2(n26), .O(n175) );
  NAND_GATE U249 ( .I1(n176), .I2(n175), .O(base_adr[6]) );
  NAND_GATE U250 ( .I1(DI_adr[5]), .I2(DI_mode), .O(n178) );
  NAND_GATE U251 ( .I1(DI_op1[5]), .I2(n26), .O(n177) );
  NAND_GATE U252 ( .I1(n178), .I2(n177), .O(base_adr[5]) );
  NAND_GATE U253 ( .I1(DI_adr[4]), .I2(DI_mode), .O(n180) );
  NAND_GATE U254 ( .I1(DI_op1[4]), .I2(n26), .O(n179) );
  NAND_GATE U255 ( .I1(n180), .I2(n179), .O(base_adr[4]) );
  NAND_GATE U256 ( .I1(DI_adr[3]), .I2(DI_mode), .O(n182) );
  NAND_GATE U257 ( .I1(DI_op1[3]), .I2(n26), .O(n181) );
  NAND_GATE U258 ( .I1(n182), .I2(n181), .O(base_adr[3]) );
  NAND_GATE U259 ( .I1(DI_adr[2]), .I2(DI_mode), .O(n184) );
  NAND_GATE U260 ( .I1(DI_op1[2]), .I2(n26), .O(n183) );
  NAND_GATE U261 ( .I1(n184), .I2(n183), .O(base_adr[2]) );
  NAND_GATE U262 ( .I1(DI_adr[1]), .I2(DI_mode), .O(n186) );
  NAND_GATE U263 ( .I1(DI_op1[1]), .I2(n26), .O(n185) );
  NAND_GATE U264 ( .I1(n186), .I2(n185), .O(base_adr[1]) );
  NAND_GATE U265 ( .I1(DI_adr[0]), .I2(DI_mode), .O(n188) );
  NAND_GATE U266 ( .I1(DI_op1[0]), .I2(n26), .O(n187) );
  NAND_GATE U267 ( .I1(n188), .I2(n187), .O(base_adr[0]) );
  AND_GATE U268 ( .I1(n3), .I2(n189), .O(n305) );
  NAND_GATE U269 ( .I1(N82), .I2(n305), .O(n193) );
  NAND_GATE U270 ( .I1(DI_bra), .I2(n3), .O(n190) );
  NOR_GATE U271 ( .I1(res_ual[0]), .I2(n190), .O(n306) );
  NAND_GATE U272 ( .I1(N10), .I2(n306), .O(n192) );
  NAND_GATE U273 ( .I1(EX_adresse[0]), .I2(n8), .O(n191) );
  NAND3_GATE U274 ( .I1(n193), .I2(n192), .I3(n191), .O(n490) );
  NAND_GATE U275 ( .I1(N83), .I2(n305), .O(n196) );
  NAND_GATE U276 ( .I1(N11), .I2(n306), .O(n195) );
  NAND_GATE U277 ( .I1(EX_adresse[1]), .I2(n8), .O(n194) );
  NAND3_GATE U278 ( .I1(n196), .I2(n195), .I3(n194), .O(n491) );
  NAND_GATE U279 ( .I1(N84), .I2(n305), .O(n199) );
  NAND_GATE U280 ( .I1(N12), .I2(n306), .O(n198) );
  NAND_GATE U281 ( .I1(EX_adresse[2]), .I2(n8), .O(n197) );
  NAND3_GATE U282 ( .I1(n199), .I2(n198), .I3(n197), .O(n492) );
  NAND_GATE U283 ( .I1(N85), .I2(n305), .O(n202) );
  NAND_GATE U284 ( .I1(N13), .I2(n306), .O(n201) );
  NAND_GATE U285 ( .I1(EX_adresse[3]), .I2(n8), .O(n200) );
  NAND3_GATE U286 ( .I1(n202), .I2(n201), .I3(n200), .O(n493) );
  NAND_GATE U287 ( .I1(N86), .I2(n305), .O(n205) );
  NAND_GATE U288 ( .I1(N14), .I2(n306), .O(n204) );
  NAND_GATE U317 ( .I1(EX_adresse[4]), .I2(n8), .O(n203) );
  NAND3_GATE U318 ( .I1(n205), .I2(n204), .I3(n203), .O(n494) );
  NAND_GATE U319 ( .I1(N87), .I2(n305), .O(n208) );
  NAND_GATE U320 ( .I1(N15), .I2(n306), .O(n207) );
  NAND_GATE U321 ( .I1(EX_adresse[5]), .I2(n8), .O(n206) );
  NAND3_GATE U322 ( .I1(n208), .I2(n207), .I3(n206), .O(n495) );
  NAND_GATE U323 ( .I1(N88), .I2(n305), .O(n211) );
  NAND_GATE U324 ( .I1(N16), .I2(n306), .O(n210) );
  NAND_GATE U325 ( .I1(EX_adresse[6]), .I2(n8), .O(n209) );
  NAND3_GATE U326 ( .I1(n211), .I2(n210), .I3(n209), .O(n496) );
  NAND_GATE U327 ( .I1(N89), .I2(n305), .O(n214) );
  NAND_GATE U328 ( .I1(N17), .I2(n306), .O(n213) );
  NAND_GATE U329 ( .I1(EX_adresse[7]), .I2(n9), .O(n212) );
  NAND3_GATE U330 ( .I1(n214), .I2(n213), .I3(n212), .O(n497) );
  NAND_GATE U331 ( .I1(N90), .I2(n305), .O(n217) );
  NAND_GATE U332 ( .I1(N18), .I2(n306), .O(n216) );
  NAND_GATE U333 ( .I1(EX_adresse[8]), .I2(n9), .O(n215) );
  NAND3_GATE U334 ( .I1(n217), .I2(n216), .I3(n215), .O(n498) );
  NAND_GATE U335 ( .I1(N91), .I2(n305), .O(n220) );
  NAND_GATE U336 ( .I1(N19), .I2(n306), .O(n219) );
  NAND_GATE U337 ( .I1(EX_adresse[9]), .I2(n9), .O(n218) );
  NAND3_GATE U338 ( .I1(n220), .I2(n219), .I3(n218), .O(n499) );
  NAND_GATE U339 ( .I1(N92), .I2(n305), .O(n244) );
  NAND_GATE U340 ( .I1(N20), .I2(n306), .O(n243) );
  NAND_GATE U341 ( .I1(EX_adresse[10]), .I2(n9), .O(n242) );
  NAND3_GATE U342 ( .I1(n244), .I2(n243), .I3(n242), .O(n500) );
  NAND_GATE U343 ( .I1(N93), .I2(n305), .O(n247) );
  NAND_GATE U344 ( .I1(N21), .I2(n306), .O(n246) );
  NAND_GATE U345 ( .I1(EX_adresse[11]), .I2(n9), .O(n245) );
  NAND3_GATE U346 ( .I1(n247), .I2(n246), .I3(n245), .O(n501) );
  NAND_GATE U347 ( .I1(N94), .I2(n305), .O(n250) );
  NAND_GATE U348 ( .I1(N22), .I2(n306), .O(n249) );
  NAND_GATE U349 ( .I1(EX_adresse[12]), .I2(n9), .O(n248) );
  NAND3_GATE U350 ( .I1(n250), .I2(n249), .I3(n248), .O(n502) );
  NAND_GATE U351 ( .I1(N95), .I2(n305), .O(n253) );
  NAND_GATE U352 ( .I1(N23), .I2(n306), .O(n252) );
  NAND_GATE U353 ( .I1(EX_adresse[13]), .I2(n9), .O(n251) );
  NAND3_GATE U354 ( .I1(n253), .I2(n252), .I3(n251), .O(n503) );
  NAND_GATE U355 ( .I1(N96), .I2(n305), .O(n256) );
  NAND_GATE U356 ( .I1(N24), .I2(n306), .O(n255) );
  NAND_GATE U357 ( .I1(EX_adresse[14]), .I2(n9), .O(n254) );
  NAND3_GATE U358 ( .I1(n256), .I2(n255), .I3(n254), .O(n504) );
  NAND_GATE U359 ( .I1(N97), .I2(n305), .O(n259) );
  NAND_GATE U360 ( .I1(N25), .I2(n306), .O(n258) );
  NAND_GATE U361 ( .I1(EX_adresse[15]), .I2(n9), .O(n257) );
  NAND3_GATE U362 ( .I1(n259), .I2(n258), .I3(n257), .O(n505) );
  NAND_GATE U363 ( .I1(N98), .I2(n305), .O(n262) );
  NAND_GATE U364 ( .I1(N26), .I2(n306), .O(n261) );
  NAND_GATE U365 ( .I1(EX_adresse[16]), .I2(n10), .O(n260) );
  NAND3_GATE U366 ( .I1(n262), .I2(n261), .I3(n260), .O(n506) );
  NAND_GATE U367 ( .I1(N99), .I2(n305), .O(n265) );
  NAND_GATE U368 ( .I1(N27), .I2(n306), .O(n264) );
  NAND_GATE U369 ( .I1(EX_adresse[17]), .I2(n10), .O(n263) );
  NAND3_GATE U370 ( .I1(n265), .I2(n264), .I3(n263), .O(n507) );
  NAND_GATE U371 ( .I1(N100), .I2(n305), .O(n268) );
  NAND_GATE U372 ( .I1(N28), .I2(n306), .O(n267) );
  NAND_GATE U373 ( .I1(EX_adresse[18]), .I2(n10), .O(n266) );
  NAND3_GATE U374 ( .I1(n268), .I2(n267), .I3(n266), .O(n508) );
  NAND_GATE U375 ( .I1(N101), .I2(n305), .O(n271) );
  NAND_GATE U376 ( .I1(N29), .I2(n306), .O(n270) );
  NAND_GATE U377 ( .I1(EX_adresse[19]), .I2(n10), .O(n269) );
  NAND3_GATE U378 ( .I1(n271), .I2(n270), .I3(n269), .O(n509) );
  NAND_GATE U379 ( .I1(N102), .I2(n305), .O(n274) );
  NAND_GATE U380 ( .I1(N30), .I2(n306), .O(n273) );
  NAND_GATE U381 ( .I1(EX_adresse[20]), .I2(n10), .O(n272) );
  NAND3_GATE U382 ( .I1(n274), .I2(n273), .I3(n272), .O(n510) );
  NAND_GATE U383 ( .I1(N103), .I2(n305), .O(n277) );
  NAND_GATE U384 ( .I1(N31), .I2(n306), .O(n276) );
  NAND_GATE U385 ( .I1(EX_adresse[21]), .I2(n10), .O(n275) );
  NAND3_GATE U386 ( .I1(n277), .I2(n276), .I3(n275), .O(n511) );
  NAND_GATE U387 ( .I1(N104), .I2(n305), .O(n280) );
  NAND_GATE U388 ( .I1(N32), .I2(n306), .O(n279) );
  NAND_GATE U389 ( .I1(EX_adresse[22]), .I2(n10), .O(n278) );
  NAND3_GATE U390 ( .I1(n280), .I2(n279), .I3(n278), .O(n512) );
  NAND_GATE U391 ( .I1(N105), .I2(n305), .O(n283) );
  NAND_GATE U392 ( .I1(N33), .I2(n306), .O(n282) );
  NAND_GATE U393 ( .I1(EX_adresse[23]), .I2(n10), .O(n281) );
  NAND3_GATE U394 ( .I1(n283), .I2(n282), .I3(n281), .O(n513) );
  NAND_GATE U395 ( .I1(N106), .I2(n305), .O(n286) );
  NAND_GATE U396 ( .I1(N34), .I2(n306), .O(n285) );
  NAND_GATE U397 ( .I1(EX_adresse[24]), .I2(n10), .O(n284) );
  NAND3_GATE U398 ( .I1(n286), .I2(n285), .I3(n284), .O(n514) );
  NAND_GATE U399 ( .I1(N107), .I2(n305), .O(n289) );
  NAND_GATE U400 ( .I1(N35), .I2(n306), .O(n288) );
  NAND_GATE U401 ( .I1(EX_adresse[25]), .I2(n11), .O(n287) );
  NAND3_GATE U402 ( .I1(n289), .I2(n288), .I3(n287), .O(n515) );
  NAND_GATE U403 ( .I1(N108), .I2(n305), .O(n292) );
  NAND_GATE U404 ( .I1(N36), .I2(n306), .O(n291) );
  NAND_GATE U405 ( .I1(EX_adresse[26]), .I2(n11), .O(n290) );
  NAND3_GATE U406 ( .I1(n292), .I2(n291), .I3(n290), .O(n516) );
  NAND_GATE U407 ( .I1(N109), .I2(n305), .O(n295) );
  NAND_GATE U408 ( .I1(N37), .I2(n306), .O(n294) );
  NAND_GATE U409 ( .I1(EX_adresse[27]), .I2(n11), .O(n293) );
  NAND3_GATE U410 ( .I1(n295), .I2(n294), .I3(n293), .O(n517) );
  NAND_GATE U411 ( .I1(N110), .I2(n305), .O(n298) );
  NAND_GATE U412 ( .I1(N38), .I2(n306), .O(n297) );
  NAND_GATE U413 ( .I1(EX_adresse[28]), .I2(n11), .O(n296) );
  NAND3_GATE U414 ( .I1(n298), .I2(n297), .I3(n296), .O(n518) );
  NAND_GATE U415 ( .I1(N111), .I2(n305), .O(n301) );
  NAND_GATE U416 ( .I1(N39), .I2(n306), .O(n300) );
  NAND_GATE U417 ( .I1(EX_adresse[29]), .I2(n11), .O(n299) );
  NAND3_GATE U418 ( .I1(n301), .I2(n300), .I3(n299), .O(n519) );
  NAND_GATE U419 ( .I1(N112), .I2(n305), .O(n304) );
  NAND_GATE U518 ( .I1(N40), .I2(n306), .O(n303) );
  NAND_GATE U519 ( .I1(EX_adresse[30]), .I2(n11), .O(n302) );
  NAND3_GATE U521 ( .I1(n304), .I2(n303), .I3(n302), .O(n520) );
  NAND_GATE U522 ( .I1(N113), .I2(n305), .O(n309) );
  NAND_GATE U523 ( .I1(N41), .I2(n306), .O(n308) );
  NAND_GATE U524 ( .I1(EX_adresse[31]), .I2(n11), .O(n307) );
  NAND3_GATE U525 ( .I1(n309), .I2(n308), .I3(n307), .O(n521) );
  NAND_GATE U526 ( .I1(res_ual[0]), .I2(n2), .O(n312) );
  NAND_GATE U527 ( .I1(N10), .I2(n1), .O(n311) );
  NAND_GATE U528 ( .I1(EX_data_ual[0]), .I2(n11), .O(n310) );
  NAND3_GATE U529 ( .I1(n312), .I2(n311), .I3(n310), .O(n522) );
  NAND_GATE U530 ( .I1(res_ual[8]), .I2(n2), .O(n315) );
  NAND_GATE U531 ( .I1(N18), .I2(n1), .O(n314) );
  NAND_GATE U532 ( .I1(EX_data_ual[8]), .I2(n11), .O(n313) );
  NAND3_GATE U533 ( .I1(n315), .I2(n314), .I3(n313), .O(n530) );
  NAND_GATE U534 ( .I1(res_ual[9]), .I2(n2), .O(n384) );
  NAND_GATE U535 ( .I1(N19), .I2(n1), .O(n383) );
  NAND_GATE U536 ( .I1(EX_data_ual[9]), .I2(n8), .O(n380) );
  NAND3_GATE U537 ( .I1(n384), .I2(n383), .I3(n380), .O(n531) );
  NAND_GATE U538 ( .I1(res_ual[10]), .I2(n2), .O(n387) );
  NAND_GATE U539 ( .I1(N20), .I2(n1), .O(n386) );
  NAND_GATE U540 ( .I1(EX_data_ual[10]), .I2(n594), .O(n385) );
  NAND3_GATE U541 ( .I1(n387), .I2(n386), .I3(n385), .O(n532) );
  NAND_GATE U542 ( .I1(res_ual[11]), .I2(n2), .O(n390) );
  NAND_GATE U543 ( .I1(N21), .I2(n1), .O(n389) );
  NAND_GATE U544 ( .I1(EX_data_ual[11]), .I2(n11), .O(n388) );
  NAND3_GATE U545 ( .I1(n390), .I2(n389), .I3(n388), .O(n533) );
  NAND_GATE U546 ( .I1(res_ual[12]), .I2(n2), .O(n393) );
  NAND_GATE U547 ( .I1(N22), .I2(n1), .O(n392) );
  NAND_GATE U548 ( .I1(EX_data_ual[12]), .I2(n10), .O(n391) );
  NAND3_GATE U549 ( .I1(n393), .I2(n392), .I3(n391), .O(n534) );
  NAND_GATE U550 ( .I1(res_ual[13]), .I2(n2), .O(n396) );
  NAND_GATE U551 ( .I1(N23), .I2(n1), .O(n395) );
  NAND_GATE U552 ( .I1(EX_data_ual[13]), .I2(n9), .O(n394) );
  NAND3_GATE U553 ( .I1(n396), .I2(n395), .I3(n394), .O(n535) );
  NAND_GATE U554 ( .I1(res_ual[14]), .I2(n2), .O(n399) );
  NAND_GATE U555 ( .I1(N24), .I2(n1), .O(n398) );
  NAND_GATE U556 ( .I1(EX_data_ual[14]), .I2(n8), .O(n397) );
  NAND3_GATE U557 ( .I1(n399), .I2(n398), .I3(n397), .O(n536) );
  NAND_GATE U558 ( .I1(res_ual[15]), .I2(n2), .O(n402) );
  NAND_GATE U559 ( .I1(N25), .I2(n1), .O(n401) );
  NAND_GATE U560 ( .I1(EX_data_ual[15]), .I2(n594), .O(n400) );
  NAND3_GATE U561 ( .I1(n402), .I2(n401), .I3(n400), .O(n537) );
  NAND_GATE U562 ( .I1(res_ual[16]), .I2(n2), .O(n405) );
  NAND_GATE U563 ( .I1(N26), .I2(n1), .O(n404) );
  NAND_GATE U564 ( .I1(EX_data_ual[16]), .I2(n11), .O(n403) );
  NAND3_GATE U565 ( .I1(n405), .I2(n404), .I3(n403), .O(n538) );
  NAND_GATE U566 ( .I1(res_ual[17]), .I2(n2), .O(n408) );
  NAND_GATE U567 ( .I1(N27), .I2(n1), .O(n407) );
  NAND_GATE U568 ( .I1(EX_data_ual[17]), .I2(n10), .O(n406) );
  NAND3_GATE U569 ( .I1(n408), .I2(n407), .I3(n406), .O(n539) );
  NAND_GATE U570 ( .I1(res_ual[18]), .I2(n2), .O(n411) );
  NAND_GATE U571 ( .I1(N28), .I2(n1), .O(n410) );
  NAND_GATE U572 ( .I1(EX_data_ual[18]), .I2(n594), .O(n409) );
  NAND3_GATE U573 ( .I1(n411), .I2(n410), .I3(n409), .O(n540) );
  NAND_GATE U574 ( .I1(res_ual[19]), .I2(n2), .O(n414) );
  NAND_GATE U575 ( .I1(N29), .I2(n1), .O(n413) );
  NAND_GATE U576 ( .I1(EX_data_ual[19]), .I2(n9), .O(n412) );
  NAND3_GATE U577 ( .I1(n414), .I2(n413), .I3(n412), .O(n541) );
  NAND_GATE U578 ( .I1(res_ual[20]), .I2(n2), .O(n417) );
  NAND_GATE U579 ( .I1(N30), .I2(n1), .O(n416) );
  NAND_GATE U580 ( .I1(EX_data_ual[20]), .I2(n11), .O(n415) );
  NAND3_GATE U581 ( .I1(n417), .I2(n416), .I3(n415), .O(n542) );
  NAND_GATE U582 ( .I1(res_ual[21]), .I2(n2), .O(n420) );
  NAND_GATE U583 ( .I1(N31), .I2(n1), .O(n419) );
  NAND_GATE U584 ( .I1(EX_data_ual[21]), .I2(n10), .O(n418) );
  NAND3_GATE U585 ( .I1(n420), .I2(n419), .I3(n418), .O(n543) );
  NAND_GATE U586 ( .I1(res_ual[22]), .I2(n2), .O(n423) );
  NAND_GATE U587 ( .I1(N32), .I2(n1), .O(n422) );
  NAND_GATE U588 ( .I1(EX_data_ual[22]), .I2(n9), .O(n421) );
  NAND3_GATE U589 ( .I1(n423), .I2(n422), .I3(n421), .O(n544) );
  NAND_GATE U590 ( .I1(res_ual[23]), .I2(n2), .O(n426) );
  NAND_GATE U591 ( .I1(N33), .I2(n1), .O(n425) );
  NAND_GATE U592 ( .I1(EX_data_ual[23]), .I2(n8), .O(n424) );
  NAND3_GATE U593 ( .I1(n426), .I2(n425), .I3(n424), .O(n545) );
  NAND_GATE U594 ( .I1(res_ual[24]), .I2(n2), .O(n429) );
  NAND_GATE U595 ( .I1(N34), .I2(n1), .O(n428) );
  NAND_GATE U596 ( .I1(EX_data_ual[24]), .I2(n594), .O(n427) );
  NAND3_GATE U597 ( .I1(n429), .I2(n428), .I3(n427), .O(n546) );
  NAND_GATE U598 ( .I1(res_ual[25]), .I2(n2), .O(n432) );
  NAND_GATE U599 ( .I1(N35), .I2(n1), .O(n431) );
  NAND_GATE U600 ( .I1(EX_data_ual[25]), .I2(n8), .O(n430) );
  NAND3_GATE U601 ( .I1(n432), .I2(n431), .I3(n430), .O(n547) );
  NAND_GATE U602 ( .I1(res_ual[26]), .I2(n2), .O(n435) );
  NAND_GATE U603 ( .I1(N36), .I2(n1), .O(n434) );
  NAND_GATE U604 ( .I1(EX_data_ual[26]), .I2(n11), .O(n433) );
  NAND3_GATE U605 ( .I1(n435), .I2(n434), .I3(n433), .O(n548) );
  NAND_GATE U606 ( .I1(res_ual[27]), .I2(n2), .O(n438) );
  NAND_GATE U607 ( .I1(N37), .I2(n1), .O(n437) );
  NAND_GATE U608 ( .I1(EX_data_ual[27]), .I2(n594), .O(n436) );
  NAND3_GATE U609 ( .I1(n438), .I2(n437), .I3(n436), .O(n549) );
  NAND_GATE U610 ( .I1(res_ual[28]), .I2(n2), .O(n441) );
  NAND_GATE U611 ( .I1(N38), .I2(n1), .O(n440) );
  NAND_GATE U612 ( .I1(EX_data_ual[28]), .I2(n594), .O(n439) );
  NAND3_GATE U613 ( .I1(n441), .I2(n440), .I3(n439), .O(n550) );
  NAND_GATE U614 ( .I1(res_ual[29]), .I2(n2), .O(n444) );
  NAND_GATE U615 ( .I1(N39), .I2(n1), .O(n443) );
  NAND_GATE U616 ( .I1(EX_data_ual[29]), .I2(n594), .O(n442) );
  NAND3_GATE U617 ( .I1(n444), .I2(n443), .I3(n442), .O(n551) );
  NAND_GATE U618 ( .I1(res_ual[30]), .I2(n2), .O(n588) );
  NAND_GATE U619 ( .I1(N40), .I2(n1), .O(n446) );
  NAND_GATE U620 ( .I1(EX_data_ual[30]), .I2(n594), .O(n445) );
  NAND3_GATE U621 ( .I1(n588), .I2(n446), .I3(n445), .O(n552) );
  NAND_GATE U622 ( .I1(res_ual[31]), .I2(n2), .O(n591) );
  NAND_GATE U623 ( .I1(N41), .I2(n1), .O(n590) );
  NAND_GATE U624 ( .I1(EX_data_ual[31]), .I2(n594), .O(n589) );
  NAND3_GATE U625 ( .I1(n591), .I2(n590), .I3(n589), .O(n553) );
  NAND_GATE U626 ( .I1(EX_bra_confirm), .I2(n12), .O(n593) );
  NAND_GATE U627 ( .I1(n4), .I2(n7), .O(n592) );
  NAND_GATE U628 ( .I1(n593), .I2(n592), .O(n554) );
endmodule


module pps_di ( clock, reset, stop_all, clear, adr_reg1, adr_reg2, use1, use2, 
        stop_di, data1, data2, EI_adr, EI_instr, EI_it_ok, DI_bra, DI_link, 
        DI_op1, DI_op2, DI_code_ual, DI_offset, DI_adr_reg_dest, DI_ecr_reg, 
        DI_mode, DI_op_mem, DI_r_w, DI_adr, DI_exc_cause, DI_level, DI_it_ok
 );
  output [5:0] adr_reg1;
  output [5:0] adr_reg2;
  input [31:0] data1;
  input [31:0] data2;
  input [31:0] EI_adr;
  input [31:0] EI_instr;
  output [31:0] DI_op1;
  output [31:0] DI_op2;
  output [27:0] DI_code_ual;
  output [31:0] DI_offset;
  output [5:0] DI_adr_reg_dest;
  output [31:0] DI_adr;
  output [31:0] DI_exc_cause;
  output [1:0] DI_level;
  input clock, reset, stop_all, clear, stop_di, EI_it_ok;
  output use1, use2, DI_bra, DI_link, DI_ecr_reg, DI_mode, DI_op_mem, DI_r_w,
         DI_it_ok;
  wire   n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958;
  assign adr_reg1[5] = 1'b0;

  FLIP_FLOP_D DI_it_ok_reg ( .D(n942), .CK(clock), .Q(DI_it_ok) );
  FLIP_FLOP_D DI_bra_reg ( .D(n941), .CK(clock), .Q(DI_bra) );
  FLIP_FLOP_D DI_link_reg ( .D(n940), .CK(clock), .Q(DI_link) );
  FLIP_FLOP_D \DI_op1_reg[31]  ( .D(n939), .CK(clock), .Q(DI_op1[31]) );
  FLIP_FLOP_D \DI_op1_reg[30]  ( .D(n938), .CK(clock), .Q(DI_op1[30]) );
  FLIP_FLOP_D \DI_op1_reg[29]  ( .D(n937), .CK(clock), .Q(DI_op1[29]) );
  FLIP_FLOP_D \DI_op1_reg[28]  ( .D(n936), .CK(clock), .Q(DI_op1[28]) );
  FLIP_FLOP_D \DI_op1_reg[27]  ( .D(n935), .CK(clock), .Q(DI_op1[27]) );
  FLIP_FLOP_D \DI_op1_reg[26]  ( .D(n934), .CK(clock), .Q(DI_op1[26]) );
  FLIP_FLOP_D \DI_op1_reg[25]  ( .D(n933), .CK(clock), .Q(DI_op1[25]) );
  FLIP_FLOP_D \DI_op1_reg[24]  ( .D(n932), .CK(clock), .Q(DI_op1[24]) );
  FLIP_FLOP_D \DI_op1_reg[23]  ( .D(n931), .CK(clock), .Q(DI_op1[23]) );
  FLIP_FLOP_D \DI_op1_reg[22]  ( .D(n930), .CK(clock), .Q(DI_op1[22]) );
  FLIP_FLOP_D \DI_op1_reg[21]  ( .D(n929), .CK(clock), .Q(DI_op1[21]) );
  FLIP_FLOP_D \DI_op1_reg[20]  ( .D(n928), .CK(clock), .Q(DI_op1[20]) );
  FLIP_FLOP_D \DI_op1_reg[19]  ( .D(n927), .CK(clock), .Q(DI_op1[19]) );
  FLIP_FLOP_D \DI_op1_reg[18]  ( .D(n926), .CK(clock), .Q(DI_op1[18]) );
  FLIP_FLOP_D \DI_op1_reg[17]  ( .D(n925), .CK(clock), .Q(DI_op1[17]) );
  FLIP_FLOP_D \DI_op1_reg[16]  ( .D(n924), .CK(clock), .Q(DI_op1[16]) );
  FLIP_FLOP_D \DI_op1_reg[15]  ( .D(n923), .CK(clock), .Q(DI_op1[15]) );
  FLIP_FLOP_D \DI_op1_reg[14]  ( .D(n922), .CK(clock), .Q(DI_op1[14]) );
  FLIP_FLOP_D \DI_op1_reg[13]  ( .D(n921), .CK(clock), .Q(DI_op1[13]) );
  FLIP_FLOP_D \DI_op1_reg[12]  ( .D(n920), .CK(clock), .Q(DI_op1[12]) );
  FLIP_FLOP_D \DI_op1_reg[11]  ( .D(n919), .CK(clock), .Q(DI_op1[11]) );
  FLIP_FLOP_D \DI_op1_reg[10]  ( .D(n918), .CK(clock), .Q(DI_op1[10]) );
  FLIP_FLOP_D \DI_op1_reg[9]  ( .D(n917), .CK(clock), .Q(DI_op1[9]) );
  FLIP_FLOP_D \DI_op1_reg[8]  ( .D(n916), .CK(clock), .Q(DI_op1[8]) );
  FLIP_FLOP_D \DI_op1_reg[7]  ( .D(n915), .CK(clock), .Q(DI_op1[7]) );
  FLIP_FLOP_D \DI_op1_reg[6]  ( .D(n914), .CK(clock), .Q(DI_op1[6]) );
  FLIP_FLOP_D \DI_op1_reg[5]  ( .D(n913), .CK(clock), .Q(DI_op1[5]) );
  FLIP_FLOP_D \DI_op1_reg[4]  ( .D(n912), .CK(clock), .Q(DI_op1[4]) );
  FLIP_FLOP_D \DI_op1_reg[3]  ( .D(n911), .CK(clock), .Q(DI_op1[3]) );
  FLIP_FLOP_D \DI_op1_reg[2]  ( .D(n910), .CK(clock), .Q(DI_op1[2]) );
  FLIP_FLOP_D \DI_op1_reg[1]  ( .D(n909), .CK(clock), .Q(DI_op1[1]) );
  FLIP_FLOP_D \DI_op1_reg[0]  ( .D(n908), .CK(clock), .Q(DI_op1[0]) );
  FLIP_FLOP_D \DI_op2_reg[31]  ( .D(n907), .CK(clock), .Q(DI_op2[31]) );
  FLIP_FLOP_D \DI_op2_reg[30]  ( .D(n906), .CK(clock), .Q(DI_op2[30]) );
  FLIP_FLOP_D \DI_op2_reg[29]  ( .D(n905), .CK(clock), .Q(DI_op2[29]) );
  FLIP_FLOP_D \DI_op2_reg[28]  ( .D(n904), .CK(clock), .Q(DI_op2[28]) );
  FLIP_FLOP_D \DI_op2_reg[27]  ( .D(n903), .CK(clock), .Q(DI_op2[27]) );
  FLIP_FLOP_D \DI_op2_reg[26]  ( .D(n902), .CK(clock), .Q(DI_op2[26]) );
  FLIP_FLOP_D \DI_op2_reg[25]  ( .D(n901), .CK(clock), .Q(DI_op2[25]) );
  FLIP_FLOP_D \DI_op2_reg[24]  ( .D(n900), .CK(clock), .Q(DI_op2[24]) );
  FLIP_FLOP_D \DI_op2_reg[23]  ( .D(n899), .CK(clock), .Q(DI_op2[23]) );
  FLIP_FLOP_D \DI_op2_reg[22]  ( .D(n898), .CK(clock), .Q(DI_op2[22]) );
  FLIP_FLOP_D \DI_op2_reg[21]  ( .D(n897), .CK(clock), .Q(DI_op2[21]) );
  FLIP_FLOP_D \DI_op2_reg[20]  ( .D(n896), .CK(clock), .Q(DI_op2[20]) );
  FLIP_FLOP_D \DI_op2_reg[19]  ( .D(n895), .CK(clock), .Q(DI_op2[19]) );
  FLIP_FLOP_D \DI_op2_reg[18]  ( .D(n894), .CK(clock), .Q(DI_op2[18]) );
  FLIP_FLOP_D \DI_op2_reg[17]  ( .D(n893), .CK(clock), .Q(DI_op2[17]) );
  FLIP_FLOP_D \DI_op2_reg[16]  ( .D(n892), .CK(clock), .Q(DI_op2[16]) );
  FLIP_FLOP_D \DI_op2_reg[15]  ( .D(n891), .CK(clock), .Q(DI_op2[15]) );
  FLIP_FLOP_D \DI_op2_reg[14]  ( .D(n890), .CK(clock), .Q(DI_op2[14]) );
  FLIP_FLOP_D \DI_op2_reg[13]  ( .D(n889), .CK(clock), .Q(DI_op2[13]) );
  FLIP_FLOP_D \DI_op2_reg[12]  ( .D(n888), .CK(clock), .Q(DI_op2[12]) );
  FLIP_FLOP_D \DI_op2_reg[11]  ( .D(n887), .CK(clock), .Q(DI_op2[11]) );
  FLIP_FLOP_D \DI_op2_reg[10]  ( .D(n886), .CK(clock), .Q(DI_op2[10]) );
  FLIP_FLOP_D \DI_op2_reg[9]  ( .D(n885), .CK(clock), .Q(DI_op2[9]) );
  FLIP_FLOP_D \DI_op2_reg[8]  ( .D(n884), .CK(clock), .Q(DI_op2[8]) );
  FLIP_FLOP_D \DI_op2_reg[7]  ( .D(n883), .CK(clock), .Q(DI_op2[7]) );
  FLIP_FLOP_D \DI_op2_reg[6]  ( .D(n882), .CK(clock), .Q(DI_op2[6]) );
  FLIP_FLOP_D \DI_op2_reg[5]  ( .D(n881), .CK(clock), .Q(DI_op2[5]) );
  FLIP_FLOP_D \DI_op2_reg[4]  ( .D(n880), .CK(clock), .Q(DI_op2[4]) );
  FLIP_FLOP_D \DI_op2_reg[3]  ( .D(n879), .CK(clock), .Q(DI_op2[3]) );
  FLIP_FLOP_D \DI_op2_reg[2]  ( .D(n878), .CK(clock), .Q(DI_op2[2]) );
  FLIP_FLOP_D \DI_op2_reg[1]  ( .D(n877), .CK(clock), .Q(DI_op2[1]) );
  FLIP_FLOP_D \DI_op2_reg[0]  ( .D(n876), .CK(clock), .Q(DI_op2[0]) );
  FLIP_FLOP_D \DI_code_ual_reg[27]  ( .D(n875), .CK(clock), .Q(DI_code_ual[27]) );
  FLIP_FLOP_D \DI_code_ual_reg[26]  ( .D(n874), .CK(clock), .Q(DI_code_ual[26]) );
  FLIP_FLOP_D \DI_code_ual_reg[25]  ( .D(n873), .CK(clock), .Q(DI_code_ual[25]) );
  FLIP_FLOP_D \DI_code_ual_reg[24]  ( .D(n872), .CK(clock), .Q(DI_code_ual[24]) );
  FLIP_FLOP_D \DI_code_ual_reg[23]  ( .D(n871), .CK(clock), .Q(DI_code_ual[23]) );
  FLIP_FLOP_D \DI_code_ual_reg[22]  ( .D(n870), .CK(clock), .Q(DI_code_ual[22]) );
  FLIP_FLOP_D \DI_code_ual_reg[21]  ( .D(n869), .CK(clock), .Q(DI_code_ual[21]) );
  FLIP_FLOP_D \DI_code_ual_reg[20]  ( .D(n868), .CK(clock), .Q(DI_code_ual[20]) );
  FLIP_FLOP_D \DI_code_ual_reg[19]  ( .D(n867), .CK(clock), .Q(DI_code_ual[19]) );
  FLIP_FLOP_D \DI_code_ual_reg[18]  ( .D(n866), .CK(clock), .Q(DI_code_ual[18]) );
  FLIP_FLOP_D \DI_code_ual_reg[17]  ( .D(n865), .CK(clock), .Q(DI_code_ual[17]) );
  FLIP_FLOP_D \DI_code_ual_reg[16]  ( .D(n864), .CK(clock), .Q(DI_code_ual[16]) );
  FLIP_FLOP_D \DI_code_ual_reg[15]  ( .D(n863), .CK(clock), .Q(DI_code_ual[15]) );
  FLIP_FLOP_D \DI_code_ual_reg[14]  ( .D(n862), .CK(clock), .Q(DI_code_ual[14]) );
  FLIP_FLOP_D \DI_code_ual_reg[13]  ( .D(n861), .CK(clock), .Q(DI_code_ual[13]) );
  FLIP_FLOP_D \DI_code_ual_reg[12]  ( .D(n860), .CK(clock), .Q(DI_code_ual[12]) );
  FLIP_FLOP_D \DI_code_ual_reg[11]  ( .D(n859), .CK(clock), .Q(DI_code_ual[11]) );
  FLIP_FLOP_D \DI_code_ual_reg[10]  ( .D(n858), .CK(clock), .Q(DI_code_ual[10]) );
  FLIP_FLOP_D \DI_code_ual_reg[9]  ( .D(n857), .CK(clock), .Q(DI_code_ual[9])
         );
  FLIP_FLOP_D \DI_code_ual_reg[8]  ( .D(n856), .CK(clock), .Q(DI_code_ual[8])
         );
  FLIP_FLOP_D \DI_code_ual_reg[7]  ( .D(n855), .CK(clock), .Q(DI_code_ual[7])
         );
  FLIP_FLOP_D \DI_code_ual_reg[6]  ( .D(n854), .CK(clock), .Q(DI_code_ual[6])
         );
  FLIP_FLOP_D \DI_code_ual_reg[5]  ( .D(n853), .CK(clock), .Q(DI_code_ual[5])
         );
  FLIP_FLOP_D \DI_code_ual_reg[4]  ( .D(n852), .CK(clock), .Q(DI_code_ual[4])
         );
  FLIP_FLOP_D \DI_code_ual_reg[3]  ( .D(n851), .CK(clock), .Q(DI_code_ual[3])
         );
  FLIP_FLOP_D \DI_code_ual_reg[2]  ( .D(n850), .CK(clock), .Q(DI_code_ual[2])
         );
  FLIP_FLOP_D \DI_code_ual_reg[1]  ( .D(n849), .CK(clock), .Q(DI_code_ual[1])
         );
  FLIP_FLOP_D \DI_code_ual_reg[0]  ( .D(n848), .CK(clock), .Q(DI_code_ual[0])
         );
  FLIP_FLOP_D \DI_offset_reg[31]  ( .D(n847), .CK(clock), .Q(DI_offset[31]) );
  FLIP_FLOP_D \DI_offset_reg[30]  ( .D(n846), .CK(clock), .Q(DI_offset[30]) );
  FLIP_FLOP_D \DI_offset_reg[29]  ( .D(n845), .CK(clock), .Q(DI_offset[29]) );
  FLIP_FLOP_D \DI_offset_reg[28]  ( .D(n844), .CK(clock), .Q(DI_offset[28]) );
  FLIP_FLOP_D \DI_offset_reg[27]  ( .D(n843), .CK(clock), .Q(DI_offset[27]) );
  FLIP_FLOP_D \DI_offset_reg[26]  ( .D(n842), .CK(clock), .Q(DI_offset[26]) );
  FLIP_FLOP_D \DI_offset_reg[25]  ( .D(n841), .CK(clock), .Q(DI_offset[25]) );
  FLIP_FLOP_D \DI_offset_reg[24]  ( .D(n840), .CK(clock), .Q(DI_offset[24]) );
  FLIP_FLOP_D \DI_offset_reg[23]  ( .D(n839), .CK(clock), .Q(DI_offset[23]) );
  FLIP_FLOP_D \DI_offset_reg[22]  ( .D(n838), .CK(clock), .Q(DI_offset[22]) );
  FLIP_FLOP_D \DI_offset_reg[21]  ( .D(n837), .CK(clock), .Q(DI_offset[21]) );
  FLIP_FLOP_D \DI_offset_reg[20]  ( .D(n836), .CK(clock), .Q(DI_offset[20]) );
  FLIP_FLOP_D \DI_offset_reg[19]  ( .D(n835), .CK(clock), .Q(DI_offset[19]) );
  FLIP_FLOP_D \DI_offset_reg[18]  ( .D(n834), .CK(clock), .Q(DI_offset[18]) );
  FLIP_FLOP_D \DI_offset_reg[17]  ( .D(n833), .CK(clock), .Q(DI_offset[17]) );
  FLIP_FLOP_D \DI_offset_reg[16]  ( .D(n832), .CK(clock), .Q(DI_offset[16]) );
  FLIP_FLOP_D \DI_offset_reg[15]  ( .D(n831), .CK(clock), .Q(DI_offset[15]) );
  FLIP_FLOP_D \DI_offset_reg[14]  ( .D(n830), .CK(clock), .Q(DI_offset[14]) );
  FLIP_FLOP_D \DI_offset_reg[13]  ( .D(n829), .CK(clock), .Q(DI_offset[13]) );
  FLIP_FLOP_D \DI_offset_reg[12]  ( .D(n828), .CK(clock), .Q(DI_offset[12]) );
  FLIP_FLOP_D \DI_offset_reg[11]  ( .D(n827), .CK(clock), .Q(DI_offset[11]) );
  FLIP_FLOP_D \DI_offset_reg[10]  ( .D(n826), .CK(clock), .Q(DI_offset[10]) );
  FLIP_FLOP_D \DI_offset_reg[9]  ( .D(n825), .CK(clock), .Q(DI_offset[9]) );
  FLIP_FLOP_D \DI_offset_reg[8]  ( .D(n824), .CK(clock), .Q(DI_offset[8]) );
  FLIP_FLOP_D \DI_offset_reg[7]  ( .D(n823), .CK(clock), .Q(DI_offset[7]) );
  FLIP_FLOP_D \DI_offset_reg[6]  ( .D(n822), .CK(clock), .Q(DI_offset[6]) );
  FLIP_FLOP_D \DI_offset_reg[5]  ( .D(n821), .CK(clock), .Q(DI_offset[5]) );
  FLIP_FLOP_D \DI_offset_reg[4]  ( .D(n820), .CK(clock), .Q(DI_offset[4]) );
  FLIP_FLOP_D \DI_offset_reg[3]  ( .D(n819), .CK(clock), .Q(DI_offset[3]) );
  FLIP_FLOP_D \DI_offset_reg[2]  ( .D(n818), .CK(clock), .Q(DI_offset[2]) );
  FLIP_FLOP_D \DI_offset_reg[1]  ( .D(n817), .CK(clock), .Q(DI_offset[1]) );
  FLIP_FLOP_D \DI_offset_reg[0]  ( .D(n816), .CK(clock), .Q(DI_offset[0]) );
  FLIP_FLOP_D \DI_adr_reg_dest_reg[5]  ( .D(n815), .CK(clock), .Q(
        DI_adr_reg_dest[5]) );
  FLIP_FLOP_D \DI_adr_reg_dest_reg[4]  ( .D(n814), .CK(clock), .Q(
        DI_adr_reg_dest[4]) );
  FLIP_FLOP_D \DI_adr_reg_dest_reg[3]  ( .D(n813), .CK(clock), .Q(
        DI_adr_reg_dest[3]) );
  FLIP_FLOP_D \DI_adr_reg_dest_reg[2]  ( .D(n812), .CK(clock), .Q(
        DI_adr_reg_dest[2]) );
  FLIP_FLOP_D \DI_adr_reg_dest_reg[1]  ( .D(n811), .CK(clock), .Q(
        DI_adr_reg_dest[1]) );
  FLIP_FLOP_D \DI_adr_reg_dest_reg[0]  ( .D(n810), .CK(clock), .Q(
        DI_adr_reg_dest[0]) );
  FLIP_FLOP_D DI_ecr_reg_reg ( .D(n809), .CK(clock), .Q(DI_ecr_reg) );
  FLIP_FLOP_D DI_mode_reg ( .D(n808), .CK(clock), .Q(DI_mode) );
  FLIP_FLOP_D DI_op_mem_reg ( .D(n807), .CK(clock), .Q(DI_op_mem) );
  FLIP_FLOP_D DI_r_w_reg ( .D(n806), .CK(clock), .Q(DI_r_w) );
  FLIP_FLOP_D \DI_adr_reg[31]  ( .D(n805), .CK(clock), .Q(DI_adr[31]) );
  FLIP_FLOP_D \DI_adr_reg[30]  ( .D(n804), .CK(clock), .Q(DI_adr[30]) );
  FLIP_FLOP_D \DI_adr_reg[29]  ( .D(n803), .CK(clock), .Q(DI_adr[29]) );
  FLIP_FLOP_D \DI_adr_reg[28]  ( .D(n802), .CK(clock), .Q(DI_adr[28]) );
  FLIP_FLOP_D \DI_adr_reg[27]  ( .D(n801), .CK(clock), .Q(DI_adr[27]) );
  FLIP_FLOP_D \DI_adr_reg[26]  ( .D(n800), .CK(clock), .Q(DI_adr[26]) );
  FLIP_FLOP_D \DI_adr_reg[25]  ( .D(n799), .CK(clock), .Q(DI_adr[25]) );
  FLIP_FLOP_D \DI_adr_reg[24]  ( .D(n798), .CK(clock), .Q(DI_adr[24]) );
  FLIP_FLOP_D \DI_adr_reg[23]  ( .D(n797), .CK(clock), .Q(DI_adr[23]) );
  FLIP_FLOP_D \DI_adr_reg[22]  ( .D(n796), .CK(clock), .Q(DI_adr[22]) );
  FLIP_FLOP_D \DI_adr_reg[21]  ( .D(n795), .CK(clock), .Q(DI_adr[21]) );
  FLIP_FLOP_D \DI_adr_reg[20]  ( .D(n794), .CK(clock), .Q(DI_adr[20]) );
  FLIP_FLOP_D \DI_adr_reg[19]  ( .D(n793), .CK(clock), .Q(DI_adr[19]) );
  FLIP_FLOP_D \DI_adr_reg[18]  ( .D(n792), .CK(clock), .Q(DI_adr[18]) );
  FLIP_FLOP_D \DI_adr_reg[17]  ( .D(n791), .CK(clock), .Q(DI_adr[17]) );
  FLIP_FLOP_D \DI_adr_reg[16]  ( .D(n790), .CK(clock), .Q(DI_adr[16]) );
  FLIP_FLOP_D \DI_adr_reg[15]  ( .D(n789), .CK(clock), .Q(DI_adr[15]) );
  FLIP_FLOP_D \DI_adr_reg[14]  ( .D(n788), .CK(clock), .Q(DI_adr[14]) );
  FLIP_FLOP_D \DI_adr_reg[13]  ( .D(n787), .CK(clock), .Q(DI_adr[13]) );
  FLIP_FLOP_D \DI_adr_reg[12]  ( .D(n786), .CK(clock), .Q(DI_adr[12]) );
  FLIP_FLOP_D \DI_adr_reg[11]  ( .D(n785), .CK(clock), .Q(DI_adr[11]) );
  FLIP_FLOP_D \DI_adr_reg[10]  ( .D(n784), .CK(clock), .Q(DI_adr[10]) );
  FLIP_FLOP_D \DI_adr_reg[9]  ( .D(n783), .CK(clock), .Q(DI_adr[9]) );
  FLIP_FLOP_D \DI_adr_reg[8]  ( .D(n782), .CK(clock), .Q(DI_adr[8]) );
  FLIP_FLOP_D \DI_adr_reg[7]  ( .D(n781), .CK(clock), .Q(DI_adr[7]) );
  FLIP_FLOP_D \DI_adr_reg[6]  ( .D(n780), .CK(clock), .Q(DI_adr[6]) );
  FLIP_FLOP_D \DI_adr_reg[5]  ( .D(n779), .CK(clock), .Q(DI_adr[5]) );
  FLIP_FLOP_D \DI_adr_reg[4]  ( .D(n778), .CK(clock), .Q(DI_adr[4]) );
  FLIP_FLOP_D \DI_adr_reg[3]  ( .D(n777), .CK(clock), .Q(DI_adr[3]) );
  FLIP_FLOP_D \DI_adr_reg[2]  ( .D(n776), .CK(clock), .Q(DI_adr[2]) );
  FLIP_FLOP_D \DI_adr_reg[1]  ( .D(n775), .CK(clock), .Q(DI_adr[1]) );
  FLIP_FLOP_D \DI_adr_reg[0]  ( .D(n774), .CK(clock), .Q(DI_adr[0]) );
  FLIP_FLOP_D \DI_exc_cause_reg[31]  ( .D(n773), .CK(clock), .Q(
        DI_exc_cause[31]) );
  FLIP_FLOP_D \DI_exc_cause_reg[30]  ( .D(n772), .CK(clock), .Q(
        DI_exc_cause[30]) );
  FLIP_FLOP_D \DI_exc_cause_reg[29]  ( .D(n771), .CK(clock), .Q(
        DI_exc_cause[29]) );
  FLIP_FLOP_D \DI_exc_cause_reg[28]  ( .D(n770), .CK(clock), .Q(
        DI_exc_cause[28]) );
  FLIP_FLOP_D \DI_exc_cause_reg[27]  ( .D(n769), .CK(clock), .Q(
        DI_exc_cause[27]) );
  FLIP_FLOP_D \DI_exc_cause_reg[26]  ( .D(n768), .CK(clock), .Q(
        DI_exc_cause[26]) );
  FLIP_FLOP_D \DI_exc_cause_reg[25]  ( .D(n767), .CK(clock), .Q(
        DI_exc_cause[25]) );
  FLIP_FLOP_D \DI_exc_cause_reg[24]  ( .D(n766), .CK(clock), .Q(
        DI_exc_cause[24]) );
  FLIP_FLOP_D \DI_exc_cause_reg[23]  ( .D(n765), .CK(clock), .Q(
        DI_exc_cause[23]) );
  FLIP_FLOP_D \DI_exc_cause_reg[22]  ( .D(n764), .CK(clock), .Q(
        DI_exc_cause[22]) );
  FLIP_FLOP_D \DI_exc_cause_reg[21]  ( .D(n763), .CK(clock), .Q(
        DI_exc_cause[21]) );
  FLIP_FLOP_D \DI_exc_cause_reg[20]  ( .D(n762), .CK(clock), .Q(
        DI_exc_cause[20]) );
  FLIP_FLOP_D \DI_exc_cause_reg[19]  ( .D(n761), .CK(clock), .Q(
        DI_exc_cause[19]) );
  FLIP_FLOP_D \DI_exc_cause_reg[18]  ( .D(n760), .CK(clock), .Q(
        DI_exc_cause[18]) );
  FLIP_FLOP_D \DI_exc_cause_reg[17]  ( .D(n759), .CK(clock), .Q(
        DI_exc_cause[17]) );
  FLIP_FLOP_D \DI_exc_cause_reg[16]  ( .D(n758), .CK(clock), .Q(
        DI_exc_cause[16]) );
  FLIP_FLOP_D \DI_exc_cause_reg[15]  ( .D(n757), .CK(clock), .Q(
        DI_exc_cause[15]) );
  FLIP_FLOP_D \DI_exc_cause_reg[14]  ( .D(n756), .CK(clock), .Q(
        DI_exc_cause[14]) );
  FLIP_FLOP_D \DI_exc_cause_reg[13]  ( .D(n755), .CK(clock), .Q(
        DI_exc_cause[13]) );
  FLIP_FLOP_D \DI_exc_cause_reg[12]  ( .D(n754), .CK(clock), .Q(
        DI_exc_cause[12]) );
  FLIP_FLOP_D \DI_exc_cause_reg[11]  ( .D(n753), .CK(clock), .Q(
        DI_exc_cause[11]) );
  FLIP_FLOP_D \DI_exc_cause_reg[10]  ( .D(n752), .CK(clock), .Q(
        DI_exc_cause[10]) );
  FLIP_FLOP_D \DI_exc_cause_reg[9]  ( .D(n751), .CK(clock), .Q(DI_exc_cause[9]) );
  FLIP_FLOP_D \DI_exc_cause_reg[8]  ( .D(n750), .CK(clock), .Q(DI_exc_cause[8]) );
  FLIP_FLOP_D \DI_exc_cause_reg[7]  ( .D(n749), .CK(clock), .Q(DI_exc_cause[7]) );
  FLIP_FLOP_D \DI_exc_cause_reg[6]  ( .D(n748), .CK(clock), .Q(DI_exc_cause[6]) );
  FLIP_FLOP_D \DI_exc_cause_reg[5]  ( .D(n747), .CK(clock), .Q(DI_exc_cause[5]) );
  FLIP_FLOP_D \DI_exc_cause_reg[4]  ( .D(n746), .CK(clock), .Q(DI_exc_cause[4]) );
  FLIP_FLOP_D \DI_exc_cause_reg[3]  ( .D(n745), .CK(clock), .Q(DI_exc_cause[3]) );
  FLIP_FLOP_D \DI_exc_cause_reg[2]  ( .D(n744), .CK(clock), .Q(DI_exc_cause[2]) );
  FLIP_FLOP_D \DI_exc_cause_reg[1]  ( .D(n743), .CK(clock), .Q(DI_exc_cause[1]) );
  FLIP_FLOP_D \DI_exc_cause_reg[0]  ( .D(n742), .CK(clock), .Q(DI_exc_cause[0]) );
  FLIP_FLOP_D \DI_level_reg[1]  ( .D(n741), .CK(clock), .Q(DI_level[1]) );
  FLIP_FLOP_D \DI_level_reg[0]  ( .D(n740), .CK(clock), .Q(DI_level[0]) );
  AND_GATE U37 ( .I1(n36), .I2(n23), .O(use1) );
  NAND5_GATE U38 ( .I1(n37), .I2(n38), .I3(n39), .I4(n40), .I5(n41), .O(n36)
         );
  OR_GATE U39 ( .I1(n33), .I2(n948), .O(n41) );
  OR_GATE U40 ( .I1(n42), .I2(n43), .O(n40) );
  NAND_GATE U41 ( .I1(n44), .I2(n27), .O(n39) );
  NAND5_GATE U42 ( .I1(n45), .I2(n32), .I3(n46), .I4(n43), .I5(n47), .O(n44)
         );
  OR_GATE U43 ( .I1(n48), .I2(n49), .O(n47) );
  OR_GATE U44 ( .I1(n34), .I2(n948), .O(n46) );
  OR3_GATE U45 ( .I1(n48), .I2(n944), .I3(n35), .O(n38) );
  NAND_GATE U46 ( .I1(n50), .I2(n51), .O(n37) );
  OR_GATE U47 ( .I1(n52), .I2(n53), .O(n50) );
  NAND_GATE U48 ( .I1(n54), .I2(n55), .O(n740) );
  NAND_GATE U49 ( .I1(n56), .I2(n17), .O(n55) );
  NAND4_GATE U50 ( .I1(n57), .I2(n58), .I3(n59), .I4(n60), .O(n56) );
  AND3_GATE U51 ( .I1(n61), .I2(n62), .I3(n63), .O(n60) );
  NAND_GATE U52 ( .I1(n52), .I2(n64), .O(n62) );
  NAND_GATE U53 ( .I1(n65), .I2(n944), .O(n61) );
  NAND_GATE U54 ( .I1(n66), .I2(n945), .O(n59) );
  OR_GATE U55 ( .I1(n943), .I2(n67), .O(n66) );
  NAND3_GATE U56 ( .I1(n68), .I2(n69), .I3(n70), .O(n58) );
  NAND3_GATE U57 ( .I1(n71), .I2(n34), .I3(n43), .O(n57) );
  NAND_GATE U58 ( .I1(DI_level[0]), .I2(n16), .O(n54) );
  NAND_GATE U59 ( .I1(n73), .I2(n74), .O(n741) );
  NAND_GATE U60 ( .I1(n75), .I2(n17), .O(n74) );
  NAND5_GATE U61 ( .I1(n26), .I2(n49), .I3(n948), .I4(n76), .I5(n77), .O(n75)
         );
  NAND_GATE U62 ( .I1(DI_level[1]), .I2(n16), .O(n73) );
  AND_GATE U63 ( .I1(DI_exc_cause[0]), .I2(n16), .O(n742) );
  AND_GATE U64 ( .I1(DI_exc_cause[1]), .I2(n16), .O(n743) );
  NAND_GATE U65 ( .I1(n78), .I2(n79), .O(n744) );
  NAND3_GATE U66 ( .I1(n80), .I2(n81), .I3(n82), .O(n79) );
  NAND_GATE U67 ( .I1(DI_exc_cause[2]), .I2(n16), .O(n78) );
  NAND_GATE U68 ( .I1(n83), .I2(n84), .O(n745) );
  NAND4_GATE U69 ( .I1(n85), .I2(n76), .I3(n18), .I4(n42), .O(n84) );
  NAND_GATE U70 ( .I1(DI_exc_cause[3]), .I2(n16), .O(n83) );
  NAND_GATE U71 ( .I1(n86), .I2(n87), .O(n746) );
  NAND4_GATE U72 ( .I1(n88), .I2(n76), .I3(n68), .I4(n18), .O(n87) );
  NAND_GATE U73 ( .I1(DI_exc_cause[4]), .I2(n15), .O(n86) );
  AND_GATE U74 ( .I1(DI_exc_cause[5]), .I2(n15), .O(n747) );
  AND_GATE U75 ( .I1(DI_exc_cause[6]), .I2(n15), .O(n748) );
  AND_GATE U76 ( .I1(DI_exc_cause[7]), .I2(n15), .O(n749) );
  AND_GATE U77 ( .I1(DI_exc_cause[8]), .I2(n15), .O(n750) );
  AND_GATE U78 ( .I1(DI_exc_cause[9]), .I2(n15), .O(n751) );
  AND_GATE U79 ( .I1(DI_exc_cause[10]), .I2(n15), .O(n752) );
  AND_GATE U80 ( .I1(DI_exc_cause[11]), .I2(n15), .O(n753) );
  AND_GATE U81 ( .I1(DI_exc_cause[12]), .I2(n15), .O(n754) );
  AND_GATE U82 ( .I1(DI_exc_cause[13]), .I2(n16), .O(n755) );
  AND_GATE U83 ( .I1(DI_exc_cause[14]), .I2(n16), .O(n756) );
  AND_GATE U84 ( .I1(DI_exc_cause[15]), .I2(n16), .O(n757) );
  AND_GATE U85 ( .I1(DI_exc_cause[16]), .I2(n8), .O(n758) );
  AND_GATE U86 ( .I1(DI_exc_cause[17]), .I2(n15), .O(n759) );
  AND_GATE U87 ( .I1(DI_exc_cause[18]), .I2(n16), .O(n760) );
  AND_GATE U88 ( .I1(DI_exc_cause[19]), .I2(n2), .O(n761) );
  AND_GATE U89 ( .I1(DI_exc_cause[20]), .I2(n3), .O(n762) );
  AND_GATE U90 ( .I1(DI_exc_cause[21]), .I2(n12), .O(n763) );
  AND_GATE U91 ( .I1(DI_exc_cause[22]), .I2(n13), .O(n764) );
  AND_GATE U92 ( .I1(DI_exc_cause[23]), .I2(n14), .O(n765) );
  AND_GATE U93 ( .I1(DI_exc_cause[24]), .I2(n8), .O(n766) );
  AND_GATE U94 ( .I1(DI_exc_cause[25]), .I2(n15), .O(n767) );
  AND_GATE U95 ( .I1(DI_exc_cause[26]), .I2(n16), .O(n768) );
  AND_GATE U96 ( .I1(DI_exc_cause[27]), .I2(n2), .O(n769) );
  AND_GATE U97 ( .I1(DI_exc_cause[28]), .I2(n3), .O(n770) );
  AND_GATE U98 ( .I1(DI_exc_cause[29]), .I2(n12), .O(n771) );
  AND_GATE U99 ( .I1(DI_exc_cause[30]), .I2(n13), .O(n772) );
  AND_GATE U100 ( .I1(DI_exc_cause[31]), .I2(n14), .O(n773) );
  NAND_GATE U101 ( .I1(n89), .I2(n90), .O(n774) );
  NAND_GATE U102 ( .I1(EI_adr[0]), .I2(n82), .O(n90) );
  NAND_GATE U103 ( .I1(DI_adr[0]), .I2(n14), .O(n89) );
  NAND_GATE U104 ( .I1(n91), .I2(n92), .O(n775) );
  NAND_GATE U105 ( .I1(EI_adr[1]), .I2(n82), .O(n92) );
  NAND_GATE U106 ( .I1(DI_adr[1]), .I2(n14), .O(n91) );
  NAND_GATE U107 ( .I1(n93), .I2(n94), .O(n776) );
  NAND_GATE U108 ( .I1(EI_adr[2]), .I2(n82), .O(n94) );
  NAND_GATE U109 ( .I1(DI_adr[2]), .I2(n14), .O(n93) );
  NAND_GATE U110 ( .I1(n95), .I2(n96), .O(n777) );
  NAND_GATE U111 ( .I1(EI_adr[3]), .I2(n82), .O(n96) );
  NAND_GATE U112 ( .I1(DI_adr[3]), .I2(n14), .O(n95) );
  NAND_GATE U113 ( .I1(n97), .I2(n98), .O(n778) );
  NAND_GATE U114 ( .I1(EI_adr[4]), .I2(n82), .O(n98) );
  NAND_GATE U115 ( .I1(DI_adr[4]), .I2(n14), .O(n97) );
  NAND_GATE U116 ( .I1(n99), .I2(n100), .O(n779) );
  NAND_GATE U117 ( .I1(EI_adr[5]), .I2(n82), .O(n100) );
  NAND_GATE U118 ( .I1(DI_adr[5]), .I2(n14), .O(n99) );
  NAND_GATE U119 ( .I1(n101), .I2(n102), .O(n780) );
  NAND_GATE U120 ( .I1(EI_adr[6]), .I2(n82), .O(n102) );
  NAND_GATE U121 ( .I1(DI_adr[6]), .I2(n14), .O(n101) );
  NAND_GATE U122 ( .I1(n103), .I2(n104), .O(n781) );
  NAND_GATE U123 ( .I1(EI_adr[7]), .I2(n82), .O(n104) );
  NAND_GATE U124 ( .I1(DI_adr[7]), .I2(n14), .O(n103) );
  NAND_GATE U125 ( .I1(n105), .I2(n106), .O(n782) );
  NAND_GATE U126 ( .I1(EI_adr[8]), .I2(n82), .O(n106) );
  NAND_GATE U127 ( .I1(DI_adr[8]), .I2(n13), .O(n105) );
  NAND_GATE U128 ( .I1(n107), .I2(n108), .O(n783) );
  NAND_GATE U129 ( .I1(EI_adr[9]), .I2(n82), .O(n108) );
  NAND_GATE U130 ( .I1(DI_adr[9]), .I2(n13), .O(n107) );
  NAND_GATE U131 ( .I1(n109), .I2(n110), .O(n784) );
  NAND_GATE U132 ( .I1(EI_adr[10]), .I2(n82), .O(n110) );
  NAND_GATE U133 ( .I1(DI_adr[10]), .I2(n13), .O(n109) );
  NAND_GATE U134 ( .I1(n111), .I2(n112), .O(n785) );
  NAND_GATE U135 ( .I1(EI_adr[11]), .I2(n82), .O(n112) );
  NAND_GATE U136 ( .I1(DI_adr[11]), .I2(n13), .O(n111) );
  NAND_GATE U137 ( .I1(n113), .I2(n114), .O(n786) );
  NAND_GATE U138 ( .I1(EI_adr[12]), .I2(n82), .O(n114) );
  NAND_GATE U139 ( .I1(DI_adr[12]), .I2(n13), .O(n113) );
  NAND_GATE U140 ( .I1(n115), .I2(n116), .O(n787) );
  NAND_GATE U141 ( .I1(EI_adr[13]), .I2(n82), .O(n116) );
  NAND_GATE U142 ( .I1(DI_adr[13]), .I2(n13), .O(n115) );
  NAND_GATE U143 ( .I1(n117), .I2(n118), .O(n788) );
  NAND_GATE U144 ( .I1(EI_adr[14]), .I2(n82), .O(n118) );
  NAND_GATE U145 ( .I1(DI_adr[14]), .I2(n13), .O(n117) );
  NAND_GATE U146 ( .I1(n119), .I2(n120), .O(n789) );
  NAND_GATE U147 ( .I1(EI_adr[15]), .I2(n82), .O(n120) );
  NAND_GATE U148 ( .I1(DI_adr[15]), .I2(n13), .O(n119) );
  NAND_GATE U149 ( .I1(n121), .I2(n122), .O(n790) );
  NAND_GATE U150 ( .I1(EI_adr[16]), .I2(n82), .O(n122) );
  NAND_GATE U151 ( .I1(DI_adr[16]), .I2(n13), .O(n121) );
  NAND_GATE U152 ( .I1(n123), .I2(n124), .O(n791) );
  NAND_GATE U153 ( .I1(EI_adr[17]), .I2(n82), .O(n124) );
  NAND_GATE U154 ( .I1(DI_adr[17]), .I2(n12), .O(n123) );
  NAND_GATE U155 ( .I1(n125), .I2(n126), .O(n792) );
  NAND_GATE U156 ( .I1(EI_adr[18]), .I2(n82), .O(n126) );
  NAND_GATE U157 ( .I1(DI_adr[18]), .I2(n12), .O(n125) );
  NAND_GATE U158 ( .I1(n127), .I2(n128), .O(n793) );
  NAND_GATE U159 ( .I1(EI_adr[19]), .I2(n82), .O(n128) );
  NAND_GATE U160 ( .I1(DI_adr[19]), .I2(n12), .O(n127) );
  NAND_GATE U161 ( .I1(n129), .I2(n130), .O(n794) );
  NAND_GATE U162 ( .I1(EI_adr[20]), .I2(n82), .O(n130) );
  NAND_GATE U163 ( .I1(DI_adr[20]), .I2(n12), .O(n129) );
  NAND_GATE U164 ( .I1(n131), .I2(n132), .O(n795) );
  NAND_GATE U165 ( .I1(EI_adr[21]), .I2(n82), .O(n132) );
  NAND_GATE U166 ( .I1(DI_adr[21]), .I2(n12), .O(n131) );
  NAND_GATE U167 ( .I1(n133), .I2(n134), .O(n796) );
  NAND_GATE U168 ( .I1(EI_adr[22]), .I2(n82), .O(n134) );
  NAND_GATE U169 ( .I1(DI_adr[22]), .I2(n12), .O(n133) );
  NAND_GATE U170 ( .I1(n135), .I2(n136), .O(n797) );
  NAND_GATE U171 ( .I1(EI_adr[23]), .I2(n82), .O(n136) );
  NAND_GATE U172 ( .I1(DI_adr[23]), .I2(n12), .O(n135) );
  NAND_GATE U173 ( .I1(n137), .I2(n138), .O(n798) );
  NAND_GATE U174 ( .I1(EI_adr[24]), .I2(n82), .O(n138) );
  NAND_GATE U175 ( .I1(DI_adr[24]), .I2(n12), .O(n137) );
  NAND_GATE U176 ( .I1(n139), .I2(n140), .O(n799) );
  NAND_GATE U177 ( .I1(EI_adr[25]), .I2(n82), .O(n140) );
  NAND_GATE U178 ( .I1(DI_adr[25]), .I2(n12), .O(n139) );
  NAND_GATE U179 ( .I1(n141), .I2(n142), .O(n800) );
  NAND_GATE U180 ( .I1(EI_adr[26]), .I2(n82), .O(n142) );
  NAND_GATE U181 ( .I1(DI_adr[26]), .I2(n14), .O(n141) );
  NAND_GATE U182 ( .I1(n143), .I2(n144), .O(n801) );
  NAND_GATE U183 ( .I1(EI_adr[27]), .I2(n82), .O(n144) );
  NAND_GATE U184 ( .I1(DI_adr[27]), .I2(n8), .O(n143) );
  NAND_GATE U185 ( .I1(n145), .I2(n146), .O(n802) );
  NAND_GATE U186 ( .I1(EI_adr[28]), .I2(n82), .O(n146) );
  NAND_GATE U187 ( .I1(DI_adr[28]), .I2(n15), .O(n145) );
  NAND_GATE U188 ( .I1(n147), .I2(n148), .O(n803) );
  NAND_GATE U189 ( .I1(EI_adr[29]), .I2(n82), .O(n148) );
  NAND_GATE U190 ( .I1(DI_adr[29]), .I2(n16), .O(n147) );
  NAND_GATE U191 ( .I1(n149), .I2(n150), .O(n804) );
  NAND_GATE U192 ( .I1(EI_adr[30]), .I2(n82), .O(n150) );
  NAND_GATE U193 ( .I1(DI_adr[30]), .I2(n12), .O(n149) );
  NAND_GATE U194 ( .I1(n151), .I2(n152), .O(n805) );
  NAND_GATE U195 ( .I1(EI_adr[31]), .I2(n82), .O(n152) );
  NAND_GATE U196 ( .I1(DI_adr[31]), .I2(n13), .O(n151) );
  NAND_GATE U197 ( .I1(n153), .I2(n154), .O(n806) );
  NAND_GATE U198 ( .I1(DI_r_w), .I2(n2), .O(n154) );
  NAND3_GATE U199 ( .I1(n155), .I2(n153), .I3(n156), .O(n807) );
  NAND_GATE U200 ( .I1(DI_op_mem), .I2(n9), .O(n156) );
  NAND_GATE U201 ( .I1(n157), .I2(n77), .O(n155) );
  NAND_GATE U202 ( .I1(n158), .I2(n159), .O(n808) );
  OR_GATE U203 ( .I1(n20), .I2(n160), .O(n159) );
  NAND_GATE U204 ( .I1(DI_mode), .I2(n3), .O(n158) );
  NAND_GATE U205 ( .I1(n162), .I2(n163), .O(n809) );
  NAND_GATE U206 ( .I1(n161), .I2(n164), .O(n163) );
  NAND5_GATE U207 ( .I1(n165), .I2(n30), .I3(n166), .I4(n28), .I5(n167), .O(
        n164) );
  AND3_GATE U208 ( .I1(n168), .I2(n169), .I3(n170), .O(n167) );
  NAND_GATE U209 ( .I1(n171), .I2(n77), .O(n170) );
  NAND_GATE U210 ( .I1(n48), .I2(n172), .O(n169) );
  OR3_GATE U211 ( .I1(n68), .I2(n171), .I3(n173), .O(n172) );
  OR_GATE U212 ( .I1(n29), .I2(n32), .O(n168) );
  NAND_GATE U213 ( .I1(n175), .I2(n176), .O(n165) );
  NAND_GATE U214 ( .I1(n70), .I2(n34), .O(n176) );
  NAND_GATE U215 ( .I1(DI_ecr_reg), .I2(n14), .O(n162) );
  NAND4_GATE U216 ( .I1(n177), .I2(n178), .I3(n179), .I4(n180), .O(n810) );
  NAND_GATE U217 ( .I1(EI_instr[11]), .I2(n181), .O(n179) );
  NAND_GATE U218 ( .I1(adr_reg2[0]), .I2(n182), .O(n178) );
  NAND_GATE U219 ( .I1(DI_adr_reg_dest[0]), .I2(n1), .O(n177) );
  NAND4_GATE U220 ( .I1(n183), .I2(n184), .I3(n185), .I4(n180), .O(n811) );
  NAND_GATE U221 ( .I1(EI_instr[12]), .I2(n181), .O(n185) );
  NAND_GATE U222 ( .I1(adr_reg2[1]), .I2(n182), .O(n184) );
  NAND_GATE U223 ( .I1(DI_adr_reg_dest[1]), .I2(n10), .O(n183) );
  NAND4_GATE U224 ( .I1(n186), .I2(n187), .I3(n188), .I4(n180), .O(n812) );
  NAND_GATE U225 ( .I1(EI_instr[13]), .I2(n181), .O(n188) );
  NAND_GATE U226 ( .I1(adr_reg2[2]), .I2(n182), .O(n187) );
  NAND_GATE U227 ( .I1(DI_adr_reg_dest[2]), .I2(n11), .O(n186) );
  NAND4_GATE U228 ( .I1(n189), .I2(n190), .I3(n191), .I4(n180), .O(n813) );
  NAND_GATE U229 ( .I1(EI_instr[14]), .I2(n181), .O(n191) );
  NAND_GATE U230 ( .I1(adr_reg2[3]), .I2(n182), .O(n190) );
  NAND_GATE U231 ( .I1(DI_adr_reg_dest[3]), .I2(n10), .O(n189) );
  NAND4_GATE U232 ( .I1(n192), .I2(n193), .I3(n194), .I4(n180), .O(n814) );
  OR3_GATE U233 ( .I1(n195), .I2(n196), .I3(n25), .O(n180) );
  NAND_GATE U234 ( .I1(EI_instr[15]), .I2(n181), .O(n194) );
  AND3_GATE U235 ( .I1(n21), .I2(n25), .I3(n196), .O(n181) );
  AND3_GATE U236 ( .I1(n197), .I2(n198), .I3(n199), .O(n196) );
  OR_GATE U237 ( .I1(n200), .I2(n31), .O(n199) );
  OR_GATE U238 ( .I1(n201), .I2(n32), .O(n198) );
  NAND_GATE U239 ( .I1(n85), .I2(n945), .O(n197) );
  NAND_GATE U240 ( .I1(adr_reg2[4]), .I2(n182), .O(n193) );
  AND_GATE U241 ( .I1(n202), .I2(n203), .O(n182) );
  AND4_GATE U242 ( .I1(n204), .I2(n205), .I3(n206), .I4(n207), .O(n202) );
  AND4_GATE U243 ( .I1(n208), .I2(n209), .I3(n210), .I4(n166), .O(n207) );
  NAND3_GATE U244 ( .I1(n70), .I2(n43), .I3(n52), .O(n166) );
  NAND_GATE U245 ( .I1(n88), .I2(n211), .O(n209) );
  NAND3_GATE U246 ( .I1(n212), .I2(n944), .I3(n213), .O(n208) );
  OR_GATE U247 ( .I1(n175), .I2(n64), .O(n212) );
  NAND_GATE U248 ( .I1(n52), .I2(n214), .O(n206) );
  NAND3_GATE U249 ( .I1(n215), .I2(n216), .I3(n217), .O(n214) );
  NAND_GATE U250 ( .I1(n69), .I2(n27), .O(n217) );
  OR_GATE U251 ( .I1(n947), .I2(n944), .O(n216) );
  OR_GATE U252 ( .I1(n948), .I2(n26), .O(n215) );
  OR_GATE U253 ( .I1(n45), .I2(n31), .O(n205) );
  NAND_GATE U254 ( .I1(n218), .I2(n34), .O(n204) );
  NAND_GATE U255 ( .I1(DI_adr_reg_dest[4]), .I2(n1), .O(n192) );
  NAND_GATE U256 ( .I1(n219), .I2(n220), .O(n815) );
  NAND4_GATE U257 ( .I1(n161), .I2(n43), .I3(n221), .I4(n34), .O(n220) );
  NAND_GATE U258 ( .I1(n222), .I2(n223), .O(n221) );
  NAND3_GATE U259 ( .I1(n48), .I2(n945), .I3(n70), .O(n223) );
  NAND3_GATE U260 ( .I1(n948), .I2(n42), .I3(n71), .O(n222) );
  OR_GATE U261 ( .I1(n224), .I2(n225), .O(n71) );
  NOR_GATE U262 ( .I1(n49), .I2(n27), .O(n225) );
  NAND_GATE U263 ( .I1(DI_adr_reg_dest[5]), .I2(n8), .O(n219) );
  NAND_GATE U264 ( .I1(n226), .I2(n227), .O(n816) );
  NAND3_GATE U265 ( .I1(n161), .I2(EI_instr[0]), .I3(n228), .O(n227) );
  NAND_GATE U266 ( .I1(DI_offset[0]), .I2(n2), .O(n226) );
  NAND_GATE U267 ( .I1(n229), .I2(n230), .O(n817) );
  NAND3_GATE U268 ( .I1(n161), .I2(EI_instr[1]), .I3(n228), .O(n230) );
  NAND_GATE U269 ( .I1(DI_offset[1]), .I2(n15), .O(n229) );
  NAND3_GATE U270 ( .I1(n231), .I2(n232), .I3(n233), .O(n818) );
  NAND_GATE U271 ( .I1(DI_offset[2]), .I2(n4), .O(n233) );
  NAND_GATE U272 ( .I1(n234), .I2(EI_instr[0]), .O(n232) );
  NAND_GATE U273 ( .I1(n235), .I2(EI_instr[2]), .O(n231) );
  NAND3_GATE U274 ( .I1(n236), .I2(n237), .I3(n238), .O(n819) );
  NAND_GATE U275 ( .I1(DI_offset[3]), .I2(n5), .O(n238) );
  NAND_GATE U276 ( .I1(n234), .I2(EI_instr[1]), .O(n237) );
  NAND_GATE U277 ( .I1(n235), .I2(EI_instr[3]), .O(n236) );
  NAND3_GATE U278 ( .I1(n239), .I2(n240), .I3(n241), .O(n820) );
  NAND_GATE U279 ( .I1(DI_offset[4]), .I2(n6), .O(n241) );
  NAND_GATE U280 ( .I1(n234), .I2(EI_instr[2]), .O(n240) );
  NAND_GATE U281 ( .I1(n235), .I2(EI_instr[4]), .O(n239) );
  NAND3_GATE U282 ( .I1(n242), .I2(n243), .I3(n244), .O(n821) );
  NAND_GATE U283 ( .I1(DI_offset[5]), .I2(n7), .O(n244) );
  NAND_GATE U284 ( .I1(n234), .I2(EI_instr[3]), .O(n243) );
  NAND_GATE U285 ( .I1(n235), .I2(EI_instr[5]), .O(n242) );
  NAND3_GATE U286 ( .I1(n245), .I2(n246), .I3(n247), .O(n822) );
  NAND_GATE U287 ( .I1(DI_offset[6]), .I2(n9), .O(n247) );
  NAND_GATE U288 ( .I1(n234), .I2(EI_instr[4]), .O(n246) );
  NAND_GATE U289 ( .I1(EI_instr[6]), .I2(n235), .O(n245) );
  NAND3_GATE U290 ( .I1(n248), .I2(n249), .I3(n250), .O(n823) );
  NAND_GATE U291 ( .I1(DI_offset[7]), .I2(n4), .O(n250) );
  NAND_GATE U292 ( .I1(n234), .I2(EI_instr[5]), .O(n249) );
  NAND_GATE U293 ( .I1(EI_instr[7]), .I2(n235), .O(n248) );
  NAND3_GATE U294 ( .I1(n251), .I2(n252), .I3(n253), .O(n824) );
  NAND_GATE U295 ( .I1(DI_offset[8]), .I2(n5), .O(n253) );
  NAND_GATE U296 ( .I1(EI_instr[6]), .I2(n234), .O(n252) );
  NAND_GATE U297 ( .I1(EI_instr[8]), .I2(n235), .O(n251) );
  NAND3_GATE U298 ( .I1(n254), .I2(n255), .I3(n256), .O(n825) );
  NAND_GATE U299 ( .I1(DI_offset[9]), .I2(n6), .O(n256) );
  NAND_GATE U300 ( .I1(EI_instr[7]), .I2(n234), .O(n255) );
  NAND_GATE U301 ( .I1(EI_instr[9]), .I2(n235), .O(n254) );
  NAND3_GATE U302 ( .I1(n257), .I2(n258), .I3(n259), .O(n826) );
  NAND_GATE U303 ( .I1(DI_offset[10]), .I2(n7), .O(n259) );
  NAND_GATE U304 ( .I1(EI_instr[8]), .I2(n234), .O(n258) );
  NAND_GATE U305 ( .I1(EI_instr[10]), .I2(n235), .O(n257) );
  NAND3_GATE U306 ( .I1(n260), .I2(n261), .I3(n262), .O(n827) );
  NAND_GATE U307 ( .I1(DI_offset[11]), .I2(n9), .O(n262) );
  NAND_GATE U308 ( .I1(EI_instr[9]), .I2(n234), .O(n261) );
  NAND_GATE U309 ( .I1(n235), .I2(EI_instr[11]), .O(n260) );
  NAND3_GATE U310 ( .I1(n263), .I2(n264), .I3(n265), .O(n828) );
  NAND_GATE U311 ( .I1(DI_offset[12]), .I2(n4), .O(n265) );
  NAND_GATE U312 ( .I1(EI_instr[10]), .I2(n234), .O(n264) );
  NAND_GATE U313 ( .I1(n235), .I2(EI_instr[12]), .O(n263) );
  NAND3_GATE U314 ( .I1(n266), .I2(n267), .I3(n268), .O(n829) );
  NAND_GATE U315 ( .I1(DI_offset[13]), .I2(n5), .O(n268) );
  NAND_GATE U316 ( .I1(n234), .I2(EI_instr[11]), .O(n267) );
  NAND_GATE U317 ( .I1(n235), .I2(EI_instr[13]), .O(n266) );
  NAND3_GATE U318 ( .I1(n269), .I2(n270), .I3(n271), .O(n830) );
  NAND_GATE U319 ( .I1(DI_offset[14]), .I2(n6), .O(n271) );
  NAND_GATE U320 ( .I1(n234), .I2(EI_instr[12]), .O(n270) );
  NAND_GATE U321 ( .I1(n235), .I2(EI_instr[14]), .O(n269) );
  NAND3_GATE U322 ( .I1(n272), .I2(n273), .I3(n274), .O(n831) );
  NAND_GATE U323 ( .I1(DI_offset[15]), .I2(n7), .O(n274) );
  NAND_GATE U324 ( .I1(n234), .I2(EI_instr[13]), .O(n272) );
  NAND3_GATE U325 ( .I1(n275), .I2(n273), .I3(n276), .O(n832) );
  NAND_GATE U326 ( .I1(DI_offset[16]), .I2(n14), .O(n276) );
  NAND_GATE U327 ( .I1(n234), .I2(EI_instr[14]), .O(n275) );
  NAND3_GATE U328 ( .I1(n277), .I2(n273), .I3(n278), .O(n833) );
  NAND_GATE U329 ( .I1(DI_offset[17]), .I2(n9), .O(n278) );
  NAND_GATE U330 ( .I1(n234), .I2(EI_instr[15]), .O(n277) );
  AND_GATE U331 ( .I1(n21), .I2(n279), .O(n234) );
  OR_GATE U332 ( .I1(n280), .I2(n281), .O(n279) );
  NAND3_GATE U333 ( .I1(n282), .I2(n283), .I3(n284), .O(n834) );
  NAND_GATE U334 ( .I1(n285), .I2(adr_reg2[0]), .O(n283) );
  NAND_GATE U335 ( .I1(DI_offset[18]), .I2(n4), .O(n282) );
  NAND3_GATE U336 ( .I1(n286), .I2(n287), .I3(n284), .O(n835) );
  NAND_GATE U337 ( .I1(n285), .I2(adr_reg2[1]), .O(n287) );
  NAND_GATE U338 ( .I1(DI_offset[19]), .I2(n5), .O(n286) );
  NAND3_GATE U339 ( .I1(n288), .I2(n289), .I3(n284), .O(n836) );
  NAND_GATE U340 ( .I1(n285), .I2(adr_reg2[2]), .O(n289) );
  NAND_GATE U341 ( .I1(DI_offset[20]), .I2(n11), .O(n288) );
  NAND3_GATE U342 ( .I1(n290), .I2(n291), .I3(n284), .O(n837) );
  NAND_GATE U343 ( .I1(n285), .I2(adr_reg2[3]), .O(n291) );
  NAND_GATE U344 ( .I1(DI_offset[21]), .I2(n11), .O(n290) );
  NAND3_GATE U345 ( .I1(n292), .I2(n293), .I3(n284), .O(n838) );
  NAND_GATE U346 ( .I1(n285), .I2(adr_reg2[4]), .O(n293) );
  NAND_GATE U347 ( .I1(DI_offset[22]), .I2(n11), .O(n292) );
  NAND3_GATE U348 ( .I1(n294), .I2(n295), .I3(n284), .O(n839) );
  NAND_GATE U349 ( .I1(adr_reg1[0]), .I2(n285), .O(n295) );
  NAND_GATE U350 ( .I1(DI_offset[23]), .I2(n11), .O(n294) );
  NAND3_GATE U351 ( .I1(n296), .I2(n297), .I3(n284), .O(n840) );
  NAND_GATE U352 ( .I1(adr_reg1[1]), .I2(n285), .O(n297) );
  NAND_GATE U353 ( .I1(DI_offset[24]), .I2(n11), .O(n296) );
  NAND3_GATE U354 ( .I1(n298), .I2(n299), .I3(n284), .O(n841) );
  NAND_GATE U355 ( .I1(adr_reg1[2]), .I2(n285), .O(n299) );
  NAND_GATE U356 ( .I1(DI_offset[25]), .I2(n11), .O(n298) );
  NAND3_GATE U357 ( .I1(n300), .I2(n301), .I3(n284), .O(n842) );
  NAND_GATE U358 ( .I1(adr_reg1[3]), .I2(n285), .O(n301) );
  NAND_GATE U359 ( .I1(DI_offset[26]), .I2(n11), .O(n300) );
  NAND3_GATE U360 ( .I1(n302), .I2(n303), .I3(n284), .O(n843) );
  NAND_GATE U361 ( .I1(adr_reg1[4]), .I2(n285), .O(n303) );
  AND_GATE U362 ( .I1(n280), .I2(n203), .O(n285) );
  NAND_GATE U363 ( .I1(DI_offset[27]), .I2(n11), .O(n302) );
  NAND3_GATE U364 ( .I1(n304), .I2(n305), .I3(n284), .O(n844) );
  NAND_GATE U365 ( .I1(n306), .I2(EI_adr[28]), .O(n305) );
  NAND_GATE U366 ( .I1(DI_offset[28]), .I2(n11), .O(n304) );
  NAND3_GATE U367 ( .I1(n307), .I2(n308), .I3(n284), .O(n845) );
  NAND_GATE U368 ( .I1(n306), .I2(EI_adr[29]), .O(n308) );
  NAND_GATE U369 ( .I1(DI_offset[29]), .I2(n10), .O(n307) );
  NAND3_GATE U370 ( .I1(n309), .I2(n310), .I3(n284), .O(n846) );
  NAND_GATE U371 ( .I1(n306), .I2(EI_adr[30]), .O(n310) );
  NAND_GATE U372 ( .I1(DI_offset[30]), .I2(n10), .O(n309) );
  NAND3_GATE U373 ( .I1(n311), .I2(n312), .I3(n284), .O(n847) );
  AND_GATE U374 ( .I1(n273), .I2(n313), .O(n284) );
  NAND3_GATE U375 ( .I1(EI_instr[15]), .I2(n21), .I3(n281), .O(n313) );
  NOR_GATE U376 ( .I1(n24), .I2(n314), .O(n281) );
  NAND_GATE U377 ( .I1(n235), .I2(EI_instr[15]), .O(n273) );
  AND_GATE U378 ( .I1(n228), .I2(n21), .O(n235) );
  NOR_GATE U379 ( .I1(n315), .I2(n314), .O(n228) );
  NAND_GATE U380 ( .I1(n306), .I2(EI_adr[31]), .O(n312) );
  AND_GATE U381 ( .I1(n280), .I2(n21), .O(n306) );
  AND_GATE U382 ( .I1(n314), .I2(n315), .O(n280) );
  AND_GATE U383 ( .I1(n316), .I2(n317), .O(n315) );
  NAND3_GATE U384 ( .I1(n318), .I2(n34), .I3(n69), .O(n317) );
  NAND_GATE U385 ( .I1(n26), .I2(n319), .O(n318) );
  OR_GATE U386 ( .I1(n945), .I2(n944), .O(n319) );
  AND3_GATE U387 ( .I1(n316), .I2(n320), .I3(n160), .O(n314) );
  NAND3_GATE U388 ( .I1(n321), .I2(n43), .I3(n224), .O(n320) );
  AND_GATE U389 ( .I1(n322), .I2(n323), .O(n316) );
  NAND_GATE U390 ( .I1(n324), .I2(n944), .O(n323) );
  OR_GATE U391 ( .I1(n28), .I2(n32), .O(n322) );
  NAND_GATE U392 ( .I1(DI_offset[31]), .I2(n10), .O(n311) );
  NAND4_GATE U393 ( .I1(n325), .I2(n326), .I3(n327), .I4(n153), .O(n848) );
  NAND_GATE U394 ( .I1(n328), .I2(n324), .O(n153) );
  NAND_GATE U395 ( .I1(n328), .I2(n329), .O(n327) );
  NAND_GATE U396 ( .I1(n210), .I2(n330), .O(n329) );
  OR_GATE U397 ( .I1(n29), .I2(n35), .O(n210) );
  NAND_GATE U398 ( .I1(n157), .I2(n52), .O(n326) );
  NAND_GATE U399 ( .I1(DI_code_ual[0]), .I2(n10), .O(n325) );
  NAND_GATE U400 ( .I1(n331), .I2(n332), .O(n849) );
  NAND_GATE U401 ( .I1(DI_code_ual[1]), .I2(n10), .O(n332) );
  NAND_GATE U402 ( .I1(n333), .I2(n18), .O(n331) );
  NAND4_GATE U403 ( .I1(n63), .I2(n334), .I3(n335), .I4(n201), .O(n333) );
  NAND3_GATE U404 ( .I1(n77), .I2(n49), .I3(n69), .O(n335) );
  NAND_GATE U405 ( .I1(n85), .I2(n42), .O(n334) );
  AND_GATE U406 ( .I1(n76), .I2(n336), .O(n63) );
  OR3_GATE U407 ( .I1(n26), .I2(n48), .I3(n31), .O(n336) );
  AND3_GATE U408 ( .I1(n23), .I2(n19), .I3(n81), .O(n76) );
  NAND_GATE U409 ( .I1(n337), .I2(n338), .O(n850) );
  NAND_GATE U410 ( .I1(n339), .I2(n68), .O(n338) );
  NAND_GATE U411 ( .I1(DI_code_ual[2]), .I2(n10), .O(n337) );
  NAND_GATE U412 ( .I1(n340), .I2(n341), .O(n851) );
  NAND_GATE U413 ( .I1(n342), .I2(n52), .O(n341) );
  NAND_GATE U414 ( .I1(DI_code_ual[3]), .I2(n10), .O(n340) );
  NAND_GATE U415 ( .I1(n343), .I2(n344), .O(n852) );
  NAND_GATE U416 ( .I1(n342), .I2(n211), .O(n344) );
  NAND_GATE U417 ( .I1(DI_code_ual[4]), .I2(n10), .O(n343) );
  NAND_GATE U418 ( .I1(n345), .I2(n346), .O(n853) );
  NAND_GATE U419 ( .I1(n342), .I2(n68), .O(n346) );
  AND_GATE U420 ( .I1(n328), .I2(n64), .O(n342) );
  NAND_GATE U421 ( .I1(DI_code_ual[5]), .I2(n10), .O(n345) );
  NAND_GATE U422 ( .I1(n347), .I2(n348), .O(n854) );
  NAND_GATE U423 ( .I1(n157), .I2(n68), .O(n348) );
  AND_GATE U424 ( .I1(n67), .I2(n21), .O(n157) );
  NAND_GATE U425 ( .I1(DI_code_ual[6]), .I2(n9), .O(n347) );
  NAND_GATE U426 ( .I1(n349), .I2(n350), .O(n855) );
  NAND3_GATE U427 ( .I1(n328), .I2(n213), .I3(n218), .O(n350) );
  NAND_GATE U428 ( .I1(DI_code_ual[7]), .I2(n9), .O(n349) );
  NAND_GATE U429 ( .I1(n351), .I2(n352), .O(n856) );
  NAND3_GATE U430 ( .I1(n328), .I2(n34), .I3(n218), .O(n352) );
  NAND_GATE U431 ( .I1(DI_code_ual[8]), .I2(n9), .O(n351) );
  NAND_GATE U432 ( .I1(n353), .I2(n354), .O(n857) );
  NAND3_GATE U433 ( .I1(n175), .I2(n34), .I3(n355), .O(n354) );
  NAND_GATE U434 ( .I1(DI_code_ual[9]), .I2(n9), .O(n353) );
  NAND_GATE U435 ( .I1(n356), .I2(n357), .O(n858) );
  NAND_GATE U436 ( .I1(n339), .I2(n321), .O(n357) );
  NAND_GATE U437 ( .I1(DI_code_ual[10]), .I2(n9), .O(n356) );
  NAND_GATE U438 ( .I1(n358), .I2(n359), .O(n859) );
  NAND_GATE U439 ( .I1(n339), .I2(n211), .O(n359) );
  NAND_GATE U440 ( .I1(DI_code_ual[11]), .I2(n9), .O(n358) );
  NAND3_GATE U441 ( .I1(n360), .I2(n361), .I3(n362), .O(n860) );
  NAND_GATE U442 ( .I1(DI_code_ual[12]), .I2(n9), .O(n362) );
  NAND3_GATE U443 ( .I1(n21), .I2(n945), .I3(n363), .O(n361) );
  NAND_GATE U444 ( .I1(n364), .I2(n68), .O(n360) );
  NAND_GATE U445 ( .I1(n365), .I2(n366), .O(n861) );
  NAND_GATE U446 ( .I1(n364), .I2(n321), .O(n366) );
  NAND_GATE U447 ( .I1(DI_code_ual[13]), .I2(n9), .O(n365) );
  NAND_GATE U448 ( .I1(n367), .I2(n368), .O(n862) );
  NAND_GATE U449 ( .I1(n364), .I2(n211), .O(n368) );
  AND_GATE U450 ( .I1(n369), .I2(n51), .O(n364) );
  NAND_GATE U451 ( .I1(DI_code_ual[14]), .I2(n9), .O(n367) );
  NAND_GATE U452 ( .I1(n370), .I2(n371), .O(n863) );
  NAND_GATE U453 ( .I1(n369), .I2(n372), .O(n371) );
  NAND_GATE U454 ( .I1(n373), .I2(n374), .O(n372) );
  NAND_GATE U455 ( .I1(n52), .I2(n51), .O(n374) );
  OR_GATE U456 ( .I1(n31), .I2(n51), .O(n373) );
  NAND_GATE U457 ( .I1(DI_code_ual[15]), .I2(n8), .O(n370) );
  NAND_GATE U458 ( .I1(n375), .I2(n376), .O(n864) );
  NAND3_GATE U459 ( .I1(n211), .I2(n27), .I3(n369), .O(n376) );
  NAND_GATE U460 ( .I1(DI_code_ual[16]), .I2(n8), .O(n375) );
  NAND_GATE U461 ( .I1(n377), .I2(n378), .O(n865) );
  NAND3_GATE U462 ( .I1(n21), .I2(n42), .I3(n363), .O(n378) );
  NAND_GATE U463 ( .I1(DI_code_ual[17]), .I2(n8), .O(n377) );
  NAND_GATE U464 ( .I1(n379), .I2(n380), .O(n866) );
  NAND3_GATE U465 ( .I1(n324), .I2(n49), .I3(n21), .O(n380) );
  NAND_GATE U466 ( .I1(DI_code_ual[18]), .I2(n8), .O(n379) );
  NAND_GATE U467 ( .I1(n381), .I2(n382), .O(n867) );
  NAND_GATE U468 ( .I1(n383), .I2(n175), .O(n382) );
  NAND_GATE U469 ( .I1(DI_code_ual[19]), .I2(n8), .O(n381) );
  NAND_GATE U470 ( .I1(n384), .I2(n385), .O(n868) );
  NAND_GATE U471 ( .I1(n339), .I2(n52), .O(n385) );
  AND3_GATE U472 ( .I1(n69), .I2(n27), .I3(n328), .O(n339) );
  NAND_GATE U473 ( .I1(DI_code_ual[20]), .I2(n8), .O(n384) );
  NAND_GATE U474 ( .I1(n386), .I2(n387), .O(n869) );
  NAND3_GATE U475 ( .I1(n88), .I2(n77), .I3(n355), .O(n387) );
  AND_GATE U476 ( .I1(n948), .I2(n946), .O(n88) );
  NAND_GATE U477 ( .I1(DI_code_ual[21]), .I2(n8), .O(n386) );
  NAND_GATE U478 ( .I1(n388), .I2(n389), .O(n870) );
  NAND3_GATE U479 ( .I1(n175), .I2(n213), .I3(n355), .O(n389) );
  NAND_GATE U480 ( .I1(DI_code_ual[22]), .I2(n8), .O(n388) );
  NAND_GATE U481 ( .I1(n390), .I2(n391), .O(n871) );
  NAND_GATE U482 ( .I1(n383), .I2(n53), .O(n391) );
  AND3_GATE U483 ( .I1(n173), .I2(n27), .I3(n21), .O(n383) );
  NAND_GATE U484 ( .I1(DI_code_ual[23]), .I2(n8), .O(n390) );
  NAND_GATE U485 ( .I1(n392), .I2(n393), .O(n872) );
  NAND_GATE U486 ( .I1(n394), .I2(n211), .O(n393) );
  NAND_GATE U487 ( .I1(DI_code_ual[24]), .I2(n16), .O(n392) );
  NAND_GATE U488 ( .I1(n395), .I2(n396), .O(n873) );
  NAND_GATE U489 ( .I1(n394), .I2(n68), .O(n396) );
  AND3_GATE U490 ( .I1(n328), .I2(n27), .I3(n175), .O(n394) );
  AND_GATE U491 ( .I1(n21), .I2(n944), .O(n328) );
  NAND_GATE U492 ( .I1(DI_code_ual[25]), .I2(n12), .O(n395) );
  NAND_GATE U493 ( .I1(n397), .I2(n398), .O(n874) );
  NAND3_GATE U494 ( .I1(n53), .I2(n34), .I3(n355), .O(n398) );
  NAND_GATE U495 ( .I1(DI_code_ual[26]), .I2(n13), .O(n397) );
  NAND_GATE U496 ( .I1(n399), .I2(n400), .O(n875) );
  NAND3_GATE U497 ( .I1(n53), .I2(n213), .I3(n355), .O(n400) );
  NAND_GATE U498 ( .I1(DI_code_ual[27]), .I2(n3), .O(n399) );
  NAND3_GATE U499 ( .I1(n401), .I2(n402), .I3(n403), .O(n876) );
  NAND_GATE U500 ( .I1(DI_op2[0]), .I2(n4), .O(n403) );
  NAND_GATE U501 ( .I1(n404), .I2(EI_instr[0]), .O(n402) );
  NAND_GATE U502 ( .I1(data2[0]), .I2(n405), .O(n401) );
  NAND3_GATE U503 ( .I1(n406), .I2(n407), .I3(n408), .O(n877) );
  NAND_GATE U504 ( .I1(DI_op2[1]), .I2(n5), .O(n408) );
  NAND_GATE U505 ( .I1(n404), .I2(EI_instr[1]), .O(n407) );
  NAND_GATE U506 ( .I1(data2[1]), .I2(n405), .O(n406) );
  NAND3_GATE U507 ( .I1(n409), .I2(n410), .I3(n411), .O(n878) );
  NAND_GATE U508 ( .I1(DI_op2[2]), .I2(n6), .O(n411) );
  NAND_GATE U509 ( .I1(n404), .I2(EI_instr[2]), .O(n410) );
  NAND_GATE U510 ( .I1(data2[2]), .I2(n405), .O(n409) );
  NAND3_GATE U511 ( .I1(n412), .I2(n413), .I3(n414), .O(n879) );
  NAND_GATE U512 ( .I1(DI_op2[3]), .I2(n7), .O(n414) );
  NAND_GATE U513 ( .I1(n404), .I2(EI_instr[3]), .O(n413) );
  NAND_GATE U514 ( .I1(data2[3]), .I2(n405), .O(n412) );
  NAND3_GATE U515 ( .I1(n415), .I2(n416), .I3(n417), .O(n880) );
  NAND_GATE U516 ( .I1(DI_op2[4]), .I2(n9), .O(n417) );
  NAND_GATE U517 ( .I1(n404), .I2(EI_instr[4]), .O(n416) );
  NAND_GATE U518 ( .I1(data2[4]), .I2(n405), .O(n415) );
  NAND3_GATE U519 ( .I1(n418), .I2(n419), .I3(n420), .O(n881) );
  NAND_GATE U520 ( .I1(DI_op2[5]), .I2(n7), .O(n420) );
  NAND_GATE U521 ( .I1(n404), .I2(EI_instr[5]), .O(n419) );
  NAND_GATE U522 ( .I1(data2[5]), .I2(n405), .O(n418) );
  NAND3_GATE U523 ( .I1(n421), .I2(n422), .I3(n423), .O(n882) );
  NAND_GATE U524 ( .I1(DI_op2[6]), .I2(n7), .O(n423) );
  NAND_GATE U525 ( .I1(n404), .I2(EI_instr[6]), .O(n422) );
  NAND_GATE U526 ( .I1(data2[6]), .I2(n405), .O(n421) );
  NAND3_GATE U527 ( .I1(n424), .I2(n425), .I3(n426), .O(n883) );
  NAND_GATE U528 ( .I1(DI_op2[7]), .I2(n7), .O(n426) );
  NAND_GATE U529 ( .I1(n404), .I2(EI_instr[7]), .O(n425) );
  NAND_GATE U530 ( .I1(data2[7]), .I2(n405), .O(n424) );
  NAND3_GATE U531 ( .I1(n427), .I2(n428), .I3(n429), .O(n884) );
  NAND_GATE U532 ( .I1(DI_op2[8]), .I2(n7), .O(n429) );
  NAND_GATE U533 ( .I1(n404), .I2(EI_instr[8]), .O(n428) );
  NAND_GATE U534 ( .I1(data2[8]), .I2(n405), .O(n427) );
  NAND3_GATE U535 ( .I1(n430), .I2(n431), .I3(n432), .O(n885) );
  NAND_GATE U536 ( .I1(DI_op2[9]), .I2(n7), .O(n432) );
  NAND_GATE U537 ( .I1(n404), .I2(EI_instr[9]), .O(n431) );
  NAND_GATE U538 ( .I1(data2[9]), .I2(n405), .O(n430) );
  NAND3_GATE U539 ( .I1(n433), .I2(n434), .I3(n435), .O(n886) );
  NAND_GATE U540 ( .I1(DI_op2[10]), .I2(n7), .O(n435) );
  NAND_GATE U541 ( .I1(n404), .I2(EI_instr[10]), .O(n434) );
  NAND_GATE U542 ( .I1(data2[10]), .I2(n405), .O(n433) );
  NAND3_GATE U543 ( .I1(n436), .I2(n437), .I3(n438), .O(n887) );
  NAND_GATE U544 ( .I1(DI_op2[11]), .I2(n7), .O(n438) );
  NAND_GATE U545 ( .I1(n404), .I2(EI_instr[11]), .O(n437) );
  NAND_GATE U546 ( .I1(data2[11]), .I2(n405), .O(n436) );
  NAND3_GATE U547 ( .I1(n439), .I2(n440), .I3(n441), .O(n888) );
  NAND_GATE U548 ( .I1(DI_op2[12]), .I2(n7), .O(n441) );
  NAND_GATE U549 ( .I1(n404), .I2(EI_instr[12]), .O(n440) );
  NAND_GATE U550 ( .I1(data2[12]), .I2(n405), .O(n439) );
  NAND3_GATE U551 ( .I1(n442), .I2(n443), .I3(n444), .O(n889) );
  NAND_GATE U552 ( .I1(DI_op2[13]), .I2(n7), .O(n444) );
  NAND_GATE U553 ( .I1(n404), .I2(EI_instr[13]), .O(n443) );
  NAND_GATE U554 ( .I1(data2[13]), .I2(n405), .O(n442) );
  NAND3_GATE U555 ( .I1(n445), .I2(n446), .I3(n447), .O(n890) );
  NAND_GATE U556 ( .I1(DI_op2[14]), .I2(n6), .O(n447) );
  NAND_GATE U557 ( .I1(n404), .I2(EI_instr[14]), .O(n446) );
  NAND_GATE U558 ( .I1(data2[14]), .I2(n405), .O(n445) );
  NAND3_GATE U559 ( .I1(n448), .I2(n449), .I3(n450), .O(n891) );
  NAND_GATE U560 ( .I1(DI_op2[15]), .I2(n6), .O(n450) );
  NAND_GATE U561 ( .I1(n404), .I2(EI_instr[15]), .O(n449) );
  NAND_GATE U562 ( .I1(data2[15]), .I2(n405), .O(n448) );
  NAND3_GATE U563 ( .I1(n451), .I2(n452), .I3(n453), .O(n892) );
  NAND_GATE U564 ( .I1(DI_op2[16]), .I2(n6), .O(n453) );
  NAND_GATE U565 ( .I1(data2[16]), .I2(n405), .O(n451) );
  NAND3_GATE U566 ( .I1(n454), .I2(n452), .I3(n455), .O(n893) );
  NAND_GATE U567 ( .I1(DI_op2[17]), .I2(n6), .O(n455) );
  NAND_GATE U568 ( .I1(data2[17]), .I2(n405), .O(n454) );
  NAND3_GATE U569 ( .I1(n456), .I2(n452), .I3(n457), .O(n894) );
  NAND_GATE U570 ( .I1(DI_op2[18]), .I2(n6), .O(n457) );
  NAND_GATE U571 ( .I1(data2[18]), .I2(n405), .O(n456) );
  NAND3_GATE U572 ( .I1(n458), .I2(n452), .I3(n459), .O(n895) );
  NAND_GATE U573 ( .I1(DI_op2[19]), .I2(n6), .O(n459) );
  NAND_GATE U574 ( .I1(data2[19]), .I2(n405), .O(n458) );
  NAND3_GATE U575 ( .I1(n460), .I2(n452), .I3(n461), .O(n896) );
  NAND_GATE U576 ( .I1(DI_op2[20]), .I2(n6), .O(n461) );
  NAND_GATE U577 ( .I1(data2[20]), .I2(n405), .O(n460) );
  NAND3_GATE U578 ( .I1(n462), .I2(n452), .I3(n463), .O(n897) );
  NAND_GATE U579 ( .I1(DI_op2[21]), .I2(n6), .O(n463) );
  NAND_GATE U580 ( .I1(data2[21]), .I2(n405), .O(n462) );
  NAND3_GATE U581 ( .I1(n464), .I2(n452), .I3(n465), .O(n898) );
  NAND_GATE U582 ( .I1(DI_op2[22]), .I2(n6), .O(n465) );
  NAND_GATE U583 ( .I1(data2[22]), .I2(n405), .O(n464) );
  NAND3_GATE U584 ( .I1(n466), .I2(n452), .I3(n467), .O(n899) );
  NAND_GATE U585 ( .I1(DI_op2[23]), .I2(n5), .O(n467) );
  NAND_GATE U586 ( .I1(data2[23]), .I2(n405), .O(n466) );
  NAND3_GATE U587 ( .I1(n468), .I2(n452), .I3(n469), .O(n900) );
  NAND_GATE U588 ( .I1(DI_op2[24]), .I2(n5), .O(n469) );
  NAND_GATE U589 ( .I1(data2[24]), .I2(n405), .O(n468) );
  NAND3_GATE U590 ( .I1(n470), .I2(n452), .I3(n471), .O(n901) );
  NAND_GATE U591 ( .I1(DI_op2[25]), .I2(n5), .O(n471) );
  NAND_GATE U592 ( .I1(data2[25]), .I2(n405), .O(n470) );
  NAND3_GATE U593 ( .I1(n472), .I2(n452), .I3(n473), .O(n902) );
  NAND_GATE U594 ( .I1(DI_op2[26]), .I2(n5), .O(n473) );
  NAND_GATE U595 ( .I1(data2[26]), .I2(n405), .O(n472) );
  NAND3_GATE U596 ( .I1(n474), .I2(n452), .I3(n475), .O(n903) );
  NAND_GATE U597 ( .I1(DI_op2[27]), .I2(n5), .O(n475) );
  NAND_GATE U598 ( .I1(data2[27]), .I2(n405), .O(n474) );
  NAND3_GATE U599 ( .I1(n476), .I2(n452), .I3(n477), .O(n904) );
  NAND_GATE U600 ( .I1(DI_op2[28]), .I2(n5), .O(n477) );
  NAND_GATE U601 ( .I1(data2[28]), .I2(n405), .O(n476) );
  NAND3_GATE U602 ( .I1(n478), .I2(n452), .I3(n479), .O(n905) );
  NAND_GATE U603 ( .I1(DI_op2[29]), .I2(n5), .O(n479) );
  NAND_GATE U604 ( .I1(data2[29]), .I2(n405), .O(n478) );
  NAND3_GATE U605 ( .I1(n480), .I2(n452), .I3(n481), .O(n906) );
  NAND_GATE U606 ( .I1(DI_op2[30]), .I2(n5), .O(n481) );
  NAND_GATE U607 ( .I1(data2[30]), .I2(n405), .O(n480) );
  NAND3_GATE U608 ( .I1(n482), .I2(n452), .I3(n483), .O(n907) );
  NAND_GATE U609 ( .I1(DI_op2[31]), .I2(n5), .O(n483) );
  NAND3_GATE U610 ( .I1(EI_instr[15]), .I2(n484), .I3(n404), .O(n452) );
  NOR_GATE U611 ( .I1(n195), .I2(n485), .O(n404) );
  NAND_GATE U612 ( .I1(n486), .I2(n487), .O(n484) );
  NAND_GATE U613 ( .I1(n175), .I2(n224), .O(n487) );
  NAND3_GATE U614 ( .I1(n211), .I2(n171), .I3(n53), .O(n486) );
  NAND_GATE U615 ( .I1(data2[31]), .I2(n405), .O(n482) );
  AND_GATE U616 ( .I1(use2), .I2(n203), .O(n405) );
  AND_GATE U617 ( .I1(n485), .I2(n23), .O(use2) );
  AND5_GATE U618 ( .I1(n488), .I2(n489), .I3(n490), .I4(n491), .I5(n492), .O(
        n485) );
  OR_GATE U619 ( .I1(n29), .I2(n42), .O(n492) );
  OR_GATE U620 ( .I1(n200), .I2(n213), .O(n491) );
  OR_GATE U621 ( .I1(n45), .I2(n32), .O(n490) );
  OR_GATE U622 ( .I1(n948), .I2(n944), .O(n45) );
  NAND_GATE U623 ( .I1(n493), .I2(n42), .O(n489) );
  NAND_GATE U624 ( .I1(n494), .I2(n495), .O(n493) );
  NAND_GATE U625 ( .I1(n324), .I2(n49), .O(n495) );
  NAND_GATE U626 ( .I1(n43), .I2(n496), .O(n488) );
  NAND4_GATE U627 ( .I1(n330), .I2(n497), .I3(n498), .I4(n499), .O(n496) );
  OR_GATE U628 ( .I1(n35), .I2(n26), .O(n499) );
  OR_GATE U629 ( .I1(n32), .I2(n70), .O(n498) );
  NOR_GATE U630 ( .I1(n51), .I2(n49), .O(n70) );
  OR_GATE U631 ( .I1(n31), .I2(n49), .O(n497) );
  NAND_GATE U632 ( .I1(n65), .I2(n945), .O(n330) );
  NAND3_GATE U633 ( .I1(n500), .I2(n501), .I3(n502), .O(n908) );
  NAND_GATE U634 ( .I1(DI_op1[0]), .I2(n4), .O(n502) );
  NAND_GATE U635 ( .I1(data1[0]), .I2(n503), .O(n501) );
  NAND_GATE U636 ( .I1(n504), .I2(EI_instr[6]), .O(n500) );
  NAND3_GATE U637 ( .I1(n505), .I2(n506), .I3(n507), .O(n909) );
  NAND_GATE U638 ( .I1(DI_op1[1]), .I2(n4), .O(n507) );
  NAND_GATE U639 ( .I1(data1[1]), .I2(n503), .O(n506) );
  NAND_GATE U640 ( .I1(n504), .I2(EI_instr[7]), .O(n505) );
  NAND3_GATE U641 ( .I1(n508), .I2(n509), .I3(n510), .O(n910) );
  NAND_GATE U642 ( .I1(DI_op1[2]), .I2(n4), .O(n510) );
  NAND_GATE U643 ( .I1(data1[2]), .I2(n503), .O(n509) );
  NAND_GATE U644 ( .I1(n504), .I2(EI_instr[8]), .O(n508) );
  NAND3_GATE U645 ( .I1(n511), .I2(n512), .I3(n513), .O(n911) );
  NAND_GATE U646 ( .I1(DI_op1[3]), .I2(n4), .O(n513) );
  NAND_GATE U647 ( .I1(data1[3]), .I2(n503), .O(n512) );
  NAND_GATE U648 ( .I1(n504), .I2(EI_instr[9]), .O(n511) );
  NAND3_GATE U649 ( .I1(n514), .I2(n515), .I3(n516), .O(n912) );
  NAND_GATE U650 ( .I1(DI_op1[4]), .I2(n4), .O(n516) );
  NAND_GATE U651 ( .I1(data1[4]), .I2(n503), .O(n515) );
  AND_GATE U652 ( .I1(n517), .I2(n21), .O(n503) );
  NAND_GATE U653 ( .I1(n504), .I2(EI_instr[10]), .O(n514) );
  AND_GATE U654 ( .I1(n518), .I2(n21), .O(n504) );
  NAND_GATE U655 ( .I1(n519), .I2(n520), .O(n913) );
  NAND_GATE U656 ( .I1(data1[5]), .I2(n521), .O(n520) );
  NAND_GATE U657 ( .I1(DI_op1[5]), .I2(n4), .O(n519) );
  NAND_GATE U658 ( .I1(n522), .I2(n523), .O(n914) );
  NAND_GATE U659 ( .I1(data1[6]), .I2(n521), .O(n523) );
  NAND_GATE U660 ( .I1(DI_op1[6]), .I2(n4), .O(n522) );
  NAND_GATE U661 ( .I1(n524), .I2(n525), .O(n915) );
  NAND_GATE U662 ( .I1(data1[7]), .I2(n521), .O(n525) );
  NAND_GATE U663 ( .I1(DI_op1[7]), .I2(n4), .O(n524) );
  NAND_GATE U664 ( .I1(n526), .I2(n527), .O(n916) );
  NAND_GATE U665 ( .I1(data1[8]), .I2(n521), .O(n527) );
  NAND_GATE U666 ( .I1(DI_op1[8]), .I2(n4), .O(n526) );
  NAND_GATE U667 ( .I1(n528), .I2(n529), .O(n917) );
  NAND_GATE U668 ( .I1(data1[9]), .I2(n521), .O(n529) );
  NAND_GATE U669 ( .I1(DI_op1[9]), .I2(n3), .O(n528) );
  NAND_GATE U670 ( .I1(n530), .I2(n531), .O(n918) );
  NAND_GATE U671 ( .I1(data1[10]), .I2(n521), .O(n531) );
  NAND_GATE U672 ( .I1(DI_op1[10]), .I2(n3), .O(n530) );
  NAND_GATE U673 ( .I1(n532), .I2(n533), .O(n919) );
  NAND_GATE U674 ( .I1(data1[11]), .I2(n521), .O(n533) );
  NAND_GATE U675 ( .I1(DI_op1[11]), .I2(n3), .O(n532) );
  NAND_GATE U676 ( .I1(n534), .I2(n535), .O(n920) );
  NAND_GATE U677 ( .I1(data1[12]), .I2(n521), .O(n535) );
  NAND_GATE U678 ( .I1(DI_op1[12]), .I2(n3), .O(n534) );
  NAND_GATE U679 ( .I1(n536), .I2(n537), .O(n921) );
  NAND_GATE U680 ( .I1(data1[13]), .I2(n521), .O(n537) );
  NAND_GATE U681 ( .I1(DI_op1[13]), .I2(n3), .O(n536) );
  NAND_GATE U682 ( .I1(n538), .I2(n539), .O(n922) );
  NAND_GATE U683 ( .I1(data1[14]), .I2(n521), .O(n539) );
  NAND_GATE U684 ( .I1(DI_op1[14]), .I2(n3), .O(n538) );
  NAND_GATE U685 ( .I1(n540), .I2(n541), .O(n923) );
  NAND_GATE U686 ( .I1(data1[15]), .I2(n521), .O(n541) );
  NAND_GATE U687 ( .I1(DI_op1[15]), .I2(n3), .O(n540) );
  NAND_GATE U688 ( .I1(n542), .I2(n543), .O(n924) );
  NAND_GATE U689 ( .I1(data1[16]), .I2(n521), .O(n543) );
  NAND_GATE U690 ( .I1(DI_op1[16]), .I2(n3), .O(n542) );
  NAND_GATE U691 ( .I1(n544), .I2(n545), .O(n925) );
  NAND_GATE U692 ( .I1(data1[17]), .I2(n521), .O(n545) );
  NAND_GATE U693 ( .I1(DI_op1[17]), .I2(n3), .O(n544) );
  NAND_GATE U694 ( .I1(n546), .I2(n547), .O(n926) );
  NAND_GATE U695 ( .I1(data1[18]), .I2(n521), .O(n547) );
  NAND_GATE U696 ( .I1(DI_op1[18]), .I2(n2), .O(n546) );
  NAND_GATE U697 ( .I1(n548), .I2(n549), .O(n927) );
  NAND_GATE U698 ( .I1(data1[19]), .I2(n521), .O(n549) );
  NAND_GATE U699 ( .I1(DI_op1[19]), .I2(n2), .O(n548) );
  NAND_GATE U700 ( .I1(n550), .I2(n551), .O(n928) );
  NAND_GATE U701 ( .I1(data1[20]), .I2(n521), .O(n551) );
  NAND_GATE U702 ( .I1(DI_op1[20]), .I2(n2), .O(n550) );
  NAND_GATE U703 ( .I1(n552), .I2(n553), .O(n929) );
  NAND_GATE U704 ( .I1(data1[21]), .I2(n521), .O(n553) );
  NAND_GATE U705 ( .I1(DI_op1[21]), .I2(n2), .O(n552) );
  NAND_GATE U706 ( .I1(n554), .I2(n555), .O(n930) );
  NAND_GATE U707 ( .I1(data1[22]), .I2(n521), .O(n555) );
  NAND_GATE U708 ( .I1(DI_op1[22]), .I2(n2), .O(n554) );
  NAND_GATE U709 ( .I1(n556), .I2(n557), .O(n931) );
  NAND_GATE U710 ( .I1(data1[23]), .I2(n521), .O(n557) );
  NAND_GATE U711 ( .I1(DI_op1[23]), .I2(n2), .O(n556) );
  NAND_GATE U712 ( .I1(n558), .I2(n559), .O(n932) );
  NAND_GATE U713 ( .I1(data1[24]), .I2(n521), .O(n559) );
  NAND_GATE U714 ( .I1(DI_op1[24]), .I2(n2), .O(n558) );
  NAND_GATE U715 ( .I1(n560), .I2(n561), .O(n933) );
  NAND_GATE U716 ( .I1(data1[25]), .I2(n521), .O(n561) );
  NAND_GATE U717 ( .I1(DI_op1[25]), .I2(n2), .O(n560) );
  NAND_GATE U718 ( .I1(n562), .I2(n563), .O(n934) );
  NAND_GATE U719 ( .I1(data1[26]), .I2(n521), .O(n563) );
  NAND_GATE U720 ( .I1(DI_op1[26]), .I2(n2), .O(n562) );
  NAND_GATE U721 ( .I1(n564), .I2(n565), .O(n935) );
  NAND_GATE U722 ( .I1(data1[27]), .I2(n521), .O(n565) );
  NAND_GATE U723 ( .I1(DI_op1[27]), .I2(n1), .O(n564) );
  NAND_GATE U724 ( .I1(n566), .I2(n567), .O(n936) );
  NAND_GATE U725 ( .I1(data1[28]), .I2(n521), .O(n567) );
  NAND_GATE U726 ( .I1(DI_op1[28]), .I2(n1), .O(n566) );
  NAND_GATE U727 ( .I1(n568), .I2(n569), .O(n937) );
  NAND_GATE U728 ( .I1(data1[29]), .I2(n521), .O(n569) );
  NAND_GATE U729 ( .I1(DI_op1[29]), .I2(n1), .O(n568) );
  NAND_GATE U730 ( .I1(n570), .I2(n571), .O(n938) );
  NAND_GATE U731 ( .I1(data1[30]), .I2(n521), .O(n571) );
  NAND_GATE U732 ( .I1(DI_op1[30]), .I2(n1), .O(n570) );
  NAND_GATE U733 ( .I1(n572), .I2(n573), .O(n939) );
  NAND_GATE U734 ( .I1(data1[31]), .I2(n521), .O(n573) );
  AND_GATE U735 ( .I1(n517), .I2(n161), .O(n521) );
  AND4_GATE U736 ( .I1(n574), .I2(n575), .I3(n576), .I4(n577), .O(n517) );
  NOR3_GATE U737 ( .I1(n174), .I2(n518), .I3(n85), .O(n577) );
  AND3_GATE U738 ( .I1(n43), .I2(n944), .I3(n65), .O(n85) );
  AND3_GATE U739 ( .I1(n33), .I2(n42), .I3(n218), .O(n518) );
  AND_GATE U740 ( .I1(n175), .I2(n51), .O(n218) );
  NOR_GATE U741 ( .I1(n948), .I2(n43), .O(n175) );
  NOR_GATE U742 ( .I1(n34), .I2(n944), .O(n173) );
  AND3_GATE U743 ( .I1(n944), .I2(n42), .I3(n64), .O(n174) );
  OR_GATE U744 ( .I1(n31), .I2(n494), .O(n575) );
  AND_GATE U745 ( .I1(n578), .I2(n579), .O(n494) );
  OR_GATE U746 ( .I1(n26), .I2(n48), .O(n579) );
  NAND_GATE U747 ( .I1(n69), .I2(n49), .O(n578) );
  OR_GATE U748 ( .I1(n29), .I2(n34), .O(n574) );
  AND_GATE U749 ( .I1(n69), .I2(n51), .O(n64) );
  NAND_GATE U750 ( .I1(DI_op1[31]), .I2(n1), .O(n572) );
  NAND3_GATE U751 ( .I1(n580), .I2(n581), .I3(n582), .O(n940) );
  NAND_GATE U752 ( .I1(DI_link), .I2(n1), .O(n582) );
  NAND3_GATE U753 ( .I1(n69), .I2(n77), .I3(n355), .O(n581) );
  AND_GATE U754 ( .I1(n21), .I2(n171), .O(n355) );
  OR_GATE U755 ( .I1(n211), .I2(n321), .O(n77) );
  NOR_GATE U756 ( .I1(n213), .I2(n945), .O(n321) );
  NOR_GATE U757 ( .I1(n34), .I2(n42), .O(n211) );
  NAND_GATE U758 ( .I1(n369), .I2(n68), .O(n580) );
  NOR_GATE U759 ( .I1(n34), .I2(n945), .O(n68) );
  AND_GATE U760 ( .I1(n21), .I2(n943), .O(n369) );
  NAND_GATE U761 ( .I1(n203), .I2(n23), .O(n195) );
  AND3_GATE U762 ( .I1(n18), .I2(n19), .I3(n81), .O(n203) );
  NAND_GATE U763 ( .I1(n583), .I2(n584), .O(n941) );
  NAND_GATE U764 ( .I1(n161), .I2(n585), .O(n584) );
  NAND_GATE U765 ( .I1(n160), .I2(n201), .O(n585) );
  NAND_GATE U766 ( .I1(n69), .I2(n171), .O(n201) );
  NOR_GATE U767 ( .I1(n27), .I2(n944), .O(n171) );
  NOR_GATE U768 ( .I1(n363), .I2(n586), .O(n160) );
  AND_GATE U769 ( .I1(n943), .I2(n587), .O(n586) );
  OR_GATE U770 ( .I1(n51), .I2(n213), .O(n587) );
  NAND_GATE U771 ( .I1(n53), .I2(n944), .O(n200) );
  NOR_GATE U772 ( .I1(n948), .I2(n946), .O(n53) );
  AND3_GATE U773 ( .I1(n43), .I2(n49), .I3(n65), .O(n363) );
  AND3_GATE U774 ( .I1(n81), .I2(n23), .I3(n82), .O(n161) );
  NOR_GATE U775 ( .I1(stop_all), .I2(reset), .O(n82) );
  NOR_GATE U776 ( .I1(clear), .I2(stop_di), .O(n81) );
  NAND_GATE U777 ( .I1(DI_bra), .I2(n1), .O(n583) );
  NAND_GATE U778 ( .I1(n588), .I2(n589), .O(n942) );
  OR4_GATE U779 ( .I1(n22), .I2(n1), .I3(clear), .I4(reset), .O(n589) );
  NAND_GATE U780 ( .I1(DI_it_ok), .I2(n1), .O(n588) );
  AND_GATE U781 ( .I1(stop_all), .I2(n19), .O(n72) );
  NAND_GATE U782 ( .I1(n576), .I2(n590), .O(adr_reg2[5]) );
  NAND3_GATE U783 ( .I1(n944), .I2(n945), .I3(n324), .O(n590) );
  AND_GATE U784 ( .I1(n65), .I2(n946), .O(n324) );
  AND3_GATE U785 ( .I1(n27), .I2(n34), .I3(n48), .O(n65) );
  NAND_GATE U786 ( .I1(n67), .I2(n52), .O(n576) );
  NOR_GATE U787 ( .I1(n42), .I2(n213), .O(n52) );
  AND4_GATE U788 ( .I1(n591), .I2(n592), .I3(n593), .I4(n594), .O(n213) );
  AND5_GATE U789 ( .I1(n595), .I2(n596), .I3(n597), .I4(n598), .I5(n599), .O(
        n594) );
  AND5_GATE U790 ( .I1(n600), .I2(n601), .I3(n602), .I4(n603), .I5(n604), .O(
        n593) );
  AND5_GATE U791 ( .I1(n605), .I2(n606), .I3(n607), .I4(n608), .I5(n609), .O(
        n592) );
  AND5_GATE U792 ( .I1(n610), .I2(n611), .I3(n612), .I4(n613), .I5(n614), .O(
        n591) );
  AND4_GATE U793 ( .I1(n615), .I2(n616), .I3(n617), .I4(n618), .O(n42) );
  AND4_GATE U794 ( .I1(n619), .I2(n595), .I3(n599), .I4(n620), .O(n618) );
  AND3_GATE U795 ( .I1(n621), .I2(n622), .I3(n623), .O(n620) );
  AND4_GATE U796 ( .I1(n604), .I2(n624), .I3(n625), .I4(n626), .O(n617) );
  AND3_GATE U797 ( .I1(n627), .I2(n628), .I3(n600), .O(n626) );
  AND5_GATE U798 ( .I1(n629), .I2(n630), .I3(n631), .I4(n632), .I5(n607), .O(
        n616) );
  AND_GATE U799 ( .I1(n633), .I2(n606), .O(n632) );
  NAND_GATE U800 ( .I1(n634), .I2(n635), .O(n606) );
  NAND_GATE U801 ( .I1(n636), .I2(n637), .O(n629) );
  AND5_GATE U802 ( .I1(n638), .I2(n611), .I3(n639), .I4(n640), .I5(n641), .O(
        n615) );
  AND_GATE U803 ( .I1(n612), .I2(n642), .O(n640) );
  NAND3_GATE U804 ( .I1(n643), .I2(n956), .I3(n644), .O(n642) );
  AND_GATE U805 ( .I1(n224), .I2(n69), .O(n67) );
  AND_GATE U806 ( .I1(n43), .I2(n948), .O(n69) );
  AND_GATE U807 ( .I1(n645), .I2(n646), .O(n48) );
  NOR_GATE U808 ( .I1(n51), .I2(n944), .O(n224) );
  AND3_GATE U809 ( .I1(n647), .I2(n648), .I3(n649), .O(n49) );
  AND4_GATE U810 ( .I1(n650), .I2(n651), .I3(n652), .I4(n653), .O(n51) );
  AND3_GATE U811 ( .I1(n654), .I2(n655), .I3(n656), .O(n653) );
  AND_GATE U812 ( .I1(EI_instr[20]), .I2(n23), .O(adr_reg2[4]) );
  AND_GATE U813 ( .I1(EI_instr[19]), .I2(n23), .O(adr_reg2[3]) );
  AND_GATE U814 ( .I1(EI_instr[18]), .I2(n23), .O(adr_reg2[2]) );
  AND_GATE U815 ( .I1(EI_instr[17]), .I2(n23), .O(adr_reg2[1]) );
  AND_GATE U816 ( .I1(EI_instr[16]), .I2(n23), .O(adr_reg2[0]) );
  AND_GATE U817 ( .I1(EI_instr[25]), .I2(n23), .O(adr_reg1[4]) );
  AND_GATE U818 ( .I1(EI_instr[24]), .I2(n23), .O(adr_reg1[3]) );
  AND_GATE U819 ( .I1(EI_instr[23]), .I2(n23), .O(adr_reg1[2]) );
  AND_GATE U820 ( .I1(EI_instr[22]), .I2(n23), .O(adr_reg1[1]) );
  AND_GATE U821 ( .I1(EI_instr[21]), .I2(n23), .O(adr_reg1[0]) );
  AND4_GATE U822 ( .I1(n655), .I2(n646), .I3(n43), .I4(n657), .O(n80) );
  AND4_GATE U823 ( .I1(n648), .I2(n613), .I3(n949), .I4(n622), .O(n657) );
  NAND_GATE U824 ( .I1(n658), .I2(n659), .O(n622) );
  AND_GATE U825 ( .I1(n660), .I2(n621), .O(n613) );
  NAND3_GATE U826 ( .I1(n661), .I2(n956), .I3(n643), .O(n621) );
  NAND_GATE U827 ( .I1(n662), .I2(n659), .O(n660) );
  AND5_GATE U828 ( .I1(n619), .I2(n663), .I3(n597), .I4(n654), .I5(n599), .O(
        n648) );
  NAND_GATE U829 ( .I1(n664), .I2(n658), .O(n599) );
  AND4_GATE U830 ( .I1(n665), .I2(n598), .I3(n628), .I4(n666), .O(n654) );
  NAND_GATE U831 ( .I1(n667), .I2(n658), .O(n666) );
  NAND_GATE U832 ( .I1(n637), .I2(n662), .O(n628) );
  NAND_GATE U833 ( .I1(n634), .I2(n668), .O(n598) );
  NAND_GATE U834 ( .I1(n634), .I2(n664), .O(n665) );
  NAND_GATE U835 ( .I1(n669), .I2(n658), .O(n597) );
  NAND_GATE U836 ( .I1(n662), .I2(n667), .O(n663) );
  AND_GATE U837 ( .I1(n635), .I2(n951), .O(n667) );
  NAND_GATE U838 ( .I1(n669), .I2(n662), .O(n619) );
  AND4_GATE U839 ( .I1(n652), .I2(n645), .I3(n649), .I4(n670), .O(n43) );
  AND3_GATE U840 ( .I1(n630), .I2(n671), .I3(n609), .O(n670) );
  NAND3_GATE U841 ( .I1(n672), .I2(n673), .I3(n636), .O(n609) );
  NAND3_GATE U842 ( .I1(n674), .I2(n956), .I3(n675), .O(n671) );
  NAND_GATE U843 ( .I1(n668), .I2(n662), .O(n630) );
  AND5_GATE U844 ( .I1(n638), .I2(n676), .I3(n677), .I4(n650), .I5(n639), .O(
        n649) );
  NAND_GATE U845 ( .I1(n636), .I2(n669), .O(n639) );
  AND3_GATE U846 ( .I1(n610), .I2(n678), .I3(n612), .O(n650) );
  NAND_GATE U847 ( .I1(n679), .I2(n953), .O(n612) );
  NAND_GATE U848 ( .I1(n644), .I2(n643), .O(n678) );
  NAND_GATE U849 ( .I1(n680), .I2(n662), .O(n610) );
  NAND_GATE U850 ( .I1(n681), .I2(n636), .O(n677) );
  NAND_GATE U851 ( .I1(n681), .I2(n634), .O(n676) );
  NAND_GATE U852 ( .I1(n634), .I2(n669), .O(n638) );
  AND_GATE U853 ( .I1(n682), .I2(n954), .O(n669) );
  AND3_GATE U854 ( .I1(n641), .I2(n683), .I3(n614), .O(n645) );
  NAND3_GATE U855 ( .I1(n658), .I2(n954), .I3(n684), .O(n614) );
  NAND_GATE U856 ( .I1(n636), .I2(n668), .O(n683) );
  NAND3_GATE U857 ( .I1(n685), .I2(n955), .I3(n675), .O(n641) );
  AND4_GATE U858 ( .I1(n611), .I2(n608), .I3(n631), .I4(n686), .O(n652) );
  NAND_GATE U859 ( .I1(n680), .I2(n636), .O(n686) );
  NAND3_GATE U860 ( .I1(n658), .I2(n687), .I3(n684), .O(n631) );
  NAND3_GATE U861 ( .I1(n662), .I2(n687), .I3(n684), .O(n608) );
  NAND_GATE U862 ( .I1(n680), .I2(n634), .O(n611) );
  AND_GATE U863 ( .I1(n688), .I2(n953), .O(n680) );
  AND4_GATE U864 ( .I1(n651), .I2(n600), .I3(n647), .I4(n689), .O(n646) );
  AND3_GATE U865 ( .I1(n627), .I2(n690), .I3(n601), .O(n689) );
  NAND_GATE U866 ( .I1(n634), .I2(n659), .O(n601) );
  AND_GATE U867 ( .I1(n691), .I2(n956), .O(n634) );
  NAND_GATE U868 ( .I1(n681), .I2(n658), .O(n690) );
  NAND_GATE U869 ( .I1(n681), .I2(n662), .O(n627) );
  AND_GATE U870 ( .I1(n682), .I2(n687), .O(n681) );
  AND_GATE U871 ( .I1(n692), .I2(n673), .O(n682) );
  AND4_GATE U872 ( .I1(n656), .I2(n603), .I3(n625), .I4(n693), .O(n647) );
  NAND_GATE U873 ( .I1(n694), .I2(n635), .O(n693) );
  NAND3_GATE U874 ( .I1(n692), .I2(n685), .I3(n695), .O(n625) );
  NAND4_GATE U875 ( .I1(n636), .I2(n696), .I3(n697), .I4(n698), .O(n603) );
  AND4_GATE U876 ( .I1(n607), .I2(n605), .I3(n633), .I4(n699), .O(n656) );
  NAND3_GATE U877 ( .I1(n692), .I2(n956), .I3(n695), .O(n699) );
  AND_GATE U878 ( .I1(n672), .I2(n955), .O(n692) );
  NAND3_GATE U879 ( .I1(n700), .I2(n685), .I3(n695), .O(n633) );
  NAND3_GATE U880 ( .I1(n700), .I2(n956), .I3(n695), .O(n605) );
  AND4_GATE U881 ( .I1(n694), .I2(n691), .I3(n687), .I4(n701), .O(n695) );
  NAND3_GATE U882 ( .I1(n955), .I2(n956), .I3(n675), .O(n607) );
  NAND_GATE U883 ( .I1(n636), .I2(n659), .O(n600) );
  AND_GATE U884 ( .I1(n702), .I2(n687), .O(n659) );
  AND4_GATE U885 ( .I1(n604), .I2(n602), .I3(n624), .I4(n703), .O(n651) );
  NAND3_GATE U886 ( .I1(n662), .I2(n954), .I3(n684), .O(n703) );
  AND3_GATE U887 ( .I1(n955), .I2(n953), .I3(n673), .O(n684) );
  NAND3_GATE U888 ( .I1(n662), .I2(n672), .I3(n688), .O(n624) );
  AND_GATE U889 ( .I1(n644), .I2(n704), .O(n688) );
  AND_GATE U890 ( .I1(n687), .I2(n955), .O(n644) );
  NAND_GATE U891 ( .I1(n679), .I2(n672), .O(n602) );
  AND4_GATE U892 ( .I1(n694), .I2(n661), .I3(n658), .I4(n950), .O(n679) );
  NOR_GATE U893 ( .I1(n698), .I2(n697), .O(n694) );
  NAND_GATE U894 ( .I1(n636), .I2(n664), .O(n604) );
  AND_GATE U895 ( .I1(n691), .I2(n685), .O(n636) );
  AND4_GATE U896 ( .I1(n595), .I2(n596), .I3(n623), .I4(n705), .O(n655) );
  NAND3_GATE U897 ( .I1(n674), .I2(n685), .I3(n675), .O(n705) );
  AND_GATE U898 ( .I1(n643), .I2(n954), .O(n675) );
  AND3_GATE U899 ( .I1(n691), .I2(n672), .I3(n704), .O(n643) );
  AND_GATE U900 ( .I1(n698), .I2(n950), .O(n704) );
  NAND_GATE U901 ( .I1(n668), .I2(n658), .O(n623) );
  AND_GATE U902 ( .I1(n702), .I2(n954), .O(n668) );
  AND_GATE U903 ( .I1(n673), .I2(n700), .O(n702) );
  AND_GATE U904 ( .I1(n674), .I2(n953), .O(n700) );
  NAND_GATE U905 ( .I1(n637), .I2(n658), .O(n596) );
  AND_GATE U906 ( .I1(n685), .I2(n957), .O(n658) );
  AND_GATE U907 ( .I1(n696), .I2(n673), .O(n637) );
  NOR3_GATE U908 ( .I1(n951), .I2(n697), .I3(n950), .O(n673) );
  AND3_GATE U909 ( .I1(n674), .I2(n954), .I3(n672), .O(n696) );
  NAND_GATE U910 ( .I1(n664), .I2(n662), .O(n595) );
  AND_GATE U911 ( .I1(n956), .I2(n957), .O(n662) );
  AND_GATE U912 ( .I1(n706), .I2(n707), .O(n691) );
  OR_GATE U913 ( .I1(n708), .I2(n709), .O(n707) );
  AND_GATE U914 ( .I1(n710), .I2(n711), .O(n685) );
  NAND_GATE U915 ( .I1(n706), .I2(n712), .O(n711) );
  NAND3_GATE U916 ( .I1(n713), .I2(n714), .I3(n715), .O(n712) );
  NAND_GATE U917 ( .I1(EI_instr[0]), .I2(n708), .O(n715) );
  NAND_GATE U918 ( .I1(EI_instr[21]), .I2(n709), .O(n714) );
  NAND_GATE U919 ( .I1(EI_instr[16]), .I2(n716), .O(n713) );
  OR_GATE U920 ( .I1(n958), .I2(n706), .O(n710) );
  AND3_GATE U921 ( .I1(n635), .I2(n698), .I3(n697), .O(n664) );
  AND_GATE U922 ( .I1(n706), .I2(n717), .O(n697) );
  OR_GATE U923 ( .I1(n716), .I2(n709), .O(n717) );
  AND_GATE U924 ( .I1(n718), .I2(n719), .O(n698) );
  NAND_GATE U925 ( .I1(n706), .I2(n720), .O(n719) );
  NAND3_GATE U926 ( .I1(n721), .I2(n722), .I3(n723), .O(n720) );
  NAND_GATE U927 ( .I1(EI_instr[4]), .I2(n708), .O(n723) );
  NAND_GATE U928 ( .I1(EI_instr[25]), .I2(n709), .O(n722) );
  NAND_GATE U929 ( .I1(EI_instr[20]), .I2(n716), .O(n721) );
  NAND_GATE U930 ( .I1(EI_instr[30]), .I2(n952), .O(n718) );
  AND3_GATE U931 ( .I1(n672), .I2(n701), .I3(n661), .O(n635) );
  AND_GATE U932 ( .I1(n687), .I2(n674), .O(n661) );
  NOR_GATE U933 ( .I1(EI_instr[27]), .I2(n724), .O(n674) );
  AND_GATE U934 ( .I1(n706), .I2(n725), .O(n724) );
  NAND3_GATE U935 ( .I1(n726), .I2(n727), .I3(n728), .O(n725) );
  NAND_GATE U936 ( .I1(EI_instr[1]), .I2(n708), .O(n728) );
  NAND_GATE U937 ( .I1(EI_instr[22]), .I2(n709), .O(n727) );
  NAND_GATE U938 ( .I1(EI_instr[17]), .I2(n716), .O(n726) );
  NOR_GATE U939 ( .I1(EI_instr[28]), .I2(n729), .O(n687) );
  AND_GATE U940 ( .I1(n706), .I2(n730), .O(n729) );
  NAND3_GATE U941 ( .I1(n731), .I2(n732), .I3(n733), .O(n730) );
  NAND_GATE U942 ( .I1(EI_instr[2]), .I2(n708), .O(n733) );
  NAND_GATE U943 ( .I1(EI_instr[23]), .I2(n709), .O(n732) );
  NAND_GATE U944 ( .I1(EI_instr[18]), .I2(n716), .O(n731) );
  NOR_GATE U945 ( .I1(EI_instr[31]), .I2(n734), .O(n701) );
  AND3_GATE U946 ( .I1(n708), .I2(n706), .I3(EI_instr[5]), .O(n734) );
  NOR_GATE U947 ( .I1(EI_instr[29]), .I2(n735), .O(n672) );
  AND_GATE U948 ( .I1(n706), .I2(n736), .O(n735) );
  NAND3_GATE U949 ( .I1(n737), .I2(n738), .I3(n739), .O(n736) );
  NAND_GATE U950 ( .I1(EI_instr[3]), .I2(n708), .O(n739) );
  NOR_GATE U951 ( .I1(EI_instr[30]), .I2(EI_instr[26]), .O(n708) );
  NAND_GATE U952 ( .I1(EI_instr[24]), .I2(n709), .O(n738) );
  AND_GATE U953 ( .I1(EI_instr[30]), .I2(n958), .O(n709) );
  NAND_GATE U954 ( .I1(EI_instr[19]), .I2(n716), .O(n737) );
  NOR_GATE U955 ( .I1(n958), .I2(EI_instr[30]), .O(n716) );
  NOR4_GATE U956 ( .I1(EI_instr[28]), .I2(EI_instr[27]), .I3(EI_instr[31]), 
        .I4(EI_instr[29]), .O(n706) );
  INV_GATE U3 ( .I1(n17), .O(n1) );
  INV_GATE U4 ( .I1(n17), .O(n2) );
  INV_GATE U5 ( .I1(n17), .O(n3) );
  INV_GATE U6 ( .I1(n17), .O(n4) );
  INV_GATE U7 ( .I1(n17), .O(n5) );
  INV_GATE U8 ( .I1(n17), .O(n6) );
  INV_GATE U9 ( .I1(n17), .O(n7) );
  INV_GATE U10 ( .I1(n17), .O(n8) );
  INV_GATE U11 ( .I1(n17), .O(n9) );
  INV_GATE U12 ( .I1(n17), .O(n10) );
  INV_GATE U13 ( .I1(n17), .O(n11) );
  INV_GATE U14 ( .I1(n17), .O(n12) );
  INV_GATE U15 ( .I1(n17), .O(n13) );
  INV_GATE U16 ( .I1(n17), .O(n14) );
  INV_GATE U17 ( .I1(n17), .O(n15) );
  INV_GATE U18 ( .I1(n17), .O(n16) );
  INV_GATE U19 ( .I1(n72), .O(n17) );
  INV_GATE U20 ( .I1(n72), .O(n18) );
  INV_GATE U21 ( .I1(reset), .O(n19) );
  INV_GATE U22 ( .I1(n161), .O(n20) );
  INV_GATE U23 ( .I1(n195), .O(n21) );
  INV_GATE U24 ( .I1(EI_it_ok), .O(n22) );
  INV_GATE U25 ( .I1(n80), .O(n23) );
  INV_GATE U26 ( .I1(n315), .O(n24) );
  INV_GATE U27 ( .I1(n202), .O(n25) );
  INV_GATE U28 ( .I1(n171), .O(n26) );
  INV_GATE U29 ( .I1(n51), .O(n27) );
  INV_GATE U30 ( .I1(n67), .O(n28) );
  INV_GATE U31 ( .I1(n64), .O(n29) );
  INV_GATE U32 ( .I1(n174), .O(n30) );
  INV_GATE U33 ( .I1(n68), .O(n31) );
  INV_GATE U34 ( .I1(n211), .O(n32) );
  INV_GATE U35 ( .I1(n173), .O(n33) );
  INV_GATE U36 ( .I1(n213), .O(n34) );
  INV_GATE U957 ( .I1(n321), .O(n35) );
  INV_GATE U958 ( .I1(n200), .O(n943) );
  INV_GATE U959 ( .I1(n49), .O(n944) );
  INV_GATE U960 ( .I1(n42), .O(n945) );
  INV_GATE U961 ( .I1(n43), .O(n946) );
  INV_GATE U962 ( .I1(n175), .O(n947) );
  INV_GATE U963 ( .I1(n48), .O(n948) );
  INV_GATE U964 ( .I1(n643), .O(n949) );
  INV_GATE U965 ( .I1(n701), .O(n950) );
  INV_GATE U966 ( .I1(n698), .O(n951) );
  INV_GATE U967 ( .I1(n706), .O(n952) );
  INV_GATE U968 ( .I1(n672), .O(n953) );
  INV_GATE U969 ( .I1(n687), .O(n954) );
  INV_GATE U970 ( .I1(n674), .O(n955) );
  INV_GATE U971 ( .I1(n685), .O(n956) );
  INV_GATE U972 ( .I1(n691), .O(n957) );
  INV_GATE U973 ( .I1(EI_instr[26]), .O(n958) );
endmodule


module pps_ei ( clock, reset, clear, stop_all, stop_ei, CTE_instr, ETC_adr, 
        PF_pc, EI_instr, EI_adr, EI_it_ok );
  input [31:0] CTE_instr;
  output [31:0] ETC_adr;
  input [31:0] PF_pc;
  output [31:0] EI_instr;
  output [31:0] EI_adr;
  input clock, reset, clear, stop_all, stop_ei;
  output EI_it_ok;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n1, n2;
  assign ETC_adr[31] = PF_pc[31];
  assign ETC_adr[30] = PF_pc[30];
  assign ETC_adr[29] = PF_pc[29];
  assign ETC_adr[28] = PF_pc[28];
  assign ETC_adr[27] = PF_pc[27];
  assign ETC_adr[26] = PF_pc[26];
  assign ETC_adr[25] = PF_pc[25];
  assign ETC_adr[24] = PF_pc[24];
  assign ETC_adr[23] = PF_pc[23];
  assign ETC_adr[22] = PF_pc[22];
  assign ETC_adr[21] = PF_pc[21];
  assign ETC_adr[20] = PF_pc[20];
  assign ETC_adr[19] = PF_pc[19];
  assign ETC_adr[18] = PF_pc[18];
  assign ETC_adr[17] = PF_pc[17];
  assign ETC_adr[16] = PF_pc[16];
  assign ETC_adr[15] = PF_pc[15];
  assign ETC_adr[14] = PF_pc[14];
  assign ETC_adr[13] = PF_pc[13];
  assign ETC_adr[12] = PF_pc[12];
  assign ETC_adr[11] = PF_pc[11];
  assign ETC_adr[10] = PF_pc[10];
  assign ETC_adr[9] = PF_pc[9];
  assign ETC_adr[8] = PF_pc[8];
  assign ETC_adr[7] = PF_pc[7];
  assign ETC_adr[6] = PF_pc[6];
  assign ETC_adr[5] = PF_pc[5];
  assign ETC_adr[4] = PF_pc[4];
  assign ETC_adr[3] = PF_pc[3];
  assign ETC_adr[2] = PF_pc[2];
  assign ETC_adr[1] = PF_pc[1];
  assign ETC_adr[0] = PF_pc[0];

  FLIP_FLOP_D EI_it_ok_reg ( .D(n204), .CK(clock), .Q(EI_it_ok) );
  FLIP_FLOP_D \EI_instr_reg[31]  ( .D(n203), .CK(clock), .Q(EI_instr[31]) );
  FLIP_FLOP_D \EI_instr_reg[30]  ( .D(n202), .CK(clock), .Q(EI_instr[30]) );
  FLIP_FLOP_D \EI_instr_reg[29]  ( .D(n201), .CK(clock), .Q(EI_instr[29]) );
  FLIP_FLOP_D \EI_instr_reg[28]  ( .D(n200), .CK(clock), .Q(EI_instr[28]) );
  FLIP_FLOP_D \EI_instr_reg[27]  ( .D(n199), .CK(clock), .Q(EI_instr[27]) );
  FLIP_FLOP_D \EI_instr_reg[26]  ( .D(n198), .CK(clock), .Q(EI_instr[26]) );
  FLIP_FLOP_D \EI_instr_reg[25]  ( .D(n197), .CK(clock), .Q(EI_instr[25]) );
  FLIP_FLOP_D \EI_instr_reg[24]  ( .D(n196), .CK(clock), .Q(EI_instr[24]) );
  FLIP_FLOP_D \EI_instr_reg[23]  ( .D(n195), .CK(clock), .Q(EI_instr[23]) );
  FLIP_FLOP_D \EI_instr_reg[22]  ( .D(n194), .CK(clock), .Q(EI_instr[22]) );
  FLIP_FLOP_D \EI_instr_reg[21]  ( .D(n193), .CK(clock), .Q(EI_instr[21]) );
  FLIP_FLOP_D \EI_instr_reg[20]  ( .D(n192), .CK(clock), .Q(EI_instr[20]) );
  FLIP_FLOP_D \EI_instr_reg[19]  ( .D(n191), .CK(clock), .Q(EI_instr[19]) );
  FLIP_FLOP_D \EI_instr_reg[18]  ( .D(n190), .CK(clock), .Q(EI_instr[18]) );
  FLIP_FLOP_D \EI_instr_reg[17]  ( .D(n189), .CK(clock), .Q(EI_instr[17]) );
  FLIP_FLOP_D \EI_instr_reg[16]  ( .D(n188), .CK(clock), .Q(EI_instr[16]) );
  FLIP_FLOP_D \EI_instr_reg[15]  ( .D(n187), .CK(clock), .Q(EI_instr[15]) );
  FLIP_FLOP_D \EI_instr_reg[14]  ( .D(n186), .CK(clock), .Q(EI_instr[14]) );
  FLIP_FLOP_D \EI_instr_reg[13]  ( .D(n185), .CK(clock), .Q(EI_instr[13]) );
  FLIP_FLOP_D \EI_instr_reg[12]  ( .D(n184), .CK(clock), .Q(EI_instr[12]) );
  FLIP_FLOP_D \EI_instr_reg[11]  ( .D(n183), .CK(clock), .Q(EI_instr[11]) );
  FLIP_FLOP_D \EI_instr_reg[10]  ( .D(n182), .CK(clock), .Q(EI_instr[10]) );
  FLIP_FLOP_D \EI_instr_reg[9]  ( .D(n181), .CK(clock), .Q(EI_instr[9]) );
  FLIP_FLOP_D \EI_instr_reg[8]  ( .D(n180), .CK(clock), .Q(EI_instr[8]) );
  FLIP_FLOP_D \EI_instr_reg[7]  ( .D(n179), .CK(clock), .Q(EI_instr[7]) );
  FLIP_FLOP_D \EI_instr_reg[6]  ( .D(n178), .CK(clock), .Q(EI_instr[6]) );
  FLIP_FLOP_D \EI_instr_reg[5]  ( .D(n177), .CK(clock), .Q(EI_instr[5]) );
  FLIP_FLOP_D \EI_instr_reg[4]  ( .D(n176), .CK(clock), .Q(EI_instr[4]) );
  FLIP_FLOP_D \EI_instr_reg[3]  ( .D(n175), .CK(clock), .Q(EI_instr[3]) );
  FLIP_FLOP_D \EI_instr_reg[2]  ( .D(n174), .CK(clock), .Q(EI_instr[2]) );
  FLIP_FLOP_D \EI_instr_reg[1]  ( .D(n173), .CK(clock), .Q(EI_instr[1]) );
  FLIP_FLOP_D \EI_instr_reg[0]  ( .D(n172), .CK(clock), .Q(EI_instr[0]) );
  FLIP_FLOP_D \EI_adr_reg[31]  ( .D(n171), .CK(clock), .Q(EI_adr[31]) );
  FLIP_FLOP_D \EI_adr_reg[30]  ( .D(n170), .CK(clock), .Q(EI_adr[30]) );
  FLIP_FLOP_D \EI_adr_reg[29]  ( .D(n169), .CK(clock), .Q(EI_adr[29]) );
  FLIP_FLOP_D \EI_adr_reg[28]  ( .D(n168), .CK(clock), .Q(EI_adr[28]) );
  FLIP_FLOP_D \EI_adr_reg[27]  ( .D(n167), .CK(clock), .Q(EI_adr[27]) );
  FLIP_FLOP_D \EI_adr_reg[26]  ( .D(n166), .CK(clock), .Q(EI_adr[26]) );
  FLIP_FLOP_D \EI_adr_reg[25]  ( .D(n165), .CK(clock), .Q(EI_adr[25]) );
  FLIP_FLOP_D \EI_adr_reg[24]  ( .D(n164), .CK(clock), .Q(EI_adr[24]) );
  FLIP_FLOP_D \EI_adr_reg[23]  ( .D(n163), .CK(clock), .Q(EI_adr[23]) );
  FLIP_FLOP_D \EI_adr_reg[22]  ( .D(n162), .CK(clock), .Q(EI_adr[22]) );
  FLIP_FLOP_D \EI_adr_reg[21]  ( .D(n161), .CK(clock), .Q(EI_adr[21]) );
  FLIP_FLOP_D \EI_adr_reg[20]  ( .D(n160), .CK(clock), .Q(EI_adr[20]) );
  FLIP_FLOP_D \EI_adr_reg[19]  ( .D(n159), .CK(clock), .Q(EI_adr[19]) );
  FLIP_FLOP_D \EI_adr_reg[18]  ( .D(n158), .CK(clock), .Q(EI_adr[18]) );
  FLIP_FLOP_D \EI_adr_reg[17]  ( .D(n157), .CK(clock), .Q(EI_adr[17]) );
  FLIP_FLOP_D \EI_adr_reg[16]  ( .D(n156), .CK(clock), .Q(EI_adr[16]) );
  FLIP_FLOP_D \EI_adr_reg[15]  ( .D(n155), .CK(clock), .Q(EI_adr[15]) );
  FLIP_FLOP_D \EI_adr_reg[14]  ( .D(n154), .CK(clock), .Q(EI_adr[14]) );
  FLIP_FLOP_D \EI_adr_reg[13]  ( .D(n153), .CK(clock), .Q(EI_adr[13]) );
  FLIP_FLOP_D \EI_adr_reg[12]  ( .D(n152), .CK(clock), .Q(EI_adr[12]) );
  FLIP_FLOP_D \EI_adr_reg[11]  ( .D(n151), .CK(clock), .Q(EI_adr[11]) );
  FLIP_FLOP_D \EI_adr_reg[10]  ( .D(n150), .CK(clock), .Q(EI_adr[10]) );
  FLIP_FLOP_D \EI_adr_reg[9]  ( .D(n149), .CK(clock), .Q(EI_adr[9]) );
  FLIP_FLOP_D \EI_adr_reg[8]  ( .D(n148), .CK(clock), .Q(EI_adr[8]) );
  FLIP_FLOP_D \EI_adr_reg[7]  ( .D(n147), .CK(clock), .Q(EI_adr[7]) );
  FLIP_FLOP_D \EI_adr_reg[6]  ( .D(n146), .CK(clock), .Q(EI_adr[6]) );
  FLIP_FLOP_D \EI_adr_reg[5]  ( .D(n145), .CK(clock), .Q(EI_adr[5]) );
  FLIP_FLOP_D \EI_adr_reg[4]  ( .D(n144), .CK(clock), .Q(EI_adr[4]) );
  FLIP_FLOP_D \EI_adr_reg[3]  ( .D(n143), .CK(clock), .Q(EI_adr[3]) );
  FLIP_FLOP_D \EI_adr_reg[2]  ( .D(n142), .CK(clock), .Q(EI_adr[2]) );
  FLIP_FLOP_D \EI_adr_reg[1]  ( .D(n141), .CK(clock), .Q(EI_adr[1]) );
  FLIP_FLOP_D \EI_adr_reg[0]  ( .D(n140), .CK(clock), .Q(EI_adr[0]) );
  NAND_GATE U5 ( .I1(n4), .I2(n5), .O(n140) );
  NAND_GATE U6 ( .I1(PF_pc[0]), .I2(n6), .O(n5) );
  NAND_GATE U7 ( .I1(EI_adr[0]), .I2(n7), .O(n4) );
  NAND_GATE U8 ( .I1(n8), .I2(n9), .O(n141) );
  NAND_GATE U9 ( .I1(PF_pc[1]), .I2(n6), .O(n9) );
  NAND_GATE U10 ( .I1(EI_adr[1]), .I2(n7), .O(n8) );
  NAND_GATE U11 ( .I1(n10), .I2(n11), .O(n142) );
  NAND_GATE U12 ( .I1(PF_pc[2]), .I2(n6), .O(n11) );
  NAND_GATE U13 ( .I1(EI_adr[2]), .I2(n7), .O(n10) );
  NAND_GATE U14 ( .I1(n12), .I2(n13), .O(n143) );
  NAND_GATE U15 ( .I1(PF_pc[3]), .I2(n6), .O(n13) );
  NAND_GATE U16 ( .I1(EI_adr[3]), .I2(n7), .O(n12) );
  NAND_GATE U17 ( .I1(n14), .I2(n15), .O(n144) );
  NAND_GATE U18 ( .I1(PF_pc[4]), .I2(n6), .O(n15) );
  NAND_GATE U19 ( .I1(EI_adr[4]), .I2(n7), .O(n14) );
  NAND_GATE U20 ( .I1(n16), .I2(n17), .O(n145) );
  NAND_GATE U21 ( .I1(PF_pc[5]), .I2(n6), .O(n17) );
  NAND_GATE U22 ( .I1(EI_adr[5]), .I2(n7), .O(n16) );
  NAND_GATE U23 ( .I1(n18), .I2(n19), .O(n146) );
  NAND_GATE U24 ( .I1(PF_pc[6]), .I2(n6), .O(n19) );
  NAND_GATE U25 ( .I1(EI_adr[6]), .I2(n7), .O(n18) );
  NAND_GATE U26 ( .I1(n20), .I2(n21), .O(n147) );
  NAND_GATE U27 ( .I1(PF_pc[7]), .I2(n6), .O(n21) );
  NAND_GATE U28 ( .I1(EI_adr[7]), .I2(n7), .O(n20) );
  NAND_GATE U29 ( .I1(n22), .I2(n23), .O(n148) );
  NAND_GATE U30 ( .I1(PF_pc[8]), .I2(n6), .O(n23) );
  NAND_GATE U31 ( .I1(EI_adr[8]), .I2(n7), .O(n22) );
  NAND_GATE U32 ( .I1(n24), .I2(n25), .O(n149) );
  NAND_GATE U33 ( .I1(PF_pc[9]), .I2(n6), .O(n25) );
  NAND_GATE U34 ( .I1(EI_adr[9]), .I2(n7), .O(n24) );
  NAND_GATE U35 ( .I1(n26), .I2(n27), .O(n150) );
  NAND_GATE U36 ( .I1(PF_pc[10]), .I2(n6), .O(n27) );
  NAND_GATE U37 ( .I1(EI_adr[10]), .I2(n7), .O(n26) );
  NAND_GATE U38 ( .I1(n28), .I2(n29), .O(n151) );
  NAND_GATE U39 ( .I1(PF_pc[11]), .I2(n6), .O(n29) );
  NAND_GATE U40 ( .I1(EI_adr[11]), .I2(n7), .O(n28) );
  NAND_GATE U41 ( .I1(n30), .I2(n31), .O(n152) );
  NAND_GATE U42 ( .I1(PF_pc[12]), .I2(n6), .O(n31) );
  NAND_GATE U43 ( .I1(EI_adr[12]), .I2(n7), .O(n30) );
  NAND_GATE U44 ( .I1(n32), .I2(n33), .O(n153) );
  NAND_GATE U45 ( .I1(PF_pc[13]), .I2(n6), .O(n33) );
  NAND_GATE U46 ( .I1(EI_adr[13]), .I2(n7), .O(n32) );
  NAND_GATE U47 ( .I1(n34), .I2(n35), .O(n154) );
  NAND_GATE U48 ( .I1(PF_pc[14]), .I2(n6), .O(n35) );
  NAND_GATE U49 ( .I1(EI_adr[14]), .I2(n7), .O(n34) );
  NAND_GATE U50 ( .I1(n36), .I2(n37), .O(n155) );
  NAND_GATE U51 ( .I1(PF_pc[15]), .I2(n6), .O(n37) );
  NAND_GATE U52 ( .I1(EI_adr[15]), .I2(n7), .O(n36) );
  NAND_GATE U53 ( .I1(n38), .I2(n39), .O(n156) );
  NAND_GATE U54 ( .I1(PF_pc[16]), .I2(n6), .O(n39) );
  NAND_GATE U55 ( .I1(EI_adr[16]), .I2(n7), .O(n38) );
  NAND_GATE U56 ( .I1(n40), .I2(n41), .O(n157) );
  NAND_GATE U57 ( .I1(PF_pc[17]), .I2(n6), .O(n41) );
  NAND_GATE U58 ( .I1(EI_adr[17]), .I2(n7), .O(n40) );
  NAND_GATE U59 ( .I1(n42), .I2(n43), .O(n158) );
  NAND_GATE U60 ( .I1(PF_pc[18]), .I2(n6), .O(n43) );
  NAND_GATE U61 ( .I1(EI_adr[18]), .I2(n7), .O(n42) );
  NAND_GATE U62 ( .I1(n44), .I2(n45), .O(n159) );
  NAND_GATE U63 ( .I1(PF_pc[19]), .I2(n6), .O(n45) );
  NAND_GATE U64 ( .I1(EI_adr[19]), .I2(n7), .O(n44) );
  NAND_GATE U65 ( .I1(n46), .I2(n47), .O(n160) );
  NAND_GATE U66 ( .I1(PF_pc[20]), .I2(n6), .O(n47) );
  NAND_GATE U67 ( .I1(EI_adr[20]), .I2(n7), .O(n46) );
  NAND_GATE U68 ( .I1(n48), .I2(n49), .O(n161) );
  NAND_GATE U69 ( .I1(PF_pc[21]), .I2(n6), .O(n49) );
  NAND_GATE U70 ( .I1(EI_adr[21]), .I2(n7), .O(n48) );
  NAND_GATE U71 ( .I1(n50), .I2(n51), .O(n162) );
  NAND_GATE U72 ( .I1(PF_pc[22]), .I2(n6), .O(n51) );
  NAND_GATE U73 ( .I1(EI_adr[22]), .I2(n7), .O(n50) );
  NAND_GATE U74 ( .I1(n52), .I2(n53), .O(n163) );
  NAND_GATE U75 ( .I1(PF_pc[23]), .I2(n6), .O(n53) );
  NAND_GATE U76 ( .I1(EI_adr[23]), .I2(n7), .O(n52) );
  NAND_GATE U77 ( .I1(n54), .I2(n55), .O(n164) );
  NAND_GATE U78 ( .I1(PF_pc[24]), .I2(n6), .O(n55) );
  NAND_GATE U79 ( .I1(EI_adr[24]), .I2(n7), .O(n54) );
  NAND_GATE U80 ( .I1(n56), .I2(n57), .O(n165) );
  NAND_GATE U81 ( .I1(PF_pc[25]), .I2(n6), .O(n57) );
  NAND_GATE U82 ( .I1(EI_adr[25]), .I2(n7), .O(n56) );
  NAND_GATE U83 ( .I1(n58), .I2(n59), .O(n166) );
  NAND_GATE U84 ( .I1(PF_pc[26]), .I2(n6), .O(n59) );
  NAND_GATE U85 ( .I1(EI_adr[26]), .I2(n7), .O(n58) );
  NAND_GATE U86 ( .I1(n60), .I2(n61), .O(n167) );
  NAND_GATE U87 ( .I1(PF_pc[27]), .I2(n6), .O(n61) );
  NAND_GATE U88 ( .I1(EI_adr[27]), .I2(n7), .O(n60) );
  NAND_GATE U89 ( .I1(n62), .I2(n63), .O(n168) );
  NAND_GATE U90 ( .I1(PF_pc[28]), .I2(n6), .O(n63) );
  NAND_GATE U91 ( .I1(EI_adr[28]), .I2(n7), .O(n62) );
  NAND_GATE U92 ( .I1(n64), .I2(n65), .O(n169) );
  NAND_GATE U93 ( .I1(PF_pc[29]), .I2(n6), .O(n65) );
  NAND_GATE U94 ( .I1(EI_adr[29]), .I2(n7), .O(n64) );
  NAND_GATE U95 ( .I1(n66), .I2(n67), .O(n170) );
  NAND_GATE U96 ( .I1(PF_pc[30]), .I2(n6), .O(n67) );
  NAND_GATE U97 ( .I1(EI_adr[30]), .I2(n7), .O(n66) );
  NAND_GATE U98 ( .I1(n68), .I2(n69), .O(n171) );
  NAND_GATE U99 ( .I1(PF_pc[31]), .I2(n6), .O(n69) );
  NOR_GATE U100 ( .I1(n7), .I2(reset), .O(n6) );
  NAND_GATE U101 ( .I1(EI_adr[31]), .I2(n7), .O(n68) );
  AND_GATE U102 ( .I1(n1), .I2(n70), .O(n7) );
  OR3_GATE U103 ( .I1(stop_ei), .I2(stop_all), .I3(clear), .O(n70) );
  NAND_GATE U104 ( .I1(n71), .I2(n72), .O(n172) );
  NAND_GATE U105 ( .I1(CTE_instr[0]), .I2(n73), .O(n72) );
  NAND_GATE U106 ( .I1(EI_instr[0]), .I2(n74), .O(n71) );
  NAND_GATE U107 ( .I1(n75), .I2(n76), .O(n173) );
  NAND_GATE U108 ( .I1(CTE_instr[1]), .I2(n73), .O(n76) );
  NAND_GATE U109 ( .I1(EI_instr[1]), .I2(n74), .O(n75) );
  NAND_GATE U110 ( .I1(n77), .I2(n78), .O(n174) );
  NAND_GATE U111 ( .I1(CTE_instr[2]), .I2(n73), .O(n78) );
  NAND_GATE U112 ( .I1(EI_instr[2]), .I2(n74), .O(n77) );
  NAND_GATE U113 ( .I1(n79), .I2(n80), .O(n175) );
  NAND_GATE U114 ( .I1(CTE_instr[3]), .I2(n73), .O(n80) );
  NAND_GATE U115 ( .I1(EI_instr[3]), .I2(n74), .O(n79) );
  NAND_GATE U116 ( .I1(n81), .I2(n82), .O(n176) );
  NAND_GATE U117 ( .I1(CTE_instr[4]), .I2(n73), .O(n82) );
  NAND_GATE U118 ( .I1(EI_instr[4]), .I2(n74), .O(n81) );
  NAND_GATE U119 ( .I1(n83), .I2(n84), .O(n177) );
  NAND_GATE U120 ( .I1(CTE_instr[5]), .I2(n73), .O(n84) );
  NAND_GATE U121 ( .I1(EI_instr[5]), .I2(n74), .O(n83) );
  NAND_GATE U122 ( .I1(n85), .I2(n86), .O(n178) );
  NAND_GATE U123 ( .I1(CTE_instr[6]), .I2(n73), .O(n86) );
  NAND_GATE U124 ( .I1(EI_instr[6]), .I2(n74), .O(n85) );
  NAND_GATE U125 ( .I1(n87), .I2(n88), .O(n179) );
  NAND_GATE U126 ( .I1(CTE_instr[7]), .I2(n73), .O(n88) );
  NAND_GATE U127 ( .I1(EI_instr[7]), .I2(n74), .O(n87) );
  NAND_GATE U128 ( .I1(n89), .I2(n90), .O(n180) );
  NAND_GATE U129 ( .I1(CTE_instr[8]), .I2(n73), .O(n90) );
  NAND_GATE U130 ( .I1(EI_instr[8]), .I2(n74), .O(n89) );
  NAND_GATE U131 ( .I1(n91), .I2(n92), .O(n181) );
  NAND_GATE U132 ( .I1(CTE_instr[9]), .I2(n73), .O(n92) );
  NAND_GATE U133 ( .I1(EI_instr[9]), .I2(n74), .O(n91) );
  NAND_GATE U134 ( .I1(n93), .I2(n94), .O(n182) );
  NAND_GATE U135 ( .I1(CTE_instr[10]), .I2(n73), .O(n94) );
  NAND_GATE U136 ( .I1(EI_instr[10]), .I2(n74), .O(n93) );
  NAND_GATE U137 ( .I1(n95), .I2(n96), .O(n183) );
  NAND_GATE U138 ( .I1(CTE_instr[11]), .I2(n73), .O(n96) );
  NAND_GATE U139 ( .I1(EI_instr[11]), .I2(n74), .O(n95) );
  NAND_GATE U140 ( .I1(n97), .I2(n98), .O(n184) );
  NAND_GATE U141 ( .I1(CTE_instr[12]), .I2(n73), .O(n98) );
  NAND_GATE U142 ( .I1(EI_instr[12]), .I2(n74), .O(n97) );
  NAND_GATE U143 ( .I1(n99), .I2(n100), .O(n185) );
  NAND_GATE U144 ( .I1(CTE_instr[13]), .I2(n73), .O(n100) );
  NAND_GATE U145 ( .I1(EI_instr[13]), .I2(n74), .O(n99) );
  NAND_GATE U146 ( .I1(n101), .I2(n102), .O(n186) );
  NAND_GATE U147 ( .I1(CTE_instr[14]), .I2(n73), .O(n102) );
  NAND_GATE U148 ( .I1(EI_instr[14]), .I2(n74), .O(n101) );
  NAND_GATE U149 ( .I1(n103), .I2(n104), .O(n187) );
  NAND_GATE U150 ( .I1(CTE_instr[15]), .I2(n73), .O(n104) );
  NAND_GATE U151 ( .I1(EI_instr[15]), .I2(n74), .O(n103) );
  NAND_GATE U152 ( .I1(n105), .I2(n106), .O(n188) );
  NAND_GATE U153 ( .I1(CTE_instr[16]), .I2(n73), .O(n106) );
  NAND_GATE U154 ( .I1(EI_instr[16]), .I2(n74), .O(n105) );
  NAND_GATE U155 ( .I1(n107), .I2(n108), .O(n189) );
  NAND_GATE U156 ( .I1(CTE_instr[17]), .I2(n73), .O(n108) );
  NAND_GATE U157 ( .I1(EI_instr[17]), .I2(n74), .O(n107) );
  NAND_GATE U158 ( .I1(n109), .I2(n110), .O(n190) );
  NAND_GATE U159 ( .I1(CTE_instr[18]), .I2(n73), .O(n110) );
  NAND_GATE U160 ( .I1(EI_instr[18]), .I2(n74), .O(n109) );
  NAND_GATE U161 ( .I1(n111), .I2(n112), .O(n191) );
  NAND_GATE U162 ( .I1(CTE_instr[19]), .I2(n73), .O(n112) );
  NAND_GATE U163 ( .I1(EI_instr[19]), .I2(n74), .O(n111) );
  NAND_GATE U164 ( .I1(n113), .I2(n114), .O(n192) );
  NAND_GATE U165 ( .I1(CTE_instr[20]), .I2(n73), .O(n114) );
  NAND_GATE U166 ( .I1(EI_instr[20]), .I2(n74), .O(n113) );
  NAND_GATE U167 ( .I1(n115), .I2(n116), .O(n193) );
  NAND_GATE U168 ( .I1(CTE_instr[21]), .I2(n73), .O(n116) );
  NAND_GATE U169 ( .I1(EI_instr[21]), .I2(n74), .O(n115) );
  NAND_GATE U170 ( .I1(n117), .I2(n118), .O(n194) );
  NAND_GATE U171 ( .I1(CTE_instr[22]), .I2(n73), .O(n118) );
  NAND_GATE U172 ( .I1(EI_instr[22]), .I2(n74), .O(n117) );
  NAND_GATE U173 ( .I1(n119), .I2(n120), .O(n195) );
  NAND_GATE U174 ( .I1(CTE_instr[23]), .I2(n73), .O(n120) );
  NAND_GATE U175 ( .I1(EI_instr[23]), .I2(n74), .O(n119) );
  NAND_GATE U176 ( .I1(n121), .I2(n122), .O(n196) );
  NAND_GATE U177 ( .I1(CTE_instr[24]), .I2(n73), .O(n122) );
  NAND_GATE U178 ( .I1(EI_instr[24]), .I2(n74), .O(n121) );
  NAND_GATE U179 ( .I1(n123), .I2(n124), .O(n197) );
  NAND_GATE U180 ( .I1(CTE_instr[25]), .I2(n73), .O(n124) );
  NAND_GATE U181 ( .I1(EI_instr[25]), .I2(n74), .O(n123) );
  NAND_GATE U182 ( .I1(n125), .I2(n126), .O(n198) );
  NAND_GATE U183 ( .I1(CTE_instr[26]), .I2(n73), .O(n126) );
  NAND_GATE U184 ( .I1(EI_instr[26]), .I2(n74), .O(n125) );
  NAND_GATE U185 ( .I1(n127), .I2(n128), .O(n199) );
  NAND_GATE U186 ( .I1(CTE_instr[27]), .I2(n73), .O(n128) );
  NAND_GATE U187 ( .I1(EI_instr[27]), .I2(n74), .O(n127) );
  NAND_GATE U188 ( .I1(n129), .I2(n130), .O(n200) );
  NAND_GATE U189 ( .I1(CTE_instr[28]), .I2(n73), .O(n130) );
  NAND_GATE U190 ( .I1(EI_instr[28]), .I2(n74), .O(n129) );
  NAND_GATE U191 ( .I1(n131), .I2(n132), .O(n201) );
  NAND_GATE U192 ( .I1(CTE_instr[29]), .I2(n73), .O(n132) );
  NAND_GATE U193 ( .I1(EI_instr[29]), .I2(n74), .O(n131) );
  NAND_GATE U194 ( .I1(n133), .I2(n134), .O(n202) );
  NAND_GATE U195 ( .I1(CTE_instr[30]), .I2(n73), .O(n134) );
  NAND_GATE U196 ( .I1(EI_instr[30]), .I2(n74), .O(n133) );
  NAND_GATE U197 ( .I1(n135), .I2(n136), .O(n203) );
  NAND_GATE U198 ( .I1(CTE_instr[31]), .I2(n73), .O(n136) );
  NAND_GATE U199 ( .I1(EI_instr[31]), .I2(n74), .O(n135) );
  OR_GATE U200 ( .I1(n73), .I2(n137), .O(n204) );
  AND_GATE U201 ( .I1(EI_it_ok), .I2(n74), .O(n137) );
  NOR3_GATE U202 ( .I1(clear), .I2(reset), .I3(n74), .O(n73) );
  AND_GATE U203 ( .I1(n1), .I2(n138), .O(n74) );
  OR_GATE U204 ( .I1(n139), .I2(stop_all), .O(n138) );
  AND_GATE U205 ( .I1(stop_ei), .I2(n2), .O(n139) );
  INV_GATE U3 ( .I1(reset), .O(n1) );
  INV_GATE U4 ( .I1(clear), .O(n2) );
endmodule


module pps_pf ( clock, reset, stop_all, bra_cmd, bra_cmd_pr, bra_adr, exch_cmd, 
        exch_adr, stop_pf, PF_pc );
  input [31:0] bra_adr;
  input [31:0] exch_adr;
  output [31:0] PF_pc;
  input clock, reset, stop_all, bra_cmd, bra_cmd_pr, exch_cmd, stop_pf;
  wire   N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28,
         N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n2, n3, n4, n5;

  FLIP_FLOP_D \pc_interne_reg[0]  ( .D(n175), .CK(clock), .Q(PF_pc[0]) );
  FLIP_FLOP_D \pc_interne_reg[1]  ( .D(n174), .CK(clock), .Q(PF_pc[1]) );
  FLIP_FLOP_D \pc_interne_reg[2]  ( .D(n173), .CK(clock), .Q(PF_pc[2]) );
  FLIP_FLOP_D \pc_interne_reg[3]  ( .D(n172), .CK(clock), .Q(PF_pc[3]) );
  FLIP_FLOP_D \pc_interne_reg[4]  ( .D(n171), .CK(clock), .Q(PF_pc[4]) );
  FLIP_FLOP_D \pc_interne_reg[5]  ( .D(n170), .CK(clock), .Q(PF_pc[5]) );
  FLIP_FLOP_D \pc_interne_reg[6]  ( .D(n169), .CK(clock), .Q(PF_pc[6]) );
  FLIP_FLOP_D \pc_interne_reg[7]  ( .D(n168), .CK(clock), .Q(PF_pc[7]) );
  FLIP_FLOP_D \pc_interne_reg[8]  ( .D(n167), .CK(clock), .Q(PF_pc[8]) );
  FLIP_FLOP_D \pc_interne_reg[9]  ( .D(n166), .CK(clock), .Q(PF_pc[9]) );
  FLIP_FLOP_D \pc_interne_reg[10]  ( .D(n165), .CK(clock), .Q(PF_pc[10]) );
  FLIP_FLOP_D \pc_interne_reg[11]  ( .D(n164), .CK(clock), .Q(PF_pc[11]) );
  FLIP_FLOP_D \pc_interne_reg[12]  ( .D(n163), .CK(clock), .Q(PF_pc[12]) );
  FLIP_FLOP_D \pc_interne_reg[13]  ( .D(n162), .CK(clock), .Q(PF_pc[13]) );
  FLIP_FLOP_D \pc_interne_reg[14]  ( .D(n161), .CK(clock), .Q(PF_pc[14]) );
  FLIP_FLOP_D \pc_interne_reg[15]  ( .D(n160), .CK(clock), .Q(PF_pc[15]) );
  FLIP_FLOP_D \pc_interne_reg[16]  ( .D(n159), .CK(clock), .Q(PF_pc[16]) );
  FLIP_FLOP_D \pc_interne_reg[17]  ( .D(n158), .CK(clock), .Q(PF_pc[17]) );
  FLIP_FLOP_D \pc_interne_reg[18]  ( .D(n157), .CK(clock), .Q(PF_pc[18]) );
  FLIP_FLOP_D \pc_interne_reg[19]  ( .D(n156), .CK(clock), .Q(PF_pc[19]) );
  FLIP_FLOP_D \pc_interne_reg[20]  ( .D(n155), .CK(clock), .Q(PF_pc[20]) );
  FLIP_FLOP_D \pc_interne_reg[21]  ( .D(n154), .CK(clock), .Q(PF_pc[21]) );
  FLIP_FLOP_D \pc_interne_reg[22]  ( .D(n153), .CK(clock), .Q(PF_pc[22]) );
  FLIP_FLOP_D \pc_interne_reg[23]  ( .D(n152), .CK(clock), .Q(PF_pc[23]) );
  FLIP_FLOP_D \pc_interne_reg[24]  ( .D(n151), .CK(clock), .Q(PF_pc[24]) );
  FLIP_FLOP_D \pc_interne_reg[25]  ( .D(n150), .CK(clock), .Q(PF_pc[25]) );
  FLIP_FLOP_D \pc_interne_reg[26]  ( .D(n149), .CK(clock), .Q(PF_pc[26]) );
  FLIP_FLOP_D \pc_interne_reg[27]  ( .D(n148), .CK(clock), .Q(PF_pc[27]) );
  FLIP_FLOP_D \pc_interne_reg[28]  ( .D(n147), .CK(clock), .Q(PF_pc[28]) );
  FLIP_FLOP_D \pc_interne_reg[29]  ( .D(n146), .CK(clock), .Q(PF_pc[29]) );
  FLIP_FLOP_D \pc_interne_reg[30]  ( .D(n145), .CK(clock), .Q(PF_pc[30]) );
  FLIP_FLOP_D \pc_interne_reg[31]  ( .D(n144), .CK(clock), .Q(PF_pc[31]) );
  NAND4_GATE U8 ( .I1(n8), .I2(n9), .I3(n10), .I4(n11), .O(n144) );
  NAND_GATE U9 ( .I1(N46), .I2(n12), .O(n11) );
  NAND_GATE U10 ( .I1(bra_adr[31]), .I2(n13), .O(n10) );
  NAND_GATE U11 ( .I1(exch_adr[31]), .I2(n14), .O(n9) );
  NAND_GATE U12 ( .I1(PF_pc[31]), .I2(n15), .O(n8) );
  NAND4_GATE U13 ( .I1(n16), .I2(n17), .I3(n18), .I4(n19), .O(n145) );
  NAND_GATE U14 ( .I1(N45), .I2(n12), .O(n19) );
  NAND_GATE U15 ( .I1(bra_adr[30]), .I2(n13), .O(n18) );
  NAND_GATE U16 ( .I1(exch_adr[30]), .I2(n14), .O(n17) );
  NAND_GATE U17 ( .I1(PF_pc[30]), .I2(n15), .O(n16) );
  NAND4_GATE U18 ( .I1(n20), .I2(n21), .I3(n22), .I4(n23), .O(n146) );
  NAND_GATE U19 ( .I1(N44), .I2(n12), .O(n23) );
  NAND_GATE U20 ( .I1(bra_adr[29]), .I2(n13), .O(n22) );
  NAND_GATE U21 ( .I1(exch_adr[29]), .I2(n14), .O(n21) );
  NAND_GATE U22 ( .I1(PF_pc[29]), .I2(n15), .O(n20) );
  NAND4_GATE U23 ( .I1(n24), .I2(n25), .I3(n26), .I4(n27), .O(n147) );
  NAND_GATE U24 ( .I1(N43), .I2(n12), .O(n27) );
  NAND_GATE U25 ( .I1(bra_adr[28]), .I2(n13), .O(n26) );
  NAND_GATE U26 ( .I1(exch_adr[28]), .I2(n14), .O(n25) );
  NAND_GATE U27 ( .I1(PF_pc[28]), .I2(n15), .O(n24) );
  NAND4_GATE U28 ( .I1(n28), .I2(n29), .I3(n30), .I4(n31), .O(n148) );
  NAND_GATE U29 ( .I1(N42), .I2(n12), .O(n31) );
  NAND_GATE U30 ( .I1(bra_adr[27]), .I2(n13), .O(n30) );
  NAND_GATE U31 ( .I1(exch_adr[27]), .I2(n14), .O(n29) );
  NAND_GATE U32 ( .I1(PF_pc[27]), .I2(n15), .O(n28) );
  NAND4_GATE U33 ( .I1(n32), .I2(n33), .I3(n34), .I4(n35), .O(n149) );
  NAND_GATE U34 ( .I1(N41), .I2(n12), .O(n35) );
  NAND_GATE U35 ( .I1(bra_adr[26]), .I2(n13), .O(n34) );
  NAND_GATE U36 ( .I1(exch_adr[26]), .I2(n14), .O(n33) );
  NAND_GATE U37 ( .I1(PF_pc[26]), .I2(n15), .O(n32) );
  NAND4_GATE U38 ( .I1(n36), .I2(n37), .I3(n38), .I4(n39), .O(n150) );
  NAND_GATE U39 ( .I1(N40), .I2(n12), .O(n39) );
  NAND_GATE U40 ( .I1(bra_adr[25]), .I2(n13), .O(n38) );
  NAND_GATE U41 ( .I1(exch_adr[25]), .I2(n14), .O(n37) );
  NAND_GATE U42 ( .I1(PF_pc[25]), .I2(n15), .O(n36) );
  NAND4_GATE U43 ( .I1(n40), .I2(n41), .I3(n42), .I4(n43), .O(n151) );
  NAND_GATE U44 ( .I1(N39), .I2(n12), .O(n43) );
  NAND_GATE U45 ( .I1(bra_adr[24]), .I2(n13), .O(n42) );
  NAND_GATE U46 ( .I1(exch_adr[24]), .I2(n14), .O(n41) );
  NAND_GATE U47 ( .I1(PF_pc[24]), .I2(n15), .O(n40) );
  NAND4_GATE U48 ( .I1(n44), .I2(n45), .I3(n46), .I4(n47), .O(n152) );
  NAND_GATE U49 ( .I1(N38), .I2(n12), .O(n47) );
  NAND_GATE U50 ( .I1(bra_adr[23]), .I2(n13), .O(n46) );
  NAND_GATE U51 ( .I1(exch_adr[23]), .I2(n14), .O(n45) );
  NAND_GATE U52 ( .I1(PF_pc[23]), .I2(n15), .O(n44) );
  NAND4_GATE U53 ( .I1(n48), .I2(n49), .I3(n50), .I4(n51), .O(n153) );
  NAND_GATE U54 ( .I1(N37), .I2(n12), .O(n51) );
  NAND_GATE U55 ( .I1(bra_adr[22]), .I2(n13), .O(n50) );
  NAND_GATE U56 ( .I1(exch_adr[22]), .I2(n14), .O(n49) );
  NAND_GATE U57 ( .I1(PF_pc[22]), .I2(n15), .O(n48) );
  NAND4_GATE U58 ( .I1(n52), .I2(n53), .I3(n54), .I4(n55), .O(n154) );
  NAND_GATE U59 ( .I1(N36), .I2(n12), .O(n55) );
  NAND_GATE U60 ( .I1(bra_adr[21]), .I2(n13), .O(n54) );
  NAND_GATE U61 ( .I1(exch_adr[21]), .I2(n14), .O(n53) );
  NAND_GATE U62 ( .I1(PF_pc[21]), .I2(n15), .O(n52) );
  NAND4_GATE U63 ( .I1(n56), .I2(n57), .I3(n58), .I4(n59), .O(n155) );
  NAND_GATE U64 ( .I1(N35), .I2(n12), .O(n59) );
  NAND_GATE U65 ( .I1(bra_adr[20]), .I2(n13), .O(n58) );
  NAND_GATE U66 ( .I1(exch_adr[20]), .I2(n14), .O(n57) );
  NAND_GATE U67 ( .I1(PF_pc[20]), .I2(n15), .O(n56) );
  NAND4_GATE U68 ( .I1(n60), .I2(n61), .I3(n62), .I4(n63), .O(n156) );
  NAND_GATE U69 ( .I1(N34), .I2(n12), .O(n63) );
  NAND_GATE U70 ( .I1(bra_adr[19]), .I2(n13), .O(n62) );
  NAND_GATE U71 ( .I1(exch_adr[19]), .I2(n14), .O(n61) );
  NAND_GATE U72 ( .I1(PF_pc[19]), .I2(n15), .O(n60) );
  NAND4_GATE U73 ( .I1(n64), .I2(n65), .I3(n66), .I4(n67), .O(n157) );
  NAND_GATE U74 ( .I1(N33), .I2(n12), .O(n67) );
  NAND_GATE U75 ( .I1(bra_adr[18]), .I2(n13), .O(n66) );
  NAND_GATE U76 ( .I1(exch_adr[18]), .I2(n14), .O(n65) );
  NAND_GATE U77 ( .I1(PF_pc[18]), .I2(n15), .O(n64) );
  NAND4_GATE U78 ( .I1(n68), .I2(n69), .I3(n70), .I4(n71), .O(n158) );
  NAND_GATE U79 ( .I1(N32), .I2(n12), .O(n71) );
  NAND_GATE U80 ( .I1(bra_adr[17]), .I2(n13), .O(n70) );
  NAND_GATE U81 ( .I1(exch_adr[17]), .I2(n14), .O(n69) );
  NAND_GATE U82 ( .I1(PF_pc[17]), .I2(n15), .O(n68) );
  NAND4_GATE U83 ( .I1(n72), .I2(n73), .I3(n74), .I4(n75), .O(n159) );
  NAND_GATE U84 ( .I1(N31), .I2(n12), .O(n75) );
  NAND_GATE U85 ( .I1(bra_adr[16]), .I2(n13), .O(n74) );
  NAND_GATE U86 ( .I1(exch_adr[16]), .I2(n14), .O(n73) );
  NAND_GATE U87 ( .I1(PF_pc[16]), .I2(n15), .O(n72) );
  NAND4_GATE U88 ( .I1(n76), .I2(n77), .I3(n78), .I4(n79), .O(n160) );
  NAND_GATE U89 ( .I1(N30), .I2(n12), .O(n79) );
  NAND_GATE U90 ( .I1(bra_adr[15]), .I2(n13), .O(n78) );
  NAND_GATE U91 ( .I1(exch_adr[15]), .I2(n14), .O(n77) );
  NAND_GATE U92 ( .I1(PF_pc[15]), .I2(n15), .O(n76) );
  NAND4_GATE U93 ( .I1(n80), .I2(n81), .I3(n82), .I4(n83), .O(n161) );
  NAND_GATE U94 ( .I1(N29), .I2(n12), .O(n83) );
  NAND_GATE U95 ( .I1(bra_adr[14]), .I2(n13), .O(n82) );
  NAND_GATE U96 ( .I1(exch_adr[14]), .I2(n14), .O(n81) );
  NAND_GATE U97 ( .I1(PF_pc[14]), .I2(n15), .O(n80) );
  NAND4_GATE U98 ( .I1(n84), .I2(n85), .I3(n86), .I4(n87), .O(n162) );
  NAND_GATE U99 ( .I1(N28), .I2(n12), .O(n87) );
  NAND_GATE U100 ( .I1(bra_adr[13]), .I2(n13), .O(n86) );
  NAND_GATE U101 ( .I1(exch_adr[13]), .I2(n14), .O(n85) );
  NAND_GATE U102 ( .I1(PF_pc[13]), .I2(n15), .O(n84) );
  NAND4_GATE U103 ( .I1(n88), .I2(n89), .I3(n90), .I4(n91), .O(n163) );
  NAND_GATE U104 ( .I1(N27), .I2(n12), .O(n91) );
  NAND_GATE U105 ( .I1(bra_adr[12]), .I2(n13), .O(n90) );
  NAND_GATE U106 ( .I1(exch_adr[12]), .I2(n14), .O(n89) );
  NAND_GATE U107 ( .I1(PF_pc[12]), .I2(n15), .O(n88) );
  NAND4_GATE U108 ( .I1(n92), .I2(n93), .I3(n94), .I4(n95), .O(n164) );
  NAND_GATE U109 ( .I1(N26), .I2(n12), .O(n95) );
  NAND_GATE U110 ( .I1(bra_adr[11]), .I2(n13), .O(n94) );
  NAND_GATE U111 ( .I1(exch_adr[11]), .I2(n14), .O(n93) );
  NAND_GATE U112 ( .I1(PF_pc[11]), .I2(n15), .O(n92) );
  NAND4_GATE U113 ( .I1(n96), .I2(n97), .I3(n98), .I4(n99), .O(n165) );
  NAND_GATE U114 ( .I1(N25), .I2(n12), .O(n99) );
  NAND_GATE U115 ( .I1(bra_adr[10]), .I2(n13), .O(n98) );
  NAND_GATE U116 ( .I1(exch_adr[10]), .I2(n14), .O(n97) );
  NAND_GATE U117 ( .I1(PF_pc[10]), .I2(n15), .O(n96) );
  NAND4_GATE U118 ( .I1(n100), .I2(n101), .I3(n102), .I4(n103), .O(n166) );
  NAND_GATE U119 ( .I1(N24), .I2(n12), .O(n103) );
  NAND_GATE U120 ( .I1(bra_adr[9]), .I2(n13), .O(n102) );
  NAND_GATE U121 ( .I1(exch_adr[9]), .I2(n14), .O(n101) );
  NAND_GATE U122 ( .I1(PF_pc[9]), .I2(n15), .O(n100) );
  NAND4_GATE U123 ( .I1(n104), .I2(n105), .I3(n106), .I4(n107), .O(n167) );
  NAND_GATE U124 ( .I1(N23), .I2(n12), .O(n107) );
  NAND_GATE U125 ( .I1(bra_adr[8]), .I2(n13), .O(n106) );
  NAND_GATE U126 ( .I1(exch_adr[8]), .I2(n14), .O(n105) );
  NAND_GATE U127 ( .I1(PF_pc[8]), .I2(n15), .O(n104) );
  NAND4_GATE U128 ( .I1(n108), .I2(n109), .I3(n110), .I4(n111), .O(n168) );
  NAND_GATE U129 ( .I1(N22), .I2(n12), .O(n111) );
  NAND_GATE U130 ( .I1(bra_adr[7]), .I2(n13), .O(n110) );
  NAND_GATE U131 ( .I1(exch_adr[7]), .I2(n14), .O(n109) );
  NAND_GATE U132 ( .I1(PF_pc[7]), .I2(n15), .O(n108) );
  NAND4_GATE U133 ( .I1(n112), .I2(n113), .I3(n114), .I4(n115), .O(n169) );
  NAND_GATE U134 ( .I1(N21), .I2(n12), .O(n115) );
  NAND_GATE U135 ( .I1(bra_adr[6]), .I2(n13), .O(n114) );
  NAND_GATE U136 ( .I1(exch_adr[6]), .I2(n14), .O(n113) );
  NAND_GATE U137 ( .I1(PF_pc[6]), .I2(n15), .O(n112) );
  NAND4_GATE U138 ( .I1(n116), .I2(n117), .I3(n118), .I4(n119), .O(n170) );
  NAND_GATE U139 ( .I1(N20), .I2(n12), .O(n119) );
  NAND_GATE U140 ( .I1(bra_adr[5]), .I2(n13), .O(n118) );
  NAND_GATE U141 ( .I1(exch_adr[5]), .I2(n14), .O(n117) );
  NAND_GATE U142 ( .I1(PF_pc[5]), .I2(n15), .O(n116) );
  NAND4_GATE U143 ( .I1(n120), .I2(n121), .I3(n122), .I4(n123), .O(n171) );
  NAND_GATE U144 ( .I1(N19), .I2(n12), .O(n123) );
  NAND_GATE U145 ( .I1(bra_adr[4]), .I2(n13), .O(n122) );
  NAND_GATE U146 ( .I1(exch_adr[4]), .I2(n14), .O(n121) );
  NAND_GATE U147 ( .I1(PF_pc[4]), .I2(n15), .O(n120) );
  NAND4_GATE U148 ( .I1(n124), .I2(n125), .I3(n126), .I4(n127), .O(n172) );
  NAND_GATE U149 ( .I1(N18), .I2(n12), .O(n127) );
  NAND_GATE U150 ( .I1(bra_adr[3]), .I2(n13), .O(n126) );
  NAND_GATE U151 ( .I1(exch_adr[3]), .I2(n14), .O(n125) );
  NAND_GATE U152 ( .I1(PF_pc[3]), .I2(n15), .O(n124) );
  NAND4_GATE U153 ( .I1(n128), .I2(n129), .I3(n130), .I4(n131), .O(n173) );
  NAND_GATE U154 ( .I1(N17), .I2(n12), .O(n131) );
  NAND_GATE U155 ( .I1(bra_adr[2]), .I2(n13), .O(n130) );
  NAND_GATE U156 ( .I1(exch_adr[2]), .I2(n14), .O(n129) );
  NAND_GATE U157 ( .I1(PF_pc[2]), .I2(n15), .O(n128) );
  NAND4_GATE U158 ( .I1(n132), .I2(n133), .I3(n134), .I4(n135), .O(n174) );
  NAND_GATE U159 ( .I1(N16), .I2(n12), .O(n135) );
  NAND_GATE U160 ( .I1(bra_adr[1]), .I2(n13), .O(n134) );
  NAND_GATE U161 ( .I1(exch_adr[1]), .I2(n14), .O(n133) );
  NAND_GATE U162 ( .I1(PF_pc[1]), .I2(n15), .O(n132) );
  NAND4_GATE U163 ( .I1(n136), .I2(n137), .I3(n138), .I4(n139), .O(n175) );
  NAND_GATE U164 ( .I1(N15), .I2(n12), .O(n139) );
  NOR_GATE U165 ( .I1(n140), .I2(n141), .O(n12) );
  NAND_GATE U166 ( .I1(bra_adr[0]), .I2(n13), .O(n138) );
  NOR_GATE U167 ( .I1(n140), .I2(n3), .O(n13) );
  OR_GATE U168 ( .I1(bra_cmd), .I2(bra_cmd_pr), .O(n141) );
  OR3_GATE U169 ( .I1(exch_cmd), .I2(reset), .I3(n15), .O(n140) );
  NAND_GATE U170 ( .I1(exch_adr[0]), .I2(n14), .O(n137) );
  NOR3_GATE U171 ( .I1(n15), .I2(reset), .I3(n4), .O(n14) );
  NAND_GATE U172 ( .I1(PF_pc[0]), .I2(n15), .O(n136) );
  AND_GATE U173 ( .I1(n2), .I2(n142), .O(n15) );
  OR_GATE U174 ( .I1(n143), .I2(stop_all), .O(n142) );
  NOR3_GATE U175 ( .I1(bra_cmd_pr), .I2(exch_cmd), .I3(n5), .O(n143) );
  pps_pf_DW01_add_0 add_89 ( .A(PF_pc), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({N46, N45, N44, N43, N42, N41, N40, N39, 
        N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, 
        N24, N23, N22, N21, N20, N19, N18, N17, N16, N15}) );
  INV_GATE U3 ( .I1(reset), .O(n2) );
  INV_GATE U4 ( .I1(n141), .O(n3) );
  INV_GATE U6 ( .I1(exch_cmd), .O(n4) );
  INV_GATE U7 ( .I1(stop_pf), .O(n5) );
endmodule


module minimips ( clock, reset, ram_req, ram_adr, ram_r_w, ram_data, ram_ack, 
        it_mat );
  output [31:0] ram_adr;
  inout [31:0] ram_data;
  input clock, reset, ram_ack, it_mat;
  output ram_req, ram_r_w;
  wire   interrupt, PR_clear, clear, it_mat_clk, stop_all, PR_bra_cmd,
         PR_bra_bad, alea, EI_it_ok, use1, use2, DI_bra, DI_link, DI_ecr_reg,
         DI_mode, DI_op_mem, DI_r_w, DI_it_ok, EX_bra_confirm, EX_ecr_reg,
         EX_op_mem, EX_r_w, EX_it_ok, MTC_r_w, MTC_req, MEM_ecr_reg, MEM_it_ok,
         write_GPR, write_SCP;
  wire   [31:0] PR_bra_adr;
  wire   [31:0] vecteur_it;
  wire   [31:0] PF_pc;
  wire   [31:0] CTE_instr;
  wire   [31:0] ETC_adr;
  wire   [31:0] EI_instr;
  wire   [31:0] EI_adr;
  wire   [5:0] adr_reg1;
  wire   [5:0] adr_reg2;
  wire   [31:0] data1;
  wire   [31:0] data2;
  wire   [31:0] DI_op1;
  wire   [31:0] DI_op2;
  wire   [27:0] DI_code_ual;
  wire   [31:0] DI_offset;
  wire   [5:0] DI_adr_reg_dest;
  wire   [31:0] DI_adr;
  wire   [31:0] DI_exc_cause;
  wire   [1:0] DI_level;
  wire   [31:0] EX_adr;
  wire   [31:0] EX_data_ual;
  wire   [31:0] EX_adresse;
  wire   [5:0] EX_adr_reg_dest;
  wire   [31:0] EX_exc_cause;
  wire   [1:0] EX_level;
  wire   [31:0] MTC_data;
  wire   [31:0] MTC_adr;
  wire   [31:0] CTM_data;
  wire   [31:0] MEM_adr;
  wire   [5:0] MEM_adr_reg_dest;
  wire   [31:0] MEM_data_ecr;
  wire   [31:0] MEM_exc_cause;
  wire   [1:0] MEM_level;
  wire   [31:0] write_data;
  wire   [4:0] write_adr;
  wire   [4:0] read_adr1;
  wire   [4:0] read_adr2;
  wire   [31:0] read_data1_GPR;
  wire   [31:0] read_data1_SCP;
  wire   [31:0] read_data2_GPR;
  wire   [31:0] read_data2_SCP;
  tri   [31:0] ram_data;
  wire   SYNOPSYS_UNCONNECTED__0;

  FLIP_FLOP_D it_mat_clk_reg ( .D(it_mat), .CK(clock), .Q(it_mat_clk) );
  OR_GATE U3 ( .I1(PR_clear), .I2(interrupt), .O(clear) );
  pps_pf U1_pf ( .clock(clock), .reset(reset), .stop_all(stop_all), .bra_cmd(
        PR_bra_cmd), .bra_cmd_pr(PR_bra_bad), .bra_adr(PR_bra_adr), .exch_cmd(
        interrupt), .exch_adr(vecteur_it), .stop_pf(alea), .PF_pc(PF_pc) );
  pps_ei U2_ei ( .clock(clock), .reset(reset), .clear(clear), .stop_all(
        stop_all), .stop_ei(alea), .CTE_instr(CTE_instr), .ETC_adr(ETC_adr), 
        .PF_pc(PF_pc), .EI_instr(EI_instr), .EI_adr(EI_adr), .EI_it_ok(
        EI_it_ok) );
  pps_di U3_di ( .clock(clock), .reset(reset), .stop_all(stop_all), .clear(
        clear), .adr_reg1({SYNOPSYS_UNCONNECTED__0, adr_reg1[4:0]}), 
        .adr_reg2(adr_reg2), .use1(use1), .use2(use2), .stop_di(alea), .data1(
        data1), .data2(data2), .EI_adr(EI_adr), .EI_instr(EI_instr), 
        .EI_it_ok(EI_it_ok), .DI_bra(DI_bra), .DI_link(DI_link), .DI_op1(
        DI_op1), .DI_op2(DI_op2), .DI_code_ual(DI_code_ual), .DI_offset(
        DI_offset), .DI_adr_reg_dest(DI_adr_reg_dest), .DI_ecr_reg(DI_ecr_reg), 
        .DI_mode(DI_mode), .DI_op_mem(DI_op_mem), .DI_r_w(DI_r_w), .DI_adr(
        DI_adr), .DI_exc_cause(DI_exc_cause), .DI_level(DI_level), .DI_it_ok(
        DI_it_ok) );
  pps_ex U4_ex ( .clock(clock), .reset(reset), .stop_all(stop_all), .clear(
        clear), .DI_bra(DI_bra), .DI_link(DI_link), .DI_op1(DI_op1), .DI_op2(
        DI_op2), .DI_code_ual(DI_code_ual), .DI_offset(DI_offset), 
        .DI_adr_reg_dest(DI_adr_reg_dest), .DI_ecr_reg(DI_ecr_reg), .DI_mode(
        DI_mode), .DI_op_mem(DI_op_mem), .DI_r_w(DI_r_w), .DI_adr(DI_adr), 
        .DI_exc_cause(DI_exc_cause), .DI_level(DI_level), .DI_it_ok(DI_it_ok), 
        .EX_adr(EX_adr), .EX_bra_confirm(EX_bra_confirm), .EX_data_ual(
        EX_data_ual), .EX_adresse(EX_adresse), .EX_adr_reg_dest(
        EX_adr_reg_dest), .EX_ecr_reg(EX_ecr_reg), .EX_op_mem(EX_op_mem), 
        .EX_r_w(EX_r_w), .EX_exc_cause(EX_exc_cause), .EX_level(EX_level), 
        .EX_it_ok(EX_it_ok) );
  pps_mem U5_mem ( .clock(clock), .reset(reset), .stop_all(stop_all), .clear(
        interrupt), .MTC_data(MTC_data), .MTC_adr(MTC_adr), .MTC_r_w(MTC_r_w), 
        .MTC_req(MTC_req), .CTM_data(CTM_data), .EX_adr(EX_adr), .EX_data_ual(
        EX_data_ual), .EX_adresse(EX_adresse), .EX_adr_reg_dest(
        EX_adr_reg_dest), .EX_ecr_reg(EX_ecr_reg), .EX_op_mem(EX_op_mem), 
        .EX_r_w(EX_r_w), .EX_exc_cause(EX_exc_cause), .EX_level(EX_level), 
        .EX_it_ok(EX_it_ok), .MEM_adr(MEM_adr), .MEM_adr_reg_dest(
        MEM_adr_reg_dest), .MEM_ecr_reg(MEM_ecr_reg), .MEM_data_ecr(
        MEM_data_ecr), .MEM_exc_cause(MEM_exc_cause), .MEM_level(MEM_level), 
        .MEM_it_ok(MEM_it_ok) );
  renvoi U6_renvoi ( .adr1({1'b0, adr_reg1[4:0]}), .adr2(adr_reg2), .use1(use1), .use2(use2), .data1(data1), .data2(data2), .alea(alea), .DI_level(DI_level), 
        .DI_adr(DI_adr_reg_dest), .DI_ecr(DI_ecr_reg), .DI_data(DI_op2), 
        .EX_level(EX_level), .EX_adr(EX_adr_reg_dest), .EX_ecr(EX_ecr_reg), 
        .EX_data(EX_data_ual), .MEM_level(MEM_level), .MEM_adr(
        MEM_adr_reg_dest), .MEM_ecr(MEM_ecr_reg), .MEM_data(MEM_data_ecr), 
        .interrupt(interrupt), .write_data(write_data), .write_adr(write_adr), 
        .write_GPR(write_GPR), .write_SCP(write_SCP), .read_adr1(read_adr1), 
        .read_adr2(read_adr2), .read_data1_GPR(read_data1_GPR), 
        .read_data2_GPR(read_data2_GPR), .read_data1_SCP(read_data1_SCP), 
        .read_data2_SCP(read_data2_SCP) );
  banc U7_banc ( .clock(clock), .reset(reset), .reg_src1(read_adr1), 
        .reg_src2(read_adr2), .reg_dest(write_adr), .donnee(write_data), 
        .cmd_ecr(write_GPR), .data_src1(read_data1_GPR), .data_src2(
        read_data2_GPR) );
  syscop U8_syscop ( .clock(clock), .reset(reset), .MEM_adr(MEM_adr), 
        .MEM_exc_cause(MEM_exc_cause), .MEM_it_ok(MEM_it_ok), .it_mat(
        it_mat_clk), .interrupt(interrupt), .vecteur_it(vecteur_it), 
        .write_data(write_data), .write_adr(write_adr), .write_SCP(write_SCP), 
        .read_adr1(read_adr1), .read_adr2(read_adr2), .read_data1(
        read_data1_SCP), .read_data2(read_data2_SCP) );
  bus_ctrl U9_bus_ctrl ( .clock(clock), .reset(reset), .interrupt(interrupt), 
        .adr_from_ei(ETC_adr), .instr_to_ei(CTE_instr), .req_from_mem(MTC_req), 
        .r_w_from_mem(MTC_r_w), .adr_from_mem(MTC_adr), .data_from_mem(
        MTC_data), .data_to_mem(CTM_data), .req_to_ram(ram_req), .adr_to_ram(
        ram_adr), .r_w_to_ram(ram_r_w), .ack_from_ram(ram_ack), 
        .data_inout_ram(ram_data), .stop_all(stop_all) );
  predict_nb_record3_1 U10_predict ( .clock(clock), .reset(reset), .PF_pc(
        PF_pc), .DI_bra(DI_bra), .DI_adr(DI_adr), .EX_bra_confirm(
        EX_bra_confirm), .EX_adr(EX_adr), .EX_adresse(EX_adresse), 
        .EX_uncleared(EX_it_ok), .PR_bra_cmd(PR_bra_cmd), .PR_bra_bad(
        PR_bra_bad), .PR_bra_adr(PR_bra_adr), .PR_clear(PR_clear) );
endmodule

